`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjEJlbRY3s2UM7QgqMREb1m/j5GRdtBtOXui81RZItJxHDO3J4vDN943yaDWqrFM
bpqKb2GR5Qh8KGyCRs+SLJrI+mOXnpsD8Cv8Kitz7U50yi6XT1TwZSCLXCIbFlXV
HF7O5UkTt7n/Xbqjtd01vOQ2RAPK2Kil/3jPivia2iZiKGNgon/aacBDen04DaZh
t2TVpY+LauzZ3HpccrJSajv1w7Wfanri792zsW5vNyVzeU4kvzu/ZTnXUy37V8+b
hvbnupwDQhkYG331/goKqCBUN0DiIrX5tYwlXy7wLztIKyEML0C+/sVUMs7FLMKs
wpR2VnGFdFR36AeC1Nkhp8sZbSls2O2ywMC2gEsD7q2tUYtZzVtkmnNbC2Mpc4tt
aOu+BlRTYA1cBykmHRAv5f5Ctr6x6M6jrzM0hgPHiJQdoIZejR+ZHbMWiSQczR7C
xxgbhOtNwC78wMOdLiqXvpuW6ByEiXGJx64hWLaafS4QCror0PD3WQHbt8ptIMwm
qbrUyv+/XrbvyDUb+ZaY3fCtAuM7luZxRY29q9h86UGOCOCVjVqSA/Ia24nvwaCx
lbWNjec8QmxNjbW9YapTmmBoXaF2URKNyO3N3bc/Kt3xjFz5l0ewExk4eJZbgI9f
XO1l6cmCu9gKA20gKXMLGpM7LTmjd6pl9OU3LM5Km27QuWW/g2/DH91mFmxQBv2K
3ZA76NHXThE/06kXdsZm8w3PEBSnUBBUPhefsnz/uaM=
`protect END_PROTECTED
