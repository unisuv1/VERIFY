`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oKYqo92xoIqT8UIz3lMvmrw+Xgh3R3d9FYDY0JyJN99n9qQPzuBHcHiAl/TNx8V6
Pgmbl4i/9sXYT/ETT7Rjurd8g5LnBw9TfP2dc+ULmmVCjA/fY0/fIowXE8Udl96A
5QYSDrpKRynSz14Z/j8oQChHQN3lxBjFEubtcihDEV7cYg956/K+bW/FuvNm0q/h
Any5LxiukW44LdX+/+aHZGTbqsgwkuC4Fu9X8a5NTwUxUBWWApw8Fiaar2jHIpmN
4LBONtxygQeh+XyRWyIQi6glrB58nVTe5/HhduckucXp1Som/+/3hmB9R4jWhCCs
R3t+YHrkBySz076Y7b0t5vkl0fEa6N8wWj7uwwM5zkSwzzlzDnxgZEQsx8uTVC66
F5ot0HyRAtEf0okizezxIGwokwLClkid2HAEbJFV6sHSg4FCEejDgYemD6jq3q5e
+JsbhLTRcvXCtBbvzVNPzTEWzDXYwJcv/cir0WJERoCWhHhpSIuMa83YNnp4VFk2
ZGIZXchpm9CuHDSEDcEPzbSwls67thogOAmlwjA/IHrl6C9zXBY4bp3mZkAeIlXN
e7cmF51PdUvAeA5cOFeLcBHiBRRBbjKsTmAi3SGtnOLWOA0ItZAgWb7C9Bif2TJg
kIGOj4ogN0MdACz5spTNcvZFMcIl5A+C4WbXNz4cV1QAvENSHO/NYIrp89V8MQQ9
1RFPWQ/J3S+aDZ7PELgaGBZ2tBHBTU/qxIW/+mpj3geY7JFWtqBj0JEpHzXWzgky
MVKqQetUdjRot2lFLp8HdInbWv5ZZrER6QX6tA2MfHERr2zwA4zf7gSQk+rHDIKN
s2A4N1wqCRvLQHDeF6bgXRv4lki4X9aKLF/+Nbr2H2MFvo6eDLyEj3sNMhuR5sui
a1WfGHAwKd1osrgpnVwsGKbXqh4pWPpWMvF2RYgcel8NXSL223FYb9TjNYjW79uy
ODYvLq4YQh+TNtY97ges8mr3yezn2lFbsuORpUAMWq3DTGQ2RiAtOCxYJbDADpD8
exTAIfqL2mCtWi5irB25oRWCHmKBcf9lNXYGWwDscYknkwKVhJHlVy6EMZ9PasND
ZvspVFtk3j3QME2yhgq1O9QMMtvOS7V2igxTjGVPeicpYRbmJj8PX1vswFR93MNJ
sTddr88M/gOxfgYjcHFF23ibWOt0uPXy1lyht236UbECqtcLlPqxZ7F1NMcfZy0C
3mzeiW+pp3f+lXhyG8x+1EvUIAYrNt2qutkGqXtxaGaotflelHT9bHXzbvIg14ia
NDVyBguhOEBsB+cK1rcAdT4/wvgClMIQqe+6qdEon9cfp4b8lWuhWmUy1NDvrwc8
MiHGeVigO0xmx8O3VpVU6hG6g3uosLDai46/boFtjhXB06xU0hFdzLHsEEHzGFwo
AIYBdStYD+OPmXzcNdVPm8kWGsZV8FO5zamwyDrgMnnmpYyjmANmlgkx+r88Zl21
wNMNjOLyufP9GZyND2kvkvS5l49Mj35zUCGx8TTqE6k=
`protect END_PROTECTED
