`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LDkboZsWLGjHcqt0MwdeKKMZC5hPiQb6dlWvQWgNkDx3WvQv1ty+hh/20IdgF9ij
09CxJfY79MORBuMpEy+09/5RTSFs1NVFNykVjcJektpdsXb10fF6h87zlV8DnJM7
GOihKazFDloRMS5I7ZEBkL2820FjvAFvGQVpr/KDfb4AN0mpgmSKbkrptR+45JPF
cu2i5DAnEnb/NfPLE5D8qgUtAspDo+K2sZtmpiU5Im6srk+ra7FTASDX4WxbenA/
b4/1yTW4CeLin1GvkOZWwbzMFo0XlwOkF/t4ZlB1Mss+Nv7WetBR8il27Zc1fiDE
CrC7vu38yRNb/idPciqgsebwZSV7wKwsjDp69gp85hTDCfBzd4+XJbpIdqhJR/YX
kaGI4I9IK7sxZ+krEahvTJG5XZAkoYpUE/QcqkYqCJtQQ8aSglX5wfGe+uQo+GAm
zQNU/foYaEVwf2NVRPfk6Xo1ds/Gkqtn4uFJmMLkkallCtVzcp7ytz/K9U01gZoj
PVANHL7Sg0sFNMAY2ffC8HehcgnVJ5N+m5Mj+qBHxiUVYYT6h0ib3yiB1PmnfJk3
NEsVNPTnZPGodfI5PGpBMZZPsqsxM3wryCJDT3Y1hqba40KbfaSyr7PTA/s8eM6t
zWpaKwj/Y4oK4v0/nZlLXLX6gQNsTrkCqY4oyjBuDJbjG7m6yIzBlsQQDLWJy4if
acXBeqEtieC0TU+C0jrhOlV3R3L9I6chXmjU5gRtMH5wO851uIJEmlsjwjy/5VL1
rqV+X6h71WYJQ0+6K0vVyzxb8oDxpcF1mBOL67vAI2+uLKRKlz2T1m6PezhIP1bH
sVheUH3A0NlXFNlk1iTjaBndPxJCMZeILLMNqDW5OarE0szoDGwiNwBjF+N/n0AN
ovtJepARtUkIV3j0Nb/gxZ61lzVn1SmNOtEzSMI26r73pThC7vMup0hTeUC7C5+o
QMH3ToGBWcrm/LnPGMhZgqZFmoqDruitIORHDpa9Bro8Jog5heirNP7pM1deb4T9
cSsbhqUUXxq7649XzSexiJ7pqPEd5NLz6WxY4L9nIGqgTB4OwwKDHaRF8YQkvbbO
4us9alsxadVNxJEvF8wjFZGBBK4oRddGXdXqYWglS0ybmzc9We/eLT+cxm8e7pkg
MZPuldCud5Oza3cRW0g8bUaG5lwZS/Z37kpo1UlnDtKORQyxLtbSTPj0K6cVoObw
LEcNUqC9UG5B3/fUy5/0y5aWhqHEwzm4i9Zb+CKbKyc3dxiM5W0MPmVEbWK0YwFQ
DjgxyBs4od84pKcxX0gvuzW/d24Nf1WaDpLNp5MxKd0kRpQ5BvUnhjcYAEqSns0I
siuxce4ddIafJcErOuIE8jwWq3HApDCjkghs+XCwW6JQZQPbATSCExTis5RxaRFH
sE3UCKNh/badlFXcmQFrL0CwC+Sk3vJItNL5ihoDK+lFoZKIr9KX+kjndAYJ1QSh
drmlzCuVQQQrwfwyVg7pEqRfgx5DpTFNj42Qx2wCfFOKbR/DV5FG++7MwJdV98dc
3cPW4ANo/Jfjt4YDbNP0Hlvtq7n10u6Yb5Z+7ShMyJKKaYC2wlsEAkU62gsxaGQ2
yBe6oziqnnGuCHgX6ZSGVrSmvAh860Ul2N8RIhnjZqWJkYUOqM2Bg1RAFSYb1tL3
Uw7+Bv1IpXCs/SWTRwHBa5BngiKXELSPLxX8vOXyApYtdQJUtkj64CHH7r2P9QGU
u/WLtAKiOHeJLo9lSCBtkKH6t17bV5W2vIvWxdQLT0Grj0XLoeOotU8GM40+62xP
qq+sxS4LscZAhBdieTaY2OU61Pichax1pHQOQELCrSAiLNzj0a7I7G2lJJ6BsOpY
WEi/tKBvD8yUeSp0M4XcU1UwkUNOLySrq31u6VXlNGX0VL1V2Fg4DGpOO739a4Bp
d+aVGiNIqaGh2/Bo5jcRECxoAXYMFcz1WpQ8CVrnKRuy/TtBFY+WZxMn1p0RMBE/
Eo1UjclOvGR4663/AbBR5RRpXMU/pBgARHdnKxFkI58Bf/bHWBlD464tUN4vmx2v
JfKvO9WvlIW+ksMeIoHb35baCWOwJs1V8uw3YmN3ZB/WXVKfPoVPeBGuGZfKV2wl
2B6uAFAkcTOFruiHdVpD68+YGRlfyQDeXK8p5GlPGhXk9nz4tR6bx7X6ZveCZ009
LA+RXtGIhfYIXbV81tEvuytiLAIx5FtWthP+EHgQHl275JEeYKg845Lqm38xwoAu
jLMCuXWngd/PeMbZtgnpIf+gofF7qgaiunyAJKXwrOba1EAdEFKt3GY6YETg9vzU
a2Tbo3Uxu7h2A8RMramdmZee//npHf0/QivPYoX6NGn+aui6QMgyL0eppn0AK2ko
cV+Oxj0TSyFZtB+NdIZd0eSthnIZsfMtGyimaqA2mdSfgE2lfc0dK4RSPZ3pcXQf
qDghIuP6tbeDC+DKrGkliMlwGNzMUtS1MBgs1qXf6h2iT/et8+UmCMzTvcSe1Vlm
CyZyz64iHanY3Muy1oMBIwMhaGWrGKf8QQiYNNBB3hkeJdTkUvTq4vbqpDIejv4M
0jXcC/aZRLkebZL0HEbqT5MVqKkYszZZcQ7WV7pNfAJYBPkaibgtzDKETKq7aQUh
NmRziDd0+eXTz7SUP41oWebZmTqwF09DeCUszbjpkHT1pb+CoPlhRfImJCou2k3w
UmtsUznSfawcfMenwuB0+4SI98hq46Vm0wIQ+F1IWvd3jey+oGN3pXXhZMkqYcWO
HOq3vl8eOMGY045otTAAYJyrtLl41jbwhCr/JAspK/o8Cv6QtopjsZfgv5Cc1K8t
YmJsvkdmazYmt/Xcw5sbdRmAghikxJcfDaHGDJQ3nQXWQaKt97/dxgVfyuhtch88
cT72CcUTgzvvv9UGtjs/1wAEbWIXM7+ePTWR/09Qe6hjKni0XNy9Tya5ksRwe8rl
Gfrnqx2wxwHCtSJwSZH7apAzFnkLIWduAvMN8led9Dn+smSfgf8/wgYlSbz0Fg28
4z38+F+JANBjYw2GNE6SyCur72yai0wFFvzC6EvFQkCOLXGZD2DlYW0dUo0Nu7zw
Q09atl3LBY7wUZ5nrHwNBvOvvR8Ptotu9JYtAwr0w/WWpQCkt2bRwP/p27FILDxF
xj0JWMQkrkp77EIAuAqJMxtFFO4/MHNnidTXqIhudq5KBpab1ltAUloPlKdYXuOZ
g0ZPTltazi0OtlBBfBAiYqALgTRwkJtbsObk109UEFd2ZdoF3y/6ReFh8YNv2Uj2
SfS3ECJeUFQuS0uidRecVgooPwq4Er9ujwabJ182YCUispKCRyI6pVsxby/XC9j+
OVEmfBNVYc38FwvGJDnyOoHPAFiIGSEdHisCt7A7F9qijZ8G/fAgXZyN6tsdX41Y
O0fmFyPA+dDiehcf4/3h4dcne/3ZcHbq78LHFMtpHElcXW8+FSmVfHEd4TAr5moH
8nDglo9z+fK3oBPLs2s741Fw3VXF6UoCF7EBJRBgUVKAQJ/+ipZm1LK2zZteozFq
Go2/huByic1qYTS2IIMpAOn4ARV9aoOai0wPYlfwR+Oj9Bkax7Cz5VH3AEszo7RW
oAnWMrSCHBHXtsoPEHAMc6qxIEJD3vdraGnHZ7z7C/5l4q3sOM5/FfGS72OC0vMm
av7a86c0pks2Pwh6w6YVeVD7o/Pietai7Ar4T8ostvEhdSlFsoEqaEpc/6J7GnrI
lY3vOorLFflx6B3TqAQL8SXrgxE6NHHXFz0XW4M8MQsHiGEKmRj+lH59CxS0pXEA
3oZF/ieag/H+Y3vkD7i8JuOW7JmvaNVAYx4BmP+ersZJsgR7IMciRk22ny4WOnAK
kLZ7s5TCZ85jWTkATF5tNaQUGYV4Lsa4RV1NRINtq9u51YVJHH2qZbZHf6jrVeA8
mI7RVN6msDs9YIZ0ioKMbb7iffAJdmeIzqDENPSVJ5vZ3mZNGKlgLYBP/tK+Gz8J
OSyxZcaRhXl40Jg8ITbZ6wZMkYHQBpOvpzCwNc1VOpABmATgG8uxVs9c3PSgP2ks
oBvjC1Vl9XHVHHLQ7B6cv3dvUizTE5mHVM1hHmQLUO4wOgymW2pYelUtJBHH7M37
bK/xRL3L4eEh+XqxX2Qqo/2HRQialfgMor1U4Khqg7uBiz+MJc2dR3d7DtoRNvIO
ekgLY9DDJ+qrIFH4t2BuukDJZ8Ngxjgb7FwQofywt4m27CyjF9j6UVCcZOVDpZsz
SylkqntAv/WopbcidKTex/8rhJyxjUqr4TMiyadVsRp+Ieo48gTZgKwup+S8XM2W
4hX3FLB9PtLhU/7c1z/lIY4kwbAeRO0oSDb4qgTeruus8Qa5JIX2zAaqXKa7M0L+
rxn4FU2jvMwS/jNlcno4sNSm9Zh59eJglwq70Hv1lZyiUD0CB3/l/ZuMxxDS/MuW
gUhUKiqU1Q6fK8Z4gecUU7UxvciVIONmOrbMvMIc4nVnSANZOB1Xc+UL9H0LV1+K
rc3Nz5hSed9Q1cl8e7gBHuxmS6+1eTLP1AK5LfGfoTA8t3T93fdr6ylaDAfWkKvl
qdkSzwJY+Qd3g73i+pOrWniGPQmiF3TZXcewxEd+i6CmMbiRIxKMRode6cMOnwc6
7kZrSxYdGff2rjY+BJy5DBuW6Ysy1FswqCPSZJgFyqVYjeVn5QR8A1tgdWJrdvDP
hSPlb2lmZlNheWBpMabL7RkGekIAWBvQP8EAnwZO0r64nzvIdyocgZel6BEWS+cp
X6l4YQJAKHwa3xiJH6LbTXjKf+aoOpI09161jup4PAW2NrX8buVI+1WBc6SJWMvi
BshasCD+ymXt4aRfAqsJ8uVJ3AB1MRD79cuEyK/fd/BVayfP/6lr7mTFL+rnYvkF
or+VPiif5JvWXVV8nish344QeVItSVUPTUCD6NTIU+t4EFJE5tljGVyTfFQswVAg
sWaeXSGbTFiXSr70FxHurUzXbJMgaonn56X1+KUb2lJJsNQgRL/3v3ooAOrtAw2K
sEn3D32chl5JAtZIoFCryDKAlMidiJgNbtauWpQUCHEWD4YAFUpT4GE/2/BnJtDf
c1bac9zOCu66loJPIV9sH/+fTcqaKTsx2+1FBgqYbLMnG80YMzli0+DCzeySSZ4f
Ot0m7TpP+zRzGRV9ta4GC83o3PSVqFvdIZAdFzCDoajNEFv9DjcBqbFogxU+2NA/
+jb38lQSbDNJ96TlysWOpw/oGIoPZqD5kFJjVrR9+mABH71w+he+tca+gZPRClet
atuYft14TQjGHBAb9jQGigAR8qMXMyhiVjlJulRiL6tfQm3G6djVJ1ZfgIbQPxB9
PQQyTbg8kqWF28h7m2mW21g2+NkqTrM9u3lIHxMWnDBmI8MlnxK8f+Ad0LcLDftm
TLNEtZDH41qaBhWoiKExZVi9yAvPKfc/wmUdizV9Xv2mY+idYB2IYmrOvM0zWEKf
lrDkj4s09PYC85nI/biJHrMTaNkK5l6wHs0UVFe9KSb7ntM8QJecdrKjV2je1vA6
l7A49enGsU+b45n7gw8NHtuDISxFqsUQaDGoqv7o9Y1cwVvWnyM6BnFLAI61N6aW
9O4Zuyam7ENguMwXscw0vjhTZ+Gz18AsTAPq4Zewpw/HzIqQpDFhvqWL+rVGJU2x
ORe9vgfGU2A2EaqcpT9q5ZMqRl+yBsSfXPqsIOQ+L7O91aDYGO8sg7BKmxJ95pq6
FgYJQU4sWiJLYg8v654e0FP045glph6YqUWphd/NRWv42dK7DlhB2j2u6WgRSSbr
bRSPKcIYNEXxuOXTIycCOICYQCarJIVYDZoPHIDlG6BRfLCa6OV0JfzdZ8H9Wwde
bT3dZPAPR1rA40vrAllXvNpgowea3tCHyK8hwUavLxqlm4Ibpq6gOYqVROhapnGT
C5h2dDYeLS2QHsl0XeWnlt9brgiS8mOu372BSMD/3ldiFceUB7zHPW0GtH3KdEr9
Ay9eHH3FtMHPkh8FIKyrJ0pg/9StICC5SNJWcIa4AhIyC1/lU+uMEzvWDQuChoR2
6z+pmKhoqBtpP99ad52yb4nbb3MBvQUDkF1O2eRVN6yh2NEdiwSdBIRxN8g88Fsr
9vNhnFY5dclJHpYpIVW4Y+nAnzBPBuI41Nnm6wVGtX+a6vYdeKmUv/THPWmlGT7d
G162DYyDw/1d7mn0MtATG0CEPFPx5jy8MDvu2NXDTdfU1YrO7a1XLHTo9/KH++iS
jm9VhTdkkJkgjCgBnZh7SYgBq6/zL8xnFt7hiCZXBClSullOFECPeZI754qCj10C
UpdKDrN8WpbSQr5vZ1vWLeOJ5CFMCQZ5UONtnEJktg63um/7YaLtC7czgKJM5YZM
W0f1CGXL4MtYhFWRZ59+IadfyUNVCCrjJhSDN0207MPkpaZ6aSeLfTKzkztnVoDm
CAyvWm7C1PVmSvbIec0twUe9yhm235eP0vnefIFHBABm532BrBQBlrBBK8ubw82c
+ImmxsA4/vh1w7Uv5KnHHXZ0Zjvjoe7/jTzlA+4kqV5fxVROewClb3qA3KmyxtGW
aibyiGkWXskeDrKUx/NDGI4woFJPJbzmQT3bPCZFvMPIPt+SjNn2wJMDrdR6vE6H
FgnGBx+tfv7qlRNiHgsL+CXQ7FhjExl/G+BljmxpCf9zONf2Q1SzYRk2jpOjNtet
mVGRtn+/xkqAcjrQE/NrrhMEL7MCA6WaTbMUpZJqJPQDCy2A/zNpfyuH+YXwRgiv
KgfXvoTZelD4TE2F65JdUKgNR+7TdzVtGwrgdH0uAZlZBfxV6uw4cRKPu6CKxpHo
xEDsft8n9OuoHerX2KiTvqsJ3AWs42pvMMQkD2fbunWh6LaKQihfGsdHnQZO0qPH
OkduWa9QoRWZGJdYQmWk6D2EnUTEr8PcCkxGqo8vrqqyZnxtHOt39fxahNkmIsk8
+MAAsOA9DgAtpSX0yO/oFDcW4VWGvMD83nwxKttGhkMl7tdwSRFGe/rPFkzI+tgr
bj26FyuDRHniLJJp/meoa5+QyqE+n3WmvdnXDMAChVrEHAtsgbjweFQZ7AJePaLa
yWC0R3TAaTL6pAvgkAhEc4e6a0NlBQmNWxj1xw+J0hf/XXMLcD19QsNKoOvtUBfy
bxNLBj5FPh6aSNABmo3qLiKlg3Vu2cUR+fZeBLrlC+sNxp5ignVjDjxOwYO4dvZ4
w7Of+IqgdQzGzmWM1XF6Tvv0nbwpDPwyfB99UDbNfBXUg3FHupWkLctZj41u9vL/
sLulBuC9qyiEJSHHMRs7WL4OU4mJqjhRaZBsrfcOlYqovbZIrfmvSVSr28zVYrEJ
yLdWtVUllRO4mf8+QPGbgfdWRn3C2CGsL6dYMmi4iA05955Jwdey8eXysIfQGVee
7AB1WkI/HuXlvLdsjpNImuy5yeBd/wPm83BvLVwW6bxgk1cTO0hRr+A+RSPd0a1k
pHECAwZ3Vi1IvRFMfzlnHLiTK9rzIPt4Yi4J9GXlCo7xp6LS1L5OtpI/asToicJe
befuaqNt25P6eO8d9SAo/Xczmz3h31XlpXufBFoh/ioer2bg3/YkJKf/aLcU7i/m
rruGZCmgzJCho5Jmz9KzWJkq6XCu9xHrpyH0ANmhGz50SKS50BXH0phJvyHp7oTj
SHc82Iakm3N3BYycW++MNKj/XRB8yWcwBvjvxXIKe1gC23U8AhVVkQIC90coyxa0
vj157MQi3LUURERG79JXB7gXYM8qs1db81x1MA/hA5LfgtV67OcTpCtY8wpVvDBM
6dEzpbiBbohCg9kZNRcyAMfjC/R8Dp9MVzSVVOpyliumt44ENJjw36EZ3UjY2lHf
GGb6On3kTOOPAO1DVr24wxisM+5IrhXcKhwAcyGwPmCTgGcYxWxiuFPLMHz/Q/H6
h49FLbv3CROhe7mXVWyNdp2T9JCmYdlBmIqEIDpbS5fXk+0fQIZF5fnRz36VNz+T
xHy1K54imMHg73sa0b5emSChtKDnvyFDKyi+KhprhqwTb0B8aprXL7FhdZXMIKQe
i22qPlb834P52om0t+7CzC9z/9lVwK5Eh026aCzjspeEZWbZK+T1eYKpWjly5pT3
yZF1JwaA0CnFTSPiZgXYFr5dtv4OYndqy/2j5vImIHst4cvG+vClVzGyzDURVbgi
y9Mb6IwD7bWaremzD3pQfTkoSybQkLCSior3LbWrfCaD0maR0MgJFN1MjPkykaqc
X6xfqIyoEdDRVormYbgSShm2VdBru5M27WuEbN9i/+jCMIqonkpAxH+gyKNhvJDw
KZHdiLs3frsQ1YiE2oQe/eW8xg8MnNsthtzI30KJYAtU5t1VM/ZlnabPvVwaMHF/
uxwVODOiSomM3+7FU5yYNbhRcybf9H1/ankFLRWspqJcHr3Yk1X8vCwlvjUzXgBj
jSnsgfhLsv4vHkb4V+bivNA7TixBtSTEqrP8MW96TRmoUserKQQjYSvXR/yLPLIb
hw1Nl33igru9k/M6Giy+uIOKyvvltEaNtJUKRmSZsX8p8YSnYo19h5m8sU17x9rA
FK34faMYjjJWmutTu/85uoZ/tDr200chRX1uclCEldJwIHOHqWYCFVMGzQxxIywT
8EdPWyIK6sCZkFXc0Ap9l+BkCTej/UsI3aLJX6Tq+mqhPwjreq6QTVNzwJxZOTpF
x9JChf3XSQRTkKNKLMEWKSJM6YXqk3IhQx99LscbuU2jk+Vw9AutzAngYs18voB/
djJsjO15sccexy3plJ+/vfcw/iP2iBQ1Nb6Fxk0HrXZ/qz+AractrSovOjviKrOG
ieHLD/AaQDlqAYEHp/4GnFh8x6m2c9S36Iz/c36LM9oq/pCHVCao+nXgzziBq0LO
x2oZzUGBiSh/q+kTh0LvRkKhT2cv68DfDuG8iugDRFYdZ3Csx92uXS6X7ww6GOgk
dFRe02ppiTwQ1Oc1eOMLazOdZBYEPRnpq/e6URv+Ob//G3DROy09d6FbOcwk7J98
IUH/c4JBsDSGayTGr2gJqZylMuNTigXyh5wMWWc6B/QS+b0IzVWaFdYEIDwLcvTv
jdTa7V73Ur7tM0GfPTr44CtJsdhLrPr4fYl69RhGzfn0SPQJZKgjBNbOUzDV4/1o
BckpaquHqlhXRXhoJwqHsAHISKj73LSCQ1uWo7RDCUwdLbcJ4GqHY4HycCoUBq5a
Ypwj+bMEdvtWmmiznVMjthSQs/zncqNmq5+sQYqXbYZH9pzZK8sJ0taonSQ4grlq
cqFn9XpLOCtOX/J/8fLI4pKfnP4KqTZpWofS14tkvi6nKZ0SOUlw0knjqShtist9
OhwhKf0JDOiUKZKGDhLevirnA8cadvOyAmrGgNmAXq6OzKarSttkUgaGp1O3XVEa
NnxaOLe4gRyocLDGSi+XkOw0XvJmBgCchScSHUW6zwBl45VthX51uEbAyXcxfcak
2qxhTQMQZjlVOb2yheCoMh/xOjBb3X5dJlFLpvxOPmP1kCzM5jgA0KGiGyBab2uf
nasNAwiR3xsRI369QlfBiz6ZO4loZncljIlPuE8h37VmDtBRjtDT9YfuxSY8VVU1
0ts4C6uOL+JqxhUS5AE3bridl08+q711WsHcJAHNrF0QvUIl8lEVlyUo1e/usMGJ
ecuvbOUTuIUVsl33RAAXtxxErgMpQe5AoHOOKEbW1sIhQA7I72ldvMZRf1yocxg/
tNAEtYhhexWwZAr7iMVD/z82JbE5xo8JhFhpsraI1z2IXOpd/a44wkZ6JBEJMQJq
DKrNdY8sws2p6LndHcrQWHbwes862BoKwEn48PcIETIWmGRmzDpOT6ZSUo5ub25K
cToQAEFOZSIzai7sen+d3UWkxLeWqtTo3Xxd560qnWAoKNaJfRg6bfRAfuCd9Jrx
Q5lNdYLntCujfaAXNC/z4PRFrBVMgmXDOMpH9LdSZHtzj+8JT/D4zftCmvcUHG2l
xHmx4ib0A89AMJLrmEATE5E1VofhwK9tgk6rl5F3GUd1qlNHwJVYrVC+XVXvIg5g
Bev8wtx3esdRYdGF2ZS6x6IseQm1qzGmb+tFI/CaZgsDO2Jgw7T8S5EOPMvsPThL
wCRJbpM3a4UT7Bjj5hRsEJFy5uJA3CqlLZBlKjZ1Q9eaWlsXOXrUZBx1/2Puz63J
+ooYYk+EhjP38P+j4hGwDLF4r6dquVev37KJQlqKRYmYXk5yQPcRbRLcBTjBzjiO
N5z1ETeWqzx8/RZvsW86ansGfCCAnaAyF8h3eu5RdEwWz/c7SL2MLHY3fv+ZL14M
6au1pOKHKz7PDIr31wwdLUlOIMAlJTw8z4agVmRhSmbegcKkVNM+MCCJKpwaPqvP
BSMf15tB4nGtgLixSUXqw+r4yptZkVObEHzGDWWoi3aKisS0vbh9gOHBVL6jbzlD
hHSUkzGDYFNOQu+lF1UiFcsjWGGS+BtGtDf3HkwNigSPHKrXqJfV9kqDDor9geRS
BijRyRgZWEEXP4/ZhT0LWCahepF+z1a+lsaAqM19DzK4by4cjZL1yebHpK4LWcSq
JHR1+ZqgwbzcvTEWOCWxNr2mhdEwQT7Hum1RGFHtuY5qfAIfHLkI2dgsCpdmeyVD
MapGq0zovUpn2iTCYp0j4T+jYlyeE755wt489GQ7vEUzl9Tsz4w6NQhdfn6PKJno
OXeqyxsF0SIbcmvliFLrxeuSfzmhzpTCbP7ihFdTsPHcZI+A/FVCIYNOrxTVefXe
6Sqn9gKGBG+QU+A6xcyZni//omA392UwAhvHO9/hu2LjgOnVwvABXU5Ye2ivGNlN
FkUdHmlgMen364c0VKJuy9Q2GzjbdVFHSxbTszBD8OlSu3Y5AE8aNNniHnR8Vepq
T6pL1hAvMpIEYG5Bi5oQZyxUWv6fzmdo2dtPa9LMW/ZHGsWPYjaC5FgPI9Q3mcgU
AL4QmSatGm9Q5NcV3sxtUjys7cIyoaNoMd0F5Q9+UKyx49kt0JuJtJB5fwwV1V7M
MnNURz3iz7kubjt6ji3nC2+2Uu5m/U8WRexIVOe3WAoEieCeJC3h63WOCc2gwgch
wUW9zEZ8dFjOr7YU4uoNLjSvi99uyPN5HW27J5C+h47ER/9repo4MqgDy0XYdd+d
IxOz2SLUVKm/8hFwbUY3UOUUbzqchFc4ycDwjmWz+MUtb/nRdbF2gcA3YLmlVEqZ
e2CZCzwTDI+0P4qf7YTH+Com94EEcewTDi3T7RKKRjhgy1t5Rg0/CQGLpWpGUqt3
TEdqemd4P0385Tl2h2EX+TGLSk1Zi0fBbgk8GSK0Zytgpny8oi/WU8ZiRwDOPPKW
hDFikC0hseQnYu3nTbADrWXfXuy/egyjN8hJMaQB5irTWGCUzOHYj5XjoDnhkGKM
gaFKzFt6T1JbjHe4WZWnjY1H4jtEj+I3SUU6pILYSesl2pz5lNB7fcE0V71tGpyk
nnfTtHEKOqgddr20bXLDDiK7epl53kxjg2tyw8Pu8cqAQEtwPcKRSSrHnH59XkRV
y5geU0w5vlfbpG9AbEQ78uVXOtzE7+1K+J9jcxCfPayHu7DyHpqqv1ZeMS6XkheG
4eYgp0C3i8/wLqPZzUsDsNrsTqJfTUBMR5NFVd3jKG/D+7n1m77Lvoh7g5qG1cck
r2G6LWTwuPHRneN3iaRntIt7rksPvqcJ1OYdwPy8a+y/xTspT/YJ6lEpLKWAmmOP
mEjOwuqNS9EaH3zr0nilMKuDo2XX5brBtPn4U5MGGx56sEG6Ca8ACxVb9z3ElJsf
IDRf8x4n2CvLlMrlNiaKqWsTNgA/FsdJ63CiIIHW5qZ8Sg4bo3gXysq2ZX1KdT/e
xQLuh3f9hNwfpaMwwZoGXDgpbgxxozlCc73q8Lrt4VLfMYenlw98x5VWhGRUvvym
mANmrzt17GN+F09NVtv+B5BwiKxtNhOiAFx10KNLDFJYd1b73HTFyONec7fi1+k5
n8eC54QO+cyNfdtChR2boIktqq/k7f7ZMtlxpFy/S4crrYBfk6MtJg+o4k8SDT86
71B/DOoZIDPgY/afM3DR77zCSnGgOVVyjJjiHDwm01TMGI7ZgyvfarWiu7SW7KVa
OdAIfBBxJH7Frtak7Wo+BOcHh3FlHERRDEzrO/ptVsKkWqsU1I7WKCfdrEU5iOuX
4xeK6smVwuQd7N8/OamjuHHztRqAo2hZgon/VJYRJm6OTxm4zlPtydsq3I5iyata
tLy17DSbraZ+mbrVHG2PRWoymsI8rdXhkNYCbt0a8WzmjXNTup4wr8fl/SWmLu7B
4wrqk7G1tK2SWVbDujmow8VSbIVmAuisl3Y4/N9qr0F+WKe/95iNFfIhMnuE/hko
7LcutxXqShKzEMyt8T/Es9v3kdDrQ1HQB5EmDat1Mf8e/mjd2PdgHs0nlsgpUiPw
PoCG8U9Ga5GG/fNyKIus1iBCdUVCSrNwdtBrtjxaJ+NRhWMrtw/iPhsHxduB7wGR
RU5CcDnFJ5YXRBQNFla1Nql3sN0eH02DsftZXHie2O2N7MZd0fvaUi9EWYSD2tin
0O8CrK/6M4KgEJ8oyuQ0Gv3XFT8n2bKtbIwjb+f3g+nqcYh1D5jKGer8aV0balzm
g8NJDrFbe3+Nd/SGm6AdJs8SV/m2CU+NzaiFUOhiLdYGMIB/aood2xEpTj7ic/SO
/14DpjhOgFYwsQS2GPA2DY6lijrOrr5/LqcqDsENmXGE/BbEm5QWIqil7yQrU5yE
N16muVDvVxTQRrK3hHD8jj7KK2wbVu7v1NHTOOyROgI8Ou/KrVCCogE/rJMsNZB3
i6Nm28hHiW9Svnkv7KEPvmi72RWHl2Alk4j+BCAw/bKkIXoYbQ/m1oJahh2szE1U
LKQxNNZ/lpUqfM+H5kZXle1cCI3EFXJPNEZFaELyyZL4KBpruQaW6kZm5hjlsvHi
Xl42EaQwjqHXTrw3KbiCd6gwDc5Qjpsn9YU2OeKQE/xczj0SZvhNRp1glrCKCtca
3M8YGSZS2zNRcjRsJd/j0xWf5eHs37e+0NW7iwUG52bZZIDflgZRDyjky+jbfWz9
8wTglxNqD9iaXTqcDD+s4ueIl0TsmXMc3UoL7Ko44nICpDWbBmJzva5dSQNvL9uC
CJYwtFT30ibolEEijQwYj7eHe6tN3ZNPG9SniKa+nSka7ZqjpXYdeYBLfQaLk6cs
D8NjnTBuVBxZV224fS+sSKM3s2TrI8CUDz66lmqufiibHirCKYP3t++mseeM8pQc
fJg8aTrRzUrGEG3oG5JGZny0gCBT5rG2D2FEt4x4li+D7rGD84euBa8kZ0P3arwz
oW6J5N9wc4CIJxmwOqe0bb8UAqsXXKvsXioapfqOFcNCZnkj99RsIRy2izfmthS4
4K15K3Qco7M2k3HIqLEriic7YMthmLAC7gEmbGLYqDO4YsH/W1+iSbJ6ZmFTDUMy
XgTXPab/hikCyiNhRHAB9UrxRvqYZEtagPdIz/SqjhwxzfEjnrgZJjNWsbO6TrCB
1kF/8TtMrLFDiJ8ZaKBk7F/aNZuUIM30oJhExJkQ7BVXcoHhxx+ifiMydpj9OfTD
ogSJyxJVWT3vOzuc63KeTR0HDdJhI2y4mCtB7GzOlJztATr+pdE/NJUQzH/bTMRw
I7dK4iUz4nWLubzhn/XWKUcbpx0kzglHM36zZ0p9OHYMfX7W/SqBWDgVocqn1pRj
/PbX/MTlFv3a4SV8PJhj4du7J2S8jndk8uX/LaqfG83D9MoOiSeC/fynEFR65v5E
85Js6v3fHhGYZCvw8rQy5SrGR9uUdsBBamwT4watuJISvqZ9cp9AfNwRRq4R2MT2
y6lIN5OA1faDxOBQ62VnzrmnMKuyTDft1Js4MIPpEfDQKQ3zeR8Q9oImnCviPZJR
G7+cXh+abkIFLaMUEFSFnK9zh0TeTHWx0hXwT3R6+9/tCEB/6H/Io3V7bxBp0zDR
ym8ZjLTE/kM3OZr3M7xE51x6OTHpRfB6i4KziRSOCODnsmP8CWEY6pnxkws9vhAs
YqeZQyq26tQAXTm0xggLonHbZxF/lNxi1OZm60uGfaRGHr05lhUN6RgfO344NrHv
4cwbWQYKDrFGN5C5rM2shdOhRyx1ekyK4bvyiRQZD07H9gUG5wPROTBLJpplPWQT
18jj4/rancXcu31HyjmyDHAmVprcFiK/PYz9La3a9o2N+AacTBJ6UKvOlAoT/UZh
sP+nBfktD1P5C0oCglrN5Aj18aiopxPpRIgLhfTmB9ZFtTfXPktm/xOgcZWUjRk4
EVCeaLZZQkLSOx3IlsDRiQ8CJKZTiaP/gxEODoNczW++Byd75tvjX7xhhl+rvI9z
unDnDN7b2Wu0tb2itgKn8KAfUU3+sWm0Bn4tA98SicJHcS6VpOy3z8cyrx+bfBh5
biNU7fowFUku2qC/wEf83TlAoB6yXZ0YVV8IHiuTlFO9vfbN6kHjuJ669n1AVaZy
ZRgzTKOBBSJUnJthUqBTNebIRompltPjuAXztfuFnaBt9LXMWPESbiWRuEowK1EX
iZtIavV5NtK1EaG/rWQzVHL3xlwQ7X1hp95ISCOFbTYeFjvcz17HfOj8+aWW4NkA
q671C1rtMTSAUvZ6OdCQ9+2n9ZH1RKOu9MZHvbgXhQOi8ZwtgPDT7hxxX20i8FiE
9A4l66Sc7DvDUbdSvBCokUmC4AiTJBN1Xj3v5SDx/WaBM+gyR4Z28l8GZFB8Wb0x
ebslCEBfLU67YtfWncIhjUK8rkwCUDu6mVYJdwsUc+EV/bQu52bkrDZF+vUAou7y
Wg5s7hw355IISLl0tx1Fe83eq4al3Sy6sLyxJjU0uDw8+dTsHK852l9zzttLLSgm
MMh5ckV+R6JUSX4QtqE//wpT7WJhCToek4R1hr2BAT38a9VUF0ISP/FQiqBivqtR
fzltLbaQgM5MgSgFiVxmvTGGzSzHq8EFnHiI1+hQohlFGYVXwMx9W/1wYsAav7Zo
X4SI6Gx1vEdYRmtouudozLT2wTVNNzFvJIZ6tDUQHNRzeqr0wTAZwV7H+6hlkaUN
iEJAT5RAmFJO4SqghsKdyX7zgfnK15ltn/seGm1mlKZya3gb21LzMnhxGnSfcYg9
xXs6yyCUV6+V8mWtpXfeTFrCsEeN63hrx8dX4F2Wuwf7JpzX6egiISs4dhaBExU9
PO9TRLCxDMdDuyadsyaZkfPv1Zbja7+WsmU2yq+vj8bWwK5V1Hh5D0LJ/T2qm6Oj
6YxP0YAYGxS0SGaxfZ3VzpSydwjWiJJTIiQJeQxTsIdt9dbYzvLQi8FH9tgRMVR5
p5bXaKrdH/Y6P2hIYZRvjL+uEkbefpIsDSkXSNaFERqYFQRXpxUxtZqRqQb2SuBX
ZwpwAsgVurhsRqScoU/QSi49z4KMVtk4icG7Aer3mk3HQISV704dkGdTKY7/FeL0
eAilXaKNTVaB2PLBWqjtNxwPJl29dErry8+Zdk3sdIya5U0fPRA9DoZSKNkn6LdI
+/T+4jWamkqO7PxBbAPbtTVEpu/gJ7LwrYgJM6lIQnplQSFt256eeBejV9W85lhF
DgzIyVIsdps5ifNNE8xvQqy7+IqcKXsU9lYuk/6XGsvwrPvv+948h4JTSiUSmCGC
fslX8drL+welCZi2voIfqEPWn+fibpNIxla9A3PddihFB+FDAKEuK2PQJMKvBI+j
j8ffo9/n8sgCMbfAxd8fJM9PdTvX0/zwxNUa7jRZuV9+RB8d2na3RlSkhSvDkxgh
vfLtuAWBAcYMnOgWQ+pkbg1ymf9bG9NGHnMDUs3FJi9sLMJY0SL6Ntg55nHh0nuq
1tOEC8TnR0IOJQFpY9jz7pGRBvU3qVGVsDQna5ondDAls/hHKhQnEDRbAr4xoXMl
PThm95IvAW23sMhl7U9o7W3FPuEfJl5W4IvxYsCvOK5Lwaqi5uWR6R/j3ePmtUwh
0e5l/AhmWxkqnksLP2MI6atjwEZwP4NVHB+7J6/V4ziROEMKT6hqW8Qy8YPjzqUA
OHyD0H85klNxURzRrHOQMHMpkfXiLj0Xd8LpBpa8tpldOnjv17sz6qzPdYIT/1F9
eSPrfPNcJyHh2iUUKbna0WuOVE/ERpYDjNYKMqgqb1Mahz+HKKRmA1Y5ATexAWih
OKk6o0gT5YwcE6BCM7J8wz8bNFSZhijjreYh5Ueh7vUybHu2zsMo5OdRhKg0JTnQ
5EMloMdhDITLF8CbtUs886NtzRpPMjFkn/6XHtzXEErWvUG2Jn0WrrvbIi6klDXm
nAI6J8zgFAvjrZwhJCBwsI2jYOj6EFVkE5QYJuRvToOW+1uOGBHAJDLyeYh5frK2
3qEB9Ck7k+AwX8/W7pF2YezBgeEWcZWaeQTVRGbDi+cKdsPai+jeW2rGJT0x1wEn
07eeObXQfTFw07opIfswhMMsTMwtRtBOEqDiY6XbH+IFV5uqci1nn4lLwAY8p/Po
YqOpkqZ1KRp/2kcKjVNrZHGmpCJEC9eegKpNWGIQ4CdGcW5kBw9+jxyXArZ0AXmh
3ZTqtiobH1oi0gekXx+Rv1M1NiqDDSnUU58uKcuasKkqv5tLle7BgtdzBKiiKxEu
u70DXu5rjJBQus4IFt+jGDKo8ClBRZyAvNX5daRZVTpKb9a9JfLU4Jm5m7B0Mllo
SX8SCtc77RyrS/JUsSg1WLGBjSXLApy8mE3mEcvWIHRtKgrYWgZc1MsctNLiZhSG
SOzXKWG34ZBsv67KiTBSaciB9btmNVEbGYAKRrSiTMtNjT9aL4rtPHLrzw+BhVP+
NNkQxUWbzFpWUClMmkSeVQRuf2pcWJhV4mTl73OsUbEFasfV8C3SP5S9KIgZbTvm
Hw574DiQv0iYsdw2yKrbu5Skg5o5LbPeZ3AKLx0CzJihBbPP+XqHb9UHqrCl0bqg
GXrRxK0YaCcgmJZ81otFdaIB3SJuKiVVft9l4jry7yvTj4LT6LQEBRTbjghYsGEo
FEo6ksZZxlQsl3M0514fG5R9etkTs1rfDcX9puJ7C7Sn8B9jojCPf0SqaXgjqQmG
ooUpD/lf9gS0XxJKt0btxREUmVedhWXneGxKqvFwyvESMT/tI+Wb2zAAW8DsHgHU
9/AA+f6BRFGOAteK1MzvA5lj6PrZayY7v6XyqQ87VA06cJgdQ4w0wAW0rUpwJr8a
LKy/uHU6hRw1gaH558KEWDmPu10fhxk/k7WwnPTIDrbX2U3i2bmlWAfMZ87yvgQe
hG61ORvY/1GzHwQ1Wu4h6jUDgRdUhRacicnkmbQlZYh+Mr5H6AaLRBU2xe/ND4Tp
xHNJK2ffAo3RyZRlplhr4zLuBwdVYIJMAiT1rnvt1i9xu/S3BIXfy3qP2/kqe6Rg
nEW5bfjIcANybdOeUDBdpcuLO+k4TGsN+7KLlEKiE/jjrhFMe/x1aqTd4mPgzEr7
wDPz+mv4cOGpKXcdbmXxCKZAHkUP5L8802PKpftJwkZEUWrRNojRpyWsgQHHPO3Z
KxqrjA4EH0QsGuh1bGmQR3gwoBJfLIuosnA5w95GZSG5QTnvNKaSg1PUXiJjRrIU
s3Z2NlbZ2BEy7ut3/Tj4ZFd2IRDthi6qBbR27P/UelV68Gtg+XMHV7Yoce1tuO8a
ef4kVgRCWxoa7kJOYwx3OD/opZYzMD5hA+Tuf2WIrrL/Jbm5OG3CasVaxhEIQ6AV
HI6EyPi1TkBPKr6ZP/lmMNvGyAMQwljnni91UIRQ1DjeJx9/ubpBkcWPknmfAav+
7E7Y8BOQRasVJXKrWXnSOGvgkfvF9VKjrcp4/XsIJezvoUli7Xcy2gCdv28ockAd
/ZIJTsCEufBCvcyXOFtuamO2L3qABKUsK275+4utHwZ3mNaT98wQ1eWYnBENPonY
UFq6PqMSlKFXxGZxyD9n35otx6OriFaSBDOeyaaQTP83Ng5F44av+NvPE2PnaLA2
W1p0H5lCGLmvroacRHT5AW7vckkPMyu3eOk6BSak65zgyGmJdgX5LRZzeteR/erW
09sNYMuGd+mZYrGp5XiqvtmQDpmxXgD5/W87X3xje+K2WF0MnXS5FLxqiEUazdQT
pPSc8lup77nhatyTiRvM8Kvv/JO97GhBodf04ytfJsLUijEnveJhIZfUlK8/lrRO
HeCiSTBBJkKyHtfTCmh6SojlE0GJhLRs1Ffn9v9DEi8FFvEYabVdZZcnAjImQYSt
5/kSArYb+aiag4kgFEkualVQO81/kOighkXjxACrFWHXa+/hV29sZAi6+hAhHQQU
t33JQ/WBlX+sdb32SwHO/wHlTfayLfKKIraHbuFzHNRZWlui59JNbgZ10RC+s1sK
z6qCV+t1AWWA30/bKHD0uUhecscFOXXOmQE/Pb40Crv+G1sLcOkMEy6G0hpZrloV
4Q4yczic6LFhqDdcfEd199dOOXrca0Q8l8UzWRFyOq8P8RYbkEdEzKgX8RszdorW
UgXCJl0T1UB6FYFtr5dq+o/iwCNsYAiydFMXK8DCmaUSvmK/zYh5WvaUOEPsRHnt
n8CxvXEwwLv1Wd7vBYVeHxU6FBVSX90E62q7GoqDUtce3ragN4iZDiK4whRbZLWR
VZScs83jbAdT+hFCkF4RrtkXH6I+3HULxkeAkGQKRNMFQlmD7qWPLFpbjecjo8uL
EI7hV58kEw10TNiXTvxWRt9F0hfopIisEHmWMgbvCmF4Emu2ibDfaHGKL6o5j7oJ
4nkuzQowUQOKLd/ybWepc63iG/GskeDPMQfy+pBrha+5UWT/H/DfMqNb25oOsgc0
F9BF8+LRQKlbFHJma9CchrnhQP4wQVELYxriCBRxSaQXHaSpJ26VEe9G/xKf4+0r
37118wWEQ1oOVpRU/NkmN3cFqUaJYutzy1anyjaGNOsaRtCVxNF1yU5UDfIKrWbr
hFqwublSSSyTn5Ru7vq6jwseIY7gJwNh4zpTbgUbhWiIPJncOFd2oUTBpfgERLrI
J90KFs48PIMF9CNnkqyMVVkPAYtNvFQMwkn1KthTY/ELAeazp+R/XHpTRwQXZobu
/Or4INzCYw/CoU2S0Yrd7Lzy5/XaVtbJcrd4Idod8KEWWtgR5kFQWb5Mfl46du+D
5j5o4wXiATGRtwSrfpXQ5mkmlJawwxCsob3AhflTCBt9f+XJRoxZlxvoo7PEf6Jw
gY/oB5GCz5mAukY55dhUTaXko1cT8V6Ix6J+cINWCUyA6JtVk7i48GfniI74RBL9
zenUStfRzJqqmVWm+AVRKx0rutXcXrSk1kF5rfK7FmnuQOXSKvIz32gJYB939Hbu
JOwZAAHr2BOmKEVLtJVcnya5aCERDiAVL5ZW7/1BVNAkQtZmkqJ2t5E9U84aQVwh
318fyrTnskHH0dkfel8yFABRVyFLf/fqBU+gDVcovuibgLNaQ2dlDLeoL0XzOCzU
72IlHahwaPQs8hC+MhCqm7o3SPQQQbkV7/0Am0KsyiphK26DZ6rZsKkYURdw01Pv
P3JufWyhPSEtsJV5obdLOSf6vJv/HzHLHAVc+kwrAd4wQ1otbHQfdjXyCttqaCcT
1oIt91i2f2MDYBsUFtRSI8El4fIHDGzP6OdQy+aDStuW0Hue+bwShb02bDCS1KIN
f/v6B+Cdt7be79RSskPYCoN9apJ/Y56u9f1t0Ns8ca87P4kYXY2BwUhF7sxHAZxa
HWpozOelOz5UJuaRT1/pto1O4vGbzWN9LDrpYXLs6h57AauSSrOlnROQ/nwD7Jom
9BiBwUNAmZzmHCBfn6/Icnhn5o0VJ3yp38gXKNOrI4MKNwJg082fCoqliJrsVD5o
QrY1mF7HbiNkGMRBeHqXKV49P21Joc21o1ogk1VrvnnVE5CuexBAB9NwsHzSDF9d
WsJnCwVqHSEzvlDLWP3byI2It5Yxx50boXmTkzQJtvMX+LLTQM/qfGYu7iEelIB3
fNXgHwQZZ8h+9zLdw6euEMdDKsunJnljAej2oPAEkRWvIUFz5Dz5FnUFf4JeHsZw
TO2hj2b3HIvSPODuZmAZHLeSIIUhbNoQdny2FztaNqr8FjBapH+tLmilU+I/bRdd
7PdMDUVVy+52Nqf0tUu8SDeypzfI2THExcOgNDhXfzmFsnSJihXE8ZZkCYGSGfp3
FS6qE8LBmPvfJESp8nt1qweCdNnDIrRUYKmOgyWwf8Qp2qaDuF16P68Fh8Ir02HH
4B3/KRP5QvWyj9xwVONZ6HkU0mpmoUg+SMgbO5VRQRLb3FQRlHRz1OSuhUGahVRM
zWhTzvA77NxSn97D4/E3s05zG2T+uqUlhoTdv+o0SgsrTRQMxqBGUllWSN0z7nWz
8VH0a2E6Jl43vBvMmiF8mBWP5J2uiWDN95a4M4L1ePPpdgoExb37KD80w6gs/dGX
3fQ2ysAMNq0PeiQoPlBdW7Qm73553LKnzMg9CSmmCE15xFIAp2UoGCmJNstb8rDZ
bnnFoP24t1ZA7cBVDRHSwfiDdnT4ZSnJkmWD2SbN5RZHWSmIXDrCM4Oqsu/yGJ8t
WALdYuFWlnwgkl5gTJo39Rx2tCBhVgsUY2lJTWoBNfgF4zwMjiNrlB/4+9h9jDi0
kgcYLKxLbbNjdKqB+RWoErBYp6/m+blnOtjSvCwAzp4xriOtg3EP5paZ4WkFeOiE
92eSSdc591cn0aYhJ1SA09tCNx+oayKp4/Jx8uTZoEqhM71tf7i6QCcfbTE4efq9
Wje+HruP39dAod17K6czucBj0blhI2XXafW2AeHe/Wz2N6yYZSN66TOYVpZT3f1r
aW+7SdLZT5983ho2dx4t3XzlAU8eeeulV78d4DeaKnsXGD9yoG4YUcR2Vt43CdvR
xTOacC6pYkom7TG28KHl4JnOpYHBGVt6g98HIc4l1vTqMcOU3wFMwtxO/uYt8Ij6
wuRG3XP0YebtzEm6TIf0dyZVlOaFq4whp8zgwAm3glMMX7d3ntC/pYbLCTufWM3L
MgYjnSp1OCgTKU/5BO1/vBuSuoZHzC9P748rFoAMGzNifzAkDboC65RMt/jaHEpX
GvtFPR8XxdsLB28SV3f7ryGWtx3ULcnOVOLnTS+JB3ZE9b+bSw5/xyMXpJX/dvHb
N0WcM8V72OwmNSZJhu61vGlqBnqj7RXQIvTeUSJkGdsVcNg+v9gysOXJhFrc5/Fj
PTZQc73OklegHXXS5EBCVEQIzDlC6YLA5eGRy6YlH2wj/VVyf6/pGHpzfdbNw+S7
OM/hFJATjqrxBrGPlEB01fGLx/qfOho9HMv6q9tzK6iRe01B0QJwVFkfU1jwuTs5
PuGAVLUT8g7osSvhpR3T/H55MItp6L6wds7xMAlcI/l3a1aVBkC7RvIoV5YoNb9u
1g9KpE6tYrFZKQp3sWXwwFa35V+zBl6Hs9dTGU3XyTfC6zAGM8D56P32iQXawykK
GESrnmpboMrejixkzO359qskXYQ0Q2bsDjgXVDaeSSZgKmSNDNSt0fDe7RJTsTbO
nX2L0to1N0PrpZubCEq9+dJlXxP8JL/Z50hpl4/EDlcuUDjarc5rdsvoXRKZ77zf
2teNdefN/ul3ivLKZtSJ4o33AZ4bZp7ya+UU9DW6fp6LlEX7ZSYR7byZ4vw2N6fM
yI7AZKVBRR7tR3JHDtymjAvcA8nYl2U13Ov6GGkXGcY55O+eqaWVOL+qLMIV0EoI
ttvRNqhTv5ARaaDh6wW6RTCjdy9ea8sbVe3P6TZA1SmmjVsR3hEsg5KqWOoOi2V3
SVyzSU8dnxgp2PAwUOJ2F/FxpttWURXtuqN8SJX+jBq/SOArQCTTKbRitj1klcX5
xklCCIKLHq81me6iqriSdBKmRh4xT1XdXDSw+u8VB64DXp+v8O+GLCK6XJhr3/P7
x8iTu06gmV7tk5yerdWeJa2SJ/SeH/RcezFD3tihgahg599vUx8yOt8eTnHzdVGd
Zjpl9Ozgv0tEOXGbxYI2B4l0EEXzDYSYwpin6PPq8aemEBEV4/X8vXB9AS3RIE2L
ddMFXL1vt/vBSiu7YIIR7PzgWejtUrntz22HqcdeaealA9oxEwseWJg2FojVzUD/
MGt8AzRL7udCh/x/UwICK6Zr0EFzbSIdp9Dbom3PtO4XB57VfxMengBsGKv+2vV3
cc5aIhO3MlYH6AAlvXvf7EvJvAERwuH3xIVtxdWKW0kxFgTsvAbSiZhZ36k9zC+9
4ky00R6Fjy7Zg8x1J9Plh8CgOISSwK2HfSVGMgMuQV5FNsKXaMJwifVOMXo8rTDo
jsoOBALPxr1ZnkwVpMwJy1CQowloE0GvyVCLS/+cTvatijhqf+nCT9AXNZtyXOtN
0iRIfkVzhFgvYqJVea7XCgV+x3xYzPuXsrAaBw35sI/JDwgDG/FKncigpzuoKEgz
Sbv36rfzOCvprrOjorEsQmyqc6sanwv9c1GBrJyY2LHkYyXdjOWRGG00r+8z6WLc
xpq8RLMIoSbCpSgJHIbzuCsEHO59Xnh5PMiOfwrYPJtWZADsro/MP9B/UgOlJoLF
2IiU0qvQ9aph4AdQpOpQxbxNO580YbuO158A3bjy7G+vdsWc9rEEO4OG0pgV3+aj
kWdN9E6Jh8jj4b6moiaDBbOesCqI9xWb2XY+/N8/RPW0ZKVjNWs63nkvi9d+x0xl
FJpTy0oT+zRRXquJw0+1DDBO4CrsMTm1Ymb/DINLDoyUClCjH3ojwau5+N/stdXW
jRPG/0/mKXRlM2QUExoMfd53114ANtPZ2bhaCBIIZG0u3hFzMtqI+eSUM7UHIDOH
y9Y8iJwPk5KqkYVhbkNzKTngjxT1MvkP/P/XjfhzCc4HlEkFGZ5+oO6i1xRCBHAk
WTAFnK75PeIZrfUDj97rQIXWPnio5+B605PEwGXaWhzHDNom5alwjYXnMxv4jbOa
ykDMgzpcFI2MipUT32v4FXV1D39ptywWOQN0O0ML7rMST7Co/khmvrH/K7BvEtCh
WkLHPYoRZtTvobbD4JAkalQr4p5/0HRiMDmRNvoUm65Gba8de8Rg3AT1RBfT7Kfq
cGYfj15rHKXE41r8BPm6wzCm2M4k05OWV8Mb2KfLjJryWB+BbyEE+155juqO+K9R
eryxaCgZiPiR5oiitttyJ2tupul+wHrN0QKOuYMfhd2AbLD+klgUgE+uB8uj2sYx
mg0yyCFRO1Rju7vV0xevV09w1diDio7bnLvokbRXfQJ24XS6zr4tDmMFajUR7ad0
dQMcdS9/ygNSDLw0ysOHWkSahFW1UX9gxZhrsJ7Ae7q7v6e0LKhjW4wE0K1/ZnS7
fGXWxWpZsc2O0FEs0OrqselRwL5aBFIg6RX0F4Xp/9u9O7UFNUqX03fmf+du2JcW
SOyjYdrZ5g6DfJM2A7p9ZaUSizx6jY/haf+0o17Vk7qA5pHK1GKtlzSVGOq7OjOu
+9EyPVFcMkrOmGs2sRuKBFmBR05nnp4sA7S8JbQlboLDtgh/f81pGpHELS2HYu50
pcuw37Kgw2IETabmfSQAgihAS00+NjFGYn6Z1lySqvAL+5drRVFb3okyORjWRjo9
XKcg2ehsc1KJrqEQQwlB0bDWHoM6OzTx/+RsplF1t7KWSKKvqG9ZVE4E2E+0FN1g
a5fWW4nyvcEv/D/WbMDo2durppKuDRmbxS3Tg2EADxkV/jfG+jVqGK0sTccRz05S
8FES+2yvXLXAsGm1jsXLj+GqWZEdeVkyGf0XqYNuTBUGqT6rnlfm++sAkA+RW9W4
RxBsRnZ2iHqGudOU3zg0dsBfRwlGv7MAOKujJK4OSmyjm5BBcnnOZPGKJsdWA9Z5
QRnTQXxVBS7vH2etR2WWhiS8aSP/dVZBTqYasWpUGTRA992uBcjVWVnp7sWg4yqv
SCHVj3GGC5zjwRoH1110mt7g7HF0Qh04RLY4peD3IX/4A/TsGZ57fNTtDU9pvOPM
ZbI7PHnxTWwHJFvRIlVwMoamXLYlNyJNmxLtIS7ko4steCwS6DDiYb7dw1dZTMX+
4US8bfhEp9uJFwu1WU5U/59kiuN4V2JzQMRNrR0mJY2RlPRRtT6Kb3usEZ7+HFY0
0RtrCr6jkrbWsnKa2zbJo1eU/GPwwu3oz5HB3cGKF1Tt8/6yNp+IDGtFqiyT65Bv
U5fboIDWBiTMemU5GkI/ms1QUfcTnocGvBL/Q+TLJxHnt4tnNYWhDL4AzWuJ2yxg
eqyL/Z/t7XVoVL/a07KMIXTTKoXGDCp7NEIjsCCPjykJI3E/vTJ6oRvsooqrTe2T
OU8Yw1hS80WisY2OFB4EmVucOdMzuuNeyak/K45a71hRUdgTWZpufziTN7UyRnHy
RkzGSykHR8fuOCmUrEUxjvu0zG4JtpYTMcZqS7u9wBzev3DcO3ABnpNntmkkabCJ
RgpQ7dMlPFOzezRNyhnt9U+5p7xIZjW1grqk5f//w4K5n9+rccTcNEdLXRYeZRZ7
zhUXh+va6Mrlx3MMp/69TbznXSTse/TliT21wVchkIVubLkM1eNxTzHX2CEFUUEW
qVwWxx5CRDOAVsjQRWCM5F2lB3jAUGduyqV+qCASkbKJoFmK3zrHY7da0rTg8dre
IwOtB6EE95pdlLglNjhVJNcD25GhSM/GdkEkGU3Ku3me1z9DwsljK+fMmqIckqv4
OPSoozfzp8MXfm6ubas9RSDRPQR0l90lGoK3mpxbZzRo+cUDsQS/6yt0luU95xWc
ktEAoPHZk94zrzXH9bEhz7kqrXkcWDuDOzIzLVTdPWAEQA5oJNG/hiTgiM7TqqkQ
QRfu/1zsthxqBhwFPJp7l28jYGZ03iy5j1NYrtArnqwmPn9kDEgApX9MVO0uoWj3
RKAmV5URsgE2t1SDxOngZC2momeafHODWqgS70tcQOQg9Xro4f9Xikz9V4s6qsMD
pBz/Yd79RZWxevEebrYD4v5TqftpNzCW9ziFiqw7OM+0E4rSEEZ/CqHTyWFt96aZ
pjLY20kFqPerPKyyfiAdzlC3tuhaa9B8VfFrRYHqJ2u1cMh+FLNJExRl0DQLX+Tl
w96FPYg1QRj3z3dSvGeokS8TlFfkgwQGJ0pEF+xbU5slQ9Bm/OSNtHNloG/wOGAi
5iEx63lfMza696YltKV50Okc5ggxassPPhO3+Wmg0eXZ2S+wXbJZAERUELafxJ/Y
FquG6R+ArDSz12LkzGzLYwzhJfux8PYNMMY5Wt4TdCDZY+8UojKT818HA/I1N0FX
Tc97z8th0q/W7kYkLQYoTaJdurrJYehKSAfe6+eLKRcCQhgGqZCEGn3IEEm3bKuY
TtyA3YumZowsQ0dwrLK26fCeNbY2HrMbFTl1AqOkwsPBrJ+JFbS/NlOK2GyiWb5m
qg5aOvehsf+5+6wAnGFP0N1hOycIZxu5bV583ihEIzy6iUz/W09VCeQs2IS1M8it
iMO2zZ4qV7KUVsiwvbt0+hLtbw9NSAV5FQOGmf+sOUM3Cj4bYH8j6c5D3X2W4gaD
cx6ckEhwYa7GE/6knepHKO1GPE4jnyL5A5F9ZnmSea41OZ+he6sdlWpBUU+e6rMG
hlENUU8WqmWEfKilq6PU33vqweYMBEnAWn9DsOFU5gZKgrH6nb92DEK/plbnWnWs
XLPHalvARdAaU1v846wLphWOwmpZQzZe159HJ5vg/FfvYpZg5sfLswubfkL4V51X
MMvRtIhoMd7kS0x0E/DfMTT0Pat56kz/KMx4dt58gHWHy67Z83mT+3+h8U+TI9TO
ong7d/clQi7HEPAujnzW+hy5w61M864Rp9qWn06k8zgReoO3VcLhM2hY2EwUsmOR
cYYYELemi7W+xYHvk+1Yp3J7Ijupoxsd8vWCBuwlXutgoordXG8TMgg8kPwrSCCP
GFijUrsU9DzITHFajd1+Kd80yYroS8aKBKEZu47mBnWQwmw3I2KzEyRrIw36PkBs
hih7SqiG/8NSzxWWrNZYIumzRg2OTKBIteVL6nv2itukpgjTQEcel7zZUgOuAYol
WT5V1oQpDAJYryNyb5v08IJd0gKJ0Qt4OF6/F5QX3fzzuXYj6AcfnQm/IrZ+k90q
72q+opmFvSoc97a1WbqA0NAiCal3Fs1ww4GjlBKok6AqKv/cKABPWitxCkHPkvc7
33L/SeG/4wVoaX1fqrBKFI2ydXlzyCIBNMcuSyP+bdGzbS07xJUzhlqvSZZ6RXyB
Der+YOa1Ev3MOSZRaJYT3lHMrpEkJJnQ08wucd6mriVKw7MvwMKnVxlnADtXGFoe
0btRrKvoNSKfteuslgfLbc9ycrtN2zJEGeg4lxTU62HA66/hCQCyRHSin7Y4ewGP
qG1TvRQqrM8+NaKjTpzX/sIfE4Xw0H5sBcjCHbsicpNZTS6VfIbF2DZlnkWW/YFv
9rafOyyKTcCd42hxhOgOotnnNbvL6tpX55VAfkbhCHB/esyqhflyivJX5edjh7zo
X0D6N/doOPjRhkN+eIMk8/rgJw4LbU8L8ngJ0PD8a92MarzlLXs+qEoAJcn7aGVQ
0NRsAmzAMahfxWZOXPx02o8wfFPRnr7c81KvqTGXTY8gKzYE6jpNXxah6pN7YQKd
Jd8op4KxMwNnKc+p+PHzr+w8WqKhmSqnLqQeJCcxsE7GJyxzNIa6ZpdvtPw4WtWf
CvLZvexs4o4yGxoS0shP5XcPDqDtoPG5QuUU4CC8gSHR1JqehU9dmI58YhfvnXtM
5qaW3/MxhqmbrkwwezCKrPMQ+fDEpiwFqfQPFOFVGJqs512Kxo7oDBRDnPJ6z7D/
xiZ2NDf1ttkuB4m2S81idheg2ViVeCuxsWHmMbG8isqf2armr/tV5lr+rfStpWr0
pV5SnTe7ybI8n2LGX4FqOqyj8O0qtkXXQxxVESKpVOo6qDoLZOm2YKsDNsiczP3i
Tr7PeZBGgU4El7kMueiVxA76eINP8eCx1raFGGhQAYo2WP1XghkTe10MVfE4gnBN
mt4QsBDVMv1BkWfG4QBtXFO2pU8xc2fadLukv23tT3xM91PHT3G8BqoHpHOagqoJ
iQTrnEzIm8FrYlNHjISTgEwcKHcSRlmJJcMbJrO4vJQme9SZik1q7bbd+++VlLwZ
d1MCoAAQPX9bKrkPQ7PenExMcvkKv8+aRRJKbZEoEtr0UCfHRJVlwdshk37iKAty
KULe1AY+9r7rEAzyuxAbynlDx+bVa6VNYHSjDq6N8tjdEml+JktOspee+/XYs1FA
hAdfFkB5IQvzLtJVx4nYrmDpMIpMTs6dwoZ8bzK1iKMfpiTOxqgBkrkW1gOtN3WR
xf7hIcgKGyeSPOuSeqziIX9RckgVOemcvkwzVVv8Z3fM6WTlmTsLkufiXMLiF6z8
0fnWrJcqpcOrzKADmyKd59q49AQLiWctCSy1zz9VNwhTxMGnwG5PSaOpPCxfEn4D
AsC+o4F8XcdbkbfALtt1UJ5SbasPWGATC3KwPZFjJKqL/2AGX7oi1XJg0Bu9oVQ8
xoFtg69zUmHcD+Sx5UthEozwIbV/ST8d8qXT5/Az6rYUDjja1a5WCxSUKdkSmmbu
s+cUDhXy527aUsKw6Qs/RICZxHlr1+/kgj7VPXvvhSATloUXrqg7+h7nO43wFvxL
fHoKJijcFuQa5sdSM21R838lpxpgwoII0NlhkEn9WXb1PtX7rvToDj5fGG7TX9qD
nbTYiORSk4UmSMvqf+bpczlJZARsPvhA2iH9d9l6zlrTFVEudgsE+uQCksMV4tq0
FBiTyAVom07oHtsdqAnC8yT/6KPnjjBmV7jliC8vIQrhOrUjgiBoT98a2iH5zgPr
Nekqdih8kfFmk3voZBf25DmpPoH7grnqTtpnUhZr/Rurak3PkrTHreLNiwAz9o8f
vkAFJGrsoZup9SMEh+ZlvmsUBBJB7tp4Q172XXcUahwGKxhQRor8lRnzJmi3HwDW
Fiwp/rdYIEPJ+Uol8eF43H0gch5lPqOsq0ngkbedLWZ26NSMrAHTw/O2f9QDDVnd
X6cUD/rkim2WgvCRvRqkBka+WO7wx32LmwFz5BoxrNGirl2XB0WNDyh1AVwlo95t
Hqd09czUz2ZDcjHM/spddubMOo/U4IGWWKEh/RnaxZoByBsNFXWo8FwwOjylbyTS
YjZ6Pm77nzyvfQYhQxLh07zzGaIiP96OYBHsJubJVqVfClIGdw0CFYSuQEEa1NJu
ybAd79mdUiYhj0U271Y3XAcVr9/CwUdK4vrYfAgH7E3olTkAVFSfWhSSSuLrgvoZ
AqpE5weDQFRsuuwU0J1tTNuuVJriCSKTgJUCCHbLIGKGeHTE9cFaL9EALeIib6b6
9Vdb6vgcHicaoo1UJDc+hU02KIf6NHbDKmDL6RRfFVO7J2INUWxbmNurxDMuWmHb
Xe+6yNw/kqcjQYVyWM3RcRnLzBOux+82XhFOyaWE3zMsZiuKHcGO/0130BYWJZDY
LcsxG2iuGe4YdVBq37JZqMo0RtZsEx9KCSO+KwHSxRACA23unRIjbRV4g4P811JP
TA/uHq21vSgaPOw4FgslBpPOdAHrD4vdEAp/J/xB1j5a7EnRX7oUsoFCrjRjDmih
RDuBBhPgeqYJLM4I/36m8sTkmrgxncoBamMhjW/IGs/77lSPNWdmt0qHxskbGitm
fImobbgsAmKguEZFk7OXlz+bF+3U77f+aqOVfIUMO4F245+qkC4bGLtvvn92TN6M
wSxGNkxtLqc9/PLtxKXHQbk5xCcZass+kdQ+wL/0IT2GSzzby4Ny7nFSPn8PBcd1
SDr7m83i6oYfBCJuxhC2DtM4xbvY1hO/kcKrrsQgnV5FwKVg3qsVnY1UZgNqVb8E
6atqTM+ZpJgGnRj+rWarb90Qk6bOaKKT+9yP082p0g3ejDFNqGTGsmJGA7ejoYVm
t0+JcxHm9iJVhvWB3GLXzUyHJRRllLvxLIXcyRD6m0t6dYFYcZbH2GsOQtvXcjGj
T+33fDAVMFQ/ZuzqKzSnihZLbRHu+oSCWhgyQL64kIfIPj+HVH9Fxm2ExE0Z9fvd
oROqh2xDp0DK+IDy6JC7mVDFOPgO6/2RU6ss9V7TdSAEaZejmqklR8zMiV8UtleW
MvXY7+KJYpMXGiJCwpCAIIjHofxWBsiOsiE8lzYVy5FgAi6BVAIm38gJ2mzc8c0h
SGRcgMX1BWU6LxbIb3Rryud8ElrJnHh2O2sXEsxWsEXtfIr+hedaWo7xTSbbRY3z
Xq8j4O4rp0h+K6kyq63RNj1N67zsUnhQ62k4g81wFGOzXkEonszqpPwtyc1daXJa
kmfK0GtQsQkVezdWkguRUdxRnisMplLd9lRqVwZTOMLv8VDtmbPB0NJSoTmAd4NC
7rFyM6H1pwRIkZr7J3pNpLgiAYsFnR6yLQb1ELqo2yZevbr+r9mn3rxf7INEwAn/
coDYtESMab8bpMZ2p8uGHLNANbl7DHD2OIkRY7z1Z6+F1CGhpH2ZvyckO90nU1Ce
Q5wk5YNgNUUdnIAl4y3TFDnmzTefj6ARGycWQW+5XRuWssAQgKs8kTCroqSkNfmT
9FDiq9/X6003blwjrW521sr5aOvS83MGd5Wr0QzmCsXo8E/2XAmepPC5JuC4X2C6
rl7lOff5DPGfJhz2X035wZKyZt/s0VfELDLkCAfidJ3EMNnnJuS+SQYXqgbKg1Ot
qRTW6a8sb5U/OkbbauluoIVH9xHfC1W45wSPPId7L1602552I9XEacXIgAznfjly
nvWZtRMpLsvgFK1QH3y6y+g1WmmMBEHAbWTuIiDa/ioKwfuULmcAeIyctRHeAY59
LlvZtWF69kx9SAVi2yu+DIq4UQd+Np5RKsUZSGLrYViTGmesNi9CMRe1tEBdWGeb
QnlFY3ppHSAf7A8XbHQTsMDJi45r43+iH7NCub54zC+dsEIqDJvAi2mWVsTpq2Lm
kOZVvJIe4hcJ7iAtnC5y2PPILbkh6D8rA7eYRruLg8O3oAb5hpG+UKKeMJTO/5Bv
1gwR3QMtran6KCImtfhxZOBdKUfjDIFqsfXIoS8eqoFouiznbBWruVnwXkDIZ8T9
/VTHNcglulfgdd+kNP3mARLzi9Yd1PKZq6+DCLBmYVcS1gdrOMEIWMgF0jZPbak+
hNGWZXJqB9WpuSqvTTQeRY1XOu8XieTbw6yRZIJKaJ2z6OkTG7nYoCLKDtQ/Dd7n
Ab7eZS2771IzhLsxg5Wnle8KVYdsyUIIHTR7+w1fh6Pyb91UoC9Fh2nh5WsKr/OK
ktxQsbopsiDuVdq4hKbBL+CAb0qNnkbmfk1pJrMAP5Ba2YeS+/IHN0FgndN9tdag
jK0YKgp004bElVyr0aSI7Vme2r7lmNKpkdGpGNHJyDdMswLTPseSGsekKaGBTewI
HLwTBX9zkuRRRiJAsS5FJN9lzCmpH5YJOgkpMZdqIJxEO3TQu2vSh2pwVjch+7t2
InYbl2jwvz3mfeCNW5xUsDW06XQuaDm4Zfz9R5fG23JoAbI33K6BJL1O55EZW4Rr
yBNhPFmVLyWpXOUPCeIwV0YAzQMYAnc3Fi6KfBLm0LyWYRVxCKaByNcDJ7eyQriw
TqlqgIGVts+2EAEbdkd2F/xTdncZd16/5L/dGSQHnk7lRYywOCpXi7C73xjsaqv2
m4ZZfnKHIPLJOH6lq3jST56Z9WgxozT4l1qxnuifNqJqWR7jzrWSGjywd8XAdW1C
VuHoM+77o9pTBBSnU3ZTsChG6tB6WWd344sCvKJ0il63WCCLHc3htjknuOfK24ox
XheoJfrdIpJlQiIPr/CjJD86BOnNDH+NGzoVH30X9YScaL0D5UOm2L7TIB98XduB
ImJ7dvPPjS+V51FWPcytBPT5IGGLrs3atibGdh+Z0USXuvSuol1YXIesLA00FjI4
9/uM3iiBogV9Acd//gG/mNHM7Xo6n8cOL9jURT8Vsh7vs6T2vCTkrZBLA27zB1EH
OjKQDOAG+GhzFkcE8Pgws14FUak4HRKfE2tvP3e/V0hDpu/MR3JTxJVdq783XbrZ
fos37BQpgVnjoZKkMwU7ERQSEsC6mOFz9ZX8vcfh/r9tJv8zAom90hAStpA9d6Yv
xbjQAzIH+nmW3H9A49ge22sTDOrgXkXFJp7baTJkTF62b7jtO600S6//6i0ztiA/
4VSEfZywJJ1QSmYoLDzPlZb1isVZOgMQmAQPlEwjNv7dggF+cCK5i1lx0XY3ev8y
B1GDpeMhobRs6ZK0nF9oXmRj6UAzXwh0eaiXppTn6B1L4xCp2Z69C89yBX9V4+5L
j/8kkNMIoFE2rylNrK845fLMzLWRaIQ3829LwRNSlf09F/ddZCPaWJsRw7b1ePQQ
KhZAUd366uvSQCr3yS9RmgD13l0dyXmlQRbvPKR03AyOa02ljlqUJrtWoweiz71t
4HHCxsBzKGwnDQgng0mwm8P2PQ+CpR1XcPz8FTRAU/jPp3+utPJoqgZuz2UJ9FrD
mJLOQrjFcnlQR8GjAx849hiqycnERF70ETHFwGzaQxwo6+6aM7+Fcj1sLVE6OAA9
AszQ7aTOuDxZfgEQrAZhrzu4BwULapxt4nt4cbY1lHgatmdT8xvoPLplHKOLj9PX
rBgdrrRBTNleNG9RqsGLQOp6Lr3G6NSLZH+sGS4ncT4PUnuSVN5bAVhiM4PTfesd
oO58WApW3G1i721unkxtCOXJVXcXkOqy5Uy9lOQ7W+1kdCaJH5kpnwP4GpNVkIQq
He7drgDvrhC8X9ut916DqjFoUo570gyDTfGwN+vtRqDGBuTGaGSZkX7f3+Q1nFQ2
Cx4JsDZamCkgtO/82u0ED8pebmpn3fz8aqDEI6wlHRU3G/fc+B7hzM13l8/qez2r
QoFO6i/ntiotLvjiYqey6la3f3ncEC3M4YVYC/4+hB2jYSpZXVIhyNMRxzMQcYKN
jCBd97GuhaGIg0RK8dS9zAtPGEjobgrC57+kOt0xQoHUl96F6dlz9QWVWRGxAVOZ
DRW/1AQob/w0BhT/jgXAuHLWdKvkeaRCedCEESRBNa88I6ggjfGXvZeE5E1fA+sT
6e43wXc9LA490i76E/SAAr0vqTpO9n7SCFsmgNnwcOH3UmKKHXXmyoz8j+/e1PG/
69bfPkH5gV3VFVoWv3M0DvjgjR25diVpz6McVHOvb7NJ0MmFG8FIcGNIu19K1iZd
7AedyCBmPbQ3xY8le2k6nqjzHIjc7CpB4MD8qSsyEXJAJRXVrtzxBuSJdQrM5PXm
AMFPoEzwdpVJ9NQYGS4iuFOu6QlYamzI6E+sC7+/qY7mIQbWc8OeBtMpe3o3dEV0
iVVa0iWasqwlk/ALzWfyIJ/0R+GShelBDNPLm51FZ7o+6bFZLXl/GjgKIc6Y78Nf
I7xv4/U7zNUv/Szbeff7aPu2+C3+OhnrZy9T3Nd1YVcLEvhsbYGKf9UmhGrs/aUR
5ewBsFmsHSF5spJEz/IMkUwp7+3NR8WXIB2hyawT2jS3EOTxnBIHK9oEZtnsxkVj
KrhTb+DhZJPoVhU3G86vAEm6jyylkZz4Jb3YXpvCOC08J2Cw0D4TpZvYKh/TWOEm
Ys8gaQyZwNTxwnX1+C/tXYCETMvPeDkeZOL9R/uEmQqUa6/1xzLpRTaF5xh2psqg
uDfFv09X4eOc1ZICP7hYVQQRR7XmcKbUaS70b9FcrWvff7OmAr3vlDDAKm2jW4Iw
OcTBcvt96sneD7YkdkBTKlXvPmIym8kA/U00OKdo7kuCbOXzB+1Ne7WhSgdmMmIF
uQrwovJtp6FpaDbsOy39qK5NJTCrHhorduE+ygbl+Dlx8m6+tFkKVFY7IzKTzQzj
o1kjuLnVyGf2OdD+AaAA8KE37KCt/yEw9ybYmn1/n/l+R2QczDRz5cA/I0JxyYK5
eS90/oOB8RorAxa50wuVf0Socsxn2hrXxQdMUysFUs7DUs/cYgp2hbkyC5vVI8Za
ygURbELFFyEq5+wkti1CodDUfVnFxb/ABLqZlR4kgstnEZYHrxREggxKCHdK2eIS
j4fxdrtN11Y0NBcr+lCD21SRlJrjOriVP9ptJlJdhGgVuotKuzphJgvYqidb8i1a
gQa9cq+1HC5Y8MaOnpwe1UID1cToOo5k62oM9RUUyYMeQvgTSAeCoj+Jxvz3mmqh
a1w0Ohw3B7snftFrNkZEgRCRaLMPLCr8lerj+4t0tMWpii+qYD3/Batta9ZDIsOl
s9iEyekZZ7wXsd3jrgN0BFcheMJc/42wE97jymV4dKIjmzDknUJg2ORk/HfU7QRs
jlQRa6cANNtWDs26PmupADXNBb8odGe9kYbjr4csVIkmLiA+/4jtqQdE8jSK6TeI
J/MWxcSNwkYJRv5pEHVk5aVSw53gdMHTUr1f5hnkldPd1/gzXUaWLNe+QeK0C7rj
/dJw5uZntOL9t8NCdfYe+WPZXuVPAset0dAxDzOnKfC5uS0KM6oX9+K9zAsemfOX
kH5fSZesuX28ZlIcfkIR5m9hOvRNEoDQx28UZMA8ZLg32c1bqAMozvdXtBOv/YcX
qWascS2D2NH0yMLmXY0tzsOfkv9rwHkNEeGCnW6tELjuv1VPpPL4iNT+gS5U9m0x
H3u9HxqdzU7P/pr+NhUZcB4iRhPEOaG8KUYgm2xNMg2Orz1B+MaMPebbjCoo0djs
OFYnLMULsxq2wRfQGNYceNKGIri7nTKGY7eimKY/9P4enpAr+DUcAWchpdUX58YJ
zApISrqyVWbrxbD9u6V5kStQP8TePFVfeDljeJriMfzBzGpa7yB1oOCc+/2L4n+z
Q/MnqTNM3IK6RP5KZMViHwBIlYK1sq2nyP6vFbnVmV6cI0t1QFc97nEIcT/zhKnu
TpYiBOWwJczxJqtzT/cK3UAXNwZ+5jD4lfVN7ei1Qcl279tezr8XVnlQjLhpxXth
xvvubwQI7EHxQReIdUtYd8j2LJG+tnUA6U4USITxe5ZdwEXuhL7IjYb3+LSYRtaI
y3xoR1DYzMH36YD/CtYG3cAOpTcsrHMr24bN7OHbiMP4b2QsI29gMHJOBVpqbOP2
1cKd+d09anhrQzE2VOK9abK/hUl+z86gunKo5P+fizyBYdWsui76gNVGEr1xUFxO
sMAj73TIQmGbpdMmRW1aIXzy3rhXwhHm7d0tHhbNLV/a4CgqgRpThvhRYgvpbLEv
n5Uk2CcuIGdVKWdeWFy0KRMO8ttD4Sgz3a/IcjP/zhZiaNWzRf5BGxnOQ+ZhNndt
6aPsl/p5Uz6+yS47cqGccdapvBEL6jl/kEQQydphgZoF01wq6gUaJeGw9IyYLqfn
H+oqr6cIyiMSbAtKk9CD4+JrappBUGNFrZW2PKacPvIxlqaXerp/0NbE8zmla/Fo
ATibPzijRqClniwLNbmUyklaKsPMPEYQEjq3n9I6513hK3ySSKkm88Zvj/OAfCLH
pqNnAs0V19ctyald3TghYO1dyjACKaEl3weAApCj3nqviXL2ycaMmoVIhZW1Sj45
E5stv8kGq0V8/FUnVTKaiWxLWbI/kuQCo/DxeBWvmslDvAj0G1qlm0DywJDj4bWF
BvfMZtNs2cFfD87bhmkDXSLkZOyBYYp5yvbkpCm41xdXHT8Ccq4HtydeJLAfnJLg
f3wVmnSH82cMgizyb3qelqcZLDB6uR8jIohLCtIyq2c8tynE5ecrOG/j78SjCtlm
AD9UJOB4lem4Na9HjSHGfa0tvpJESGlhd6qIzFXcWVJ7C5K4f+bYzJxIsRrYJTnC
fxUfbY1RtAvNXsETGui7p62ePXf4yRxOv2HMnE5/MI+C7RJC0q+6zAInemebASmb
LAlYPlw/0yQdaZdjC3muA35cS1mDktOMMKnmvvYMM2zJf6Osd0JpMHIz6WGLAmbw
R9NvCif5bUkBWcbRF9ei+5/qfNeL8JMBswkFYfV3QGjbMUheq1sE2xVoIKDyIgk9
W1VSI2R86FJuPZIB7TgPljbQapzkllclpbPliDx/Rh41iUfCm5V/+6EAnsbm+YDn
SxnzhJS0qVJnXho7DPeh2a78vy+XX8cjzktrXNE7dkUJ7jXSgZX0QfGnXWQKb5jX
8vT59BYcd+kPockRYPuiXphrNGhBxeFKvOjvDQWI916Tb014qZ0UskAdTWFaNahR
G0r6DK+kZBbpwtwh72N0MJP/RZana95UZg9smqWsUH1G3ilbAFCzdZClbohpHxfP
7h+Bv8tpHqPsAv0lu5kHBNm0GMRUit2yHm2tsFMYwsZtRX4zZ5kMe9eqyQNIgdC4
/KY/vA8Y6NRpnT5nEbF89c4NZrVEMEHUrTxOBnn4ejdR5qiF2Ldr2xz64u05Dtus
EyeyZizz2XheMzRDKa0C+dXAddTIf1gbrxbEOGFs/j3Up+bjJDESARdDf74hM7qM
yzBgVorrdx94oqhUPb4DegQzxIMoA9J5W+6CNKr2xQCPEH4en0UX1TB4YOVezI7y
pYTCcxCofSH2rVLECaI5O7RamL1QOYgi2zCy4kWP5lk2GkzyK1jA0jjHZ0PihAmD
jbighI9iuYFVTnNDvH1Ep2xxlzaxGWxiTBxKdd+du4UWf/ZGUoerDDYhRq2zhhWX
+Jzkjbw88fBpU9gkubWEowlp24dx7TBjv5TVT8zUwu/6BdAP4p1RqrkWCjMJzFPI
nwm98cz03De5H2rTHN3G/8FuqVBCTQhg4Y6GJ2R5BT3vrrI4QQ0oudUp7lgHbK20
LlumsNap++MO61khuh7VUQoTolLQYdVAJemK0eBWOlLfMMvBi+p+/W1aUpS87oAE
QDm/LqkwkbLNscRHk9ad6TZs8G8Wenk7ZsGt2I50D5hkDclWQrLFXpJ341Kr8X9z
XGv6Sx6wVihlKANcbYbtZL1XlWOgEbwQvn4p8WHgJ+dMd51VSrLjwV9J1nHY7rbw
OfPJEFSqdeFO+Eq3hc9PDQ3wGJ0zQ81jxNQeS9ETEPu6PPjLH5GQtkfEV+BZ2mt6
33yVyvV2fz1iJx5f34e+upLtbHnFgZEzrg72JmN3hRo5NPQCmgE5tXv4VHC/SWZw
9BIPRDPiFeds2GM3F2IeAKvWkgnDTNTrMegizEotKs+6XxT9NesTkteJBcaCjb27
UH8NCG9c9AH5vM6716oIaXdYQlk9xZSgrTrLSWbCQTbw0dbN5Y1BH6kXJvz7fS3b
wQx657VcDsye0szSwdHq78kG/pGt2U0o/BoLjPcQeMtPjbu9P+s+XXUyLQ0W/jzV
7N32Qa0zu2U53tSfF5cn2LoUgrsaYi0xDdTK3uZHUFuEBliFGY0LoihoZ37EDS1M
CVMvOUDJ91WZN83EuZGnA4Mf3UuiZAvzusmhP+KGinK5laQ+3qRm5ckvjluTHmUj
2IBPVA0kpWAop52GitPCYNnMcHe7gU4zMhShyHvV31QpZPEbKigy1IVy9DdQ5P9L
cOzFmj4Y9EpBNn1kkiLR0SPY1weX5bakKY0AWGtN+q1TkHpdDy51bZFGKCeZ1f16
dqJmFwKqOoUr52GdXpmUkj6lnFwHBUc5ekTFufLm0Hsfld2rgbvoCZ+1kU7tBJ9c
IOcT4342dGwBh7iM0Nf2qs1CqvCXJj3os1laq341BEv2JXHCXX0SPUsuste63/IA
w2k3Lcthu3jgVOwhQO+eQRydB0CVRodcyD3dIbD3SrP4nqCTzP6z9yLyrvQMfy2H
0avE30zl8/jl/paSbzLs73rnDdOWmriVJEeM0F95OlQQxeoM0/Mx7zCm4Wb0vf1g
C+XbxHUAEfzINQtuWO+sdMoYWKMSNtwJwukjP/suVOVn63XaAGVUMihEuQINbo0u
3nUg8NkR2V8M0yuXI82uEHfSxZyBWHbxtROT7D5bVgTTck61zY0sjY8zTlT4XS8b
2mZddC0vEK8J6STeRc1z29SdB3J9bamgbwL0r8+dNSbNgkj7dneX2blEbLIKF/A9
WaaTgpsHodA6VWTy+HXdtT19deya5bUaqvhUii1lGnWXYW8wLzHD3XgWrs1nDFVd
FOvt7L8GLLLp7GKTXUeBHHlwK/63ErSFpbF+NF8Wpb/tAagvQJCRxQ+MPPJgiFjZ
k/Hi+FOg9+kXS00fJPpt2dOVtAO0/9xIFoPR5WdTZR/rfxEBCaxSfdLRVWEQTX7D
N6SKWPdkp5z6P+V3j3tpv+qGo7sHiWH2fdhwAuWBqVyul0py7VvQQheU9zMXdTb4
8ksBGZ9mR+yJrD7ECOYzhxpktZK/MdeO/SLsHpR44viv2zHwL2WZegJUMAA3h1PU
JM00XqnqXltVrK/GY5ExrqmjQD+ALcwwM5vfk4wIz7dia57VvHTCrZoOd/kXpt3y
CISoJdTXNmpsQ0Dcz0iiHpaXcFeFKu3H8InHSXn+fSPMd6lr9B9mfRS9XH/M672x
imbAeiD+lALvxiyPLNmlocnzylcEKiMJ9UVyrdLKOU7eqtIdSMdwQFpM3KAa0LtP
uEgqVq+fixxVZj3zxrXY5wHZoSTDxrXubj87o13OY1R7gTCsCpc7pTQDCtDECSNP
ZZoiuZ8SLPhZhOt23imwujJxcp7YXc3d+++o5n6g07Le9jbjJ5X39jQVAiDJjzsj
TrZg3M4EP4alai1Qh3i80f+xR3JtU5Cnbi46dlNvjJkcRLoEkOYD5NckrMhO1HF2
CcSZsf7yW1nxAVqt9HUej9yOq1PganESjXr5+rv2SfFe4HGmc3uFmhf9Ho9MS5pU
ZtHzqr1Fg7o2UAms/mCi1A/JPAwZGOGboN1+p6M1Nb5fpxIrefFEZKrVwe/SwuIc
b2SCnLxYPCd6ARbgEyO6qTQhX0gmZZPahkBHULHQuiWcn270cJ00U/eS4onjCIEs
ULQLIZprpOpemo071ueXDsRsXZ26Jx7jepiFl58vm4+2neWbFTzuPfrj1j9Qwz+1
n/Es10lnK/FEobiqPJEGWYJwDAPycO5EHK5p/tyMbXJXOnxtvfy/N0cIfVSGF4YI
v/jkppzq3iNs61IfKicsxoFiX6UehDD97XBUHzazAB6tFbKOzNctoXBnFUKxED9u
LBbIwy93vxZUeSnYAxuX8w6Dm9SMXGBpfYdjr/Fv9g+5RSdVefR18lcG1ilvczuk
yjU2EMKX+ZsUPgAhgr8jgSivnkbTCh467N4PwpsfGzP2FqAGLW7GIStAIqep/G7N
etJWNZlK9ICKMk0quE0OMOy4eukSbVunhNZsE9IGmYrie4LoUiXbpy7Wo2EME6qS
OdIDPi5gCuatCc8+dutGYtoX4SqadeCmztCm1MQbwKyWYfbUS+glye0x737+8Y3p
uAoUsFjn0nkIMnfSq5UjtD3BaebaQpKcv1nMbPSc7THw2IXXU1wP+Ol0QfEpHG6z
Q1a+/EdD6H598hF3L5Y/4agg/wbkmU/oS6Hw9453X3e6GrqYxqmeVbxoAD73SWvq
pu/Db7Yh3TkETc9Zwt4JJnf+sWG1H/ctfAn8OkILHKKWGefE6YsfGr8tRCmU5V5u
+thJRlWMMf7xml9653q7Uw5vVDMJOsVsn0P3TDeP3240UhULPjiKi6Ll4g87XIsr
8K2ROPuSHdgGyGVQusl+8rusAGMJtPydPQpIAIi994BYdO8VlCtbqgm3/BdJAMW9
HxtiqVfZCJl8rbH48kCzRz4RQZKY8RLaFyMkQr3MGDDuv20HAhFjuVvK1cFcu6bL
nY8ufFFCIYk56WS604Gg9cucLcwOuHDdXL9l8gqkk4GDouGf4EBTWbJBtOYIf3or
o3iH5yAByKqJYJ0xiO+GEkdfL1mCRz9vmXEz+r6TcmxZ8rou+vCLhUWzmWp7pEvQ
fthzMMzx/dydStvNZwyJDfka62AYwRoloKDCziOACiLplxflHpJya+RnC5AXpxvd
8iNS8vaoTZcfAQhWVlRVyZKicKGZiC62jsP1hV0rWlFX852ZouPiPmeynqrXPmvI
Tlj2k1tP1tUf9AE5JvFuM7Zo+v6+dzibxsc3TLsccoaaXEYxnRatsS78SsVh/UNd
2t6VEnpvgXOmxWec/N/dwdPlbQZfry17odFckHGqIQcaZmP6a11sCvzn8PeltKu9
VHOtJ2vtetem2PiLqU2wua8nz9UZRaiNMilZZTGqDhuL+ev08GbNv989KVO/ayVT
5qcHdSMVx7xVBaVMkvvMvfEzL5gcmbWHfVlDdlnSnPpfijtjfICkzX+IfiWcn+0q
8zmcs3racDQfmmfFs0RKcJql2sw3HcWH4XdlQ9aegMvxPFgBzi9OWVdL69THEI3l
+4Uvh9cm5IgvGTXETMgcgz0VIfdZzcp9smTASg4i1wONx3uGwt2xDoj2qfE3iSop
6s1jKfComzX9sUPYoeFSSytKYRHov5oG1nB1ptVwmTuf3BJtFv3sxGiw4OHSsBtO
e8EY9Byr6+fT5KMWrGtYGhrEzN9PMy8gR/jZm1+Rtd9dNKiakdFSvRUXrpPQh/Iz
O8DiCkrl3vvoGDYgWalXBKTnGFWEgfwK2SPVUabmflqCnXmleFVVoRPuUjBwSSlw
8ABTPZnZgTn3w9xKwxaSa/PnLLpqyDE/oz0KOPRciLPHy1s/2tL6a0GF59uAPgHQ
LIfSXqwWspFVrVqeMwrXhiXvRwgYWGe4kjWkEffgC6w7N8v+7cC1OoHvKPD+UK0f
tkUfGt+JmnxtiTK0P7m7ddUQCoMuoignphJ/kAZDFBdTFPDEuu0TEDK0OS1pUZDh
BLHDIVtIiOT0g4AA0MowOI9LSY9J5zGgxclpg0O+qHM3cSk4tkV+YXDkf3F7JsHF
EUcrYYmKzieyCfXl7WUihyuOw/ewJ1SsDL0gXmc0m+GZRvsNvDdFAUtEIvMDvKWR
7y7477g/HiG7IWW/NC8qeuFZ892siWdlzMRm17514rP2kTmRjBt8phsWxZmD+lZP
8WSFmaRi3TVASXwwH01UZCvBSD4vWrQ57ACk3xsKGRhhZn6Gi9kGiB39Ed4pmSsV
itCwHiRgCPhHMEzp+ivt5FYkLShE9mplZIhYCRFnQgv91ojOOiBn7pJKXKA2Iz1Q
rXFLMhaRLWGzvoe26DQQ9OP/7TBdz+QafABlqBDHdX4befLjwrOLPbRgRieeWLd8
zH+TVexl3qOICiphDFqYNWsjjBkR9tpspgI+E4TXCXwj4R5S6na8ObTmqKNjntjW
tN8/DKEeY1OThK1L4aGzm9l63gjkJGGcbr/eU76SBwWRI5nz+TrNc/Cgta++orEk
bg9RcEMpHeH7A0sYhRwqUdgkmvUYAk20AidBKRGa16KgArsQScbVAw/iDfw9XYMR
TFMk60Z4vui/PdYTpzVc0Cd0FPVF3KMpj5AJxVo5ydPTOCYaDARpHAuoINwa7I48
wWjFzbRJfe85cDWupwMZ1ZTbByRmaBfu1/F9nNcWtEJjgmrvJbIQ2zfco1lSitP2
y6D1XEqVD98OMCxLvo2LLrlj9C9v+VLMrt53sy5hFAgsbmqy6l9B5uSJc7p7qBOr
WXZI0jHko4Ng3Z5EPKbyqM9jMEWQ37oEwY5rW2Q0OG9jBlzAicsyPJkaJ72x5NfW
4uSx6xvxPdhJGt97Q5Y9Lv2Ok6tQTzQaf7pp9/l/CeIXJey/wZHO97ubv3KGep1w
aHFCPVk1rrev6fzfHV4yomsQKESx87U0m8Z+fUotr7LgmXr19zSPGrILh/cOGqXr
dR+BMsGaYr0lLckJdluM7Vlpw3H+mHidBQW7Y43j4ZOzjBFuYCIDSPUzY2vaUsYU
x24bYvxcQLce5t7cqSdalzXHlDJtF6xRbgAUMmBpHcLSe/2AV/VoRTRWcbLxSXIT
eld2nUrl1e0hxMbRLxNeIp7GNVz7bmlouhwTSMyXjUIvLgl9beqvBCbsgEMiDx8x
oi1R/GGhuxuQSeipRvIr+NyglqOi1ClWsYeSRIuUCyU9CrtHT3VoIKZjPsh5ELN+
A5Ug85ZMZq5h0SmP3QRtsLae99yXqWRoeQtw60wAobyg5Vi6pZqD6LRLc9IiLUuA
LmTcJpg7ersYrj7dIE2Q2ZIfsakpssJdcZzp8KcVPoe0NTVB8L28lddiDqadkqpA
yY6pGzVlxRBiYkVoL3p4HshEFR+Sil6ivqvtsCYikNt0Gj09wtWRhEfD1jkIPxoq
5Eygr8vTk5FnccWnocZE7rZZ26AqsfFdhpbNN3RKE6zFeJKP5RyKQhg7FB74xmfr
7rWpecmIkkUZGLulalbXhTVzdfZBRAC8m67vEnX0klJKfUCRG4X7aGMd5xJ80vXs
1Y8PQl6uEtjb9uQt1QpmEXuYxR1Q08emH4OZZ3+2E5wh1M39czBC6xhjZhdqgGVN
pc6lhh1iRwEA76syyIRI4p34v5KWcVM/SDAn5wZF26kSFiRRc9uDYCjo8OBuXmru
nmglKMDyiMi96fyU+v16TMUxAJowrThDXQFuBy/Vf7wQmxNKrUQOHegDFtJCXVEc
2xcvr7cAdKoobi8GAhGyxT2Ap/ezhocieuHs85x2336HE2Oz2Z+I2n9auiR97uG1
aSTKAf3AR1kYZ0uSsY+OrrRax9/UvpFGUl0WbaNjc8XgPxRnj7bdtZUW5ef+pgXJ
R3t5Ngrmg/F40xDVCxwCtdN06sLC9i4iPCuF2QQS9LTaWBNzGicLkpmQX+N77stL
STv7WtFz6uJ3SyDCaXr39r7F0H1xk4dINTdt6rkWG+4Ov6nlzOA2CZLsPP+5E4iO
9D/jswbmAkcqRTzHR6RokZ3rmnksF7MG3NEkX0CHmFZeUIKgsmk8nqRrmRUXfKyj
SG72NKp3Iuj15CxB0ke4LDsv2L0ZnMlktrv9NbHvzfc6YuLUIOT/pdKp5NpBTGMx
L5V4u0E7eKXNjQ5ivTjo+p09Ycc8Swzk8+x7VNFYnBFf8cSJptAxUw/5b5EQOJj6
adZidQ2JhYwPEOUfBM20gjRYqfDaO/rFxp8jYkmjXt+ZpFMNgt6u4N5AnQm4NXQs
0sBcRKpLsh+1Ijf+v3gVo8HzJ+7vZpuDgtshRKOZDUG4fwRcqt/FIXotYL2lGZSD
S4rQgAQT0UyGCBg1pjGMjS4O29P6M5gjARi05c4VZBy7MdfPiWFaPDuzF8CIR9nz
gcprqc+jw2508bHrg8YY79DOBeJ97kmLZ5RVOM66eVsxwLdUtbl0ZACiBIW6ASPo
iHwXYvGbmHTZgfEbOOsGgHabPhQCfmkGagf9NRfvE4iZkzNbyY8oT0XJGRoAJo3l
+OEDeT17L6gxykE2aX5ubfMqBSymx0lLoG787T2ei1FRGfJFFWY6VOT2JL0A/F70
FGbnFsaCKjUoF+ohQvJxSnrAR6p2RsaHjVAu3R6ecxWcTtojUgx0cw5IR74tDNPd
2M1t2bgjHkuJWukujKPk4jHz07tnyZyTv49of/F+/tFHzv4cPmVq8XVE8jrhznsx
es6jwAhn1h5uK3Wys3s32VgAVFgUAwOT0FkDm9WvtgqpZEKR+iLXonRZq/UU5Wzq
S4J3EK1NNb/7JNpf/+5zgUsTv/VbbFDp/zdv/OYS5qY+5fPNch1wdSrrFPEUX1bx
XdvJxNSnOF8KKyJiiIWkae8KCxzpOh3XRLurlL/783sSgJN02YJ8v8wZWB23q8/R
kAWpXe7zdTWtwikIxL5FL5MnYYdpUcTQZ+cVdD44JJvVtyPoYX+TY/nfytfWY449
48fmILWttM7AB4/z+bTshO0dGRj0BOmoojNX1SxFB7iN+S7p3hNpIIYBRxVY3orL
d7xjWCZ7HJFG5yEGd/rj+BAH8/eOAFmXA2yhXQbqETsGYMB73LPhya8/vXuWjnLb
kysfsx8vjabUD3xq5Rep5lrCLpczp+a1bOYE/SgG7xmMRO38nNpVo7vCkIwFmFdR
vJNYZdxfPlkwzuAW6WpItosE1JSs/FEm/1S7MmbRoLsmgWGzWDVk00/qwp7lV66M
YEv5d0aTK53qv0uBbKjXlg2Z9nBYE5eS5OBZknO0Z7lO7R57TXv4dGr2wo16q+QX
rsydDkqAe6SsZ9rLSH7R+2laEvoBnrI0xIB5POWgGM9qqPoD2TRg+QS3LQM9M9cM
Rxoy7mz5Tjhb7NW/X8nli/xocJStEkSzuOlKb9ipsXEhYXGkKYDAqRDn4JNcrqi9
igU1mMmZDbRWPrNEwdPl1A4XF+pmCHdu5Jaf1lgfM1F6JAfmL4QLaNjukLLRU4AF
LldcVVpbPn9N2adOoOgC7lbTCUcDXVL9dHVewsx2MCqwUbzFAPqd1Mi+QS1yMaN3
reMeDJSZc7PZb/YijkKfhtuPS6qneCY/aEBj+djenszHNBJj/l5O+yYVWw36Yiao
mhzXpEJDzKoMndyXKV7jA/oEVsPUFhIC11mhh5ggsmqgqtlmzrdRn4pJ9WAu3NjF
ra0+moNaJ9HEjYrRS3Hh9mi9b+VilOv3YNZE479JHkyBWhnOisL7mttKtGd25JE4
A9YNsgqHbuDGxxxeTKNA2dgfW1BL9/he0v/iP9qAIiMlriaxPffIlz6lYfRtv2Aq
n40odbmBj7kZOScBhUobtXFDI/+dSHfDCZ3DJ2Jew2GNcgzCFmZQQMaVJUDZ0863
YobJi3hOm97+szYDg9aGyN0i6Ao7cMFfOplgWTpS9P/wE/QYLC6Xu5toMV2K2/uj
z9maGYExGfroIinbPqRpyVl7v0cNq5GqAltRDJf2TbxMmPiWVfyJIfQnM3CLiJjZ
ZSSjK16SCG460RV61e0GhRLanwFYCTRvVDEl5cjdncbr36gy/uMyHV/S3wEfuFiz
gNHwjhD5NvjFEPk0e1dF6Eo9NnIo/P45FvQ/sSKPfOWCwVhF9kiSWP13kh8d7Zcl
MesWdDdoc2vBiR9aBu1+P//OPvMNOqHe0VfQB53cBjOzBx51C9U9nZHM20enfCZ2
GL4xgEqF1PJdneQzG2abEL83FmfPTCnfovD6uW51P+RLo34rqEXyEPLJqGCyhRUb
sSeT/2jGwvN4GJ5jFDeP5iW8JYap0T6Im883RdLugGA2Lkjuh8tVMgfPuxxNjjXq
CU7v3CLb88TzYIGfhSL1HhPoBfedHNRkLCVEW9BOtRQXm0hXfqpSg2qCLyWFjsIK
sh1ZtkT0GTQUK4wcLU9LfvF0DCK5WDeV39jIJlu41Wa3Xg8fXp7Xl7vWk8zmH254
x3oc69NElbiEBhgm/59FNZFssMdrBKgCKAjBZ/I2B9Pb3FJ+TwTceqWfUfIl16Pr
wAe9lIWSYeiw6RnK9TDgfmVCyyIvRSh+opvFOtHokeZo1Y2/EPYZlyvkW9OHIhvC
5eMessaW3njA6or8MyaOLuUxOLOIxOjItbtM9azyDQNh6WPoHerKGWs7PwNoJLgu
1oxXT8KyitoOnIuGZ3GE1X0Goe2Wr5fC28VD5MQ2NrfGbDSF9zdIzGGUZvpIGQaZ
LXvInDV15ao+d7ayHLF63I+gTmncZJQQR99IsMxlIDg0ysIMVD3sYsATZ5jTnQar
YyctA+gvU0p6oHh9btIUkpK3vb7w28uVxWPXMZFFkAMnwj6PzwHJj9sr1N0vN2a4
AgxreV12MQE/Uu331rwd2/sOU11wAFGjWLfZG+R02LQqvEXEMCANN3UOrQgS6xn6
GHVX+sdUVFRtnwXfxIKZvrz85akqg5y3yPBgnT2jKULM3bnkuoZ/x/rEVOw2NFIg
U9dQxEGpat43yPBfOSzPB/3n0HRWw1sGF8ZQiVT9OIPRm9E9Gr/xxafsjpvyWJ8U
b9wbnLcmOrvCLI8UBO2/RGEYqB4iOt1L3M8/OMOTDKrjSocj7WZgzrzPG7XUP0dN
0JqTONzEEUS4CJ3JA9Aiq7TsypSixCOOhx1NKjzGLfozVQ0tPQYDxUB8el8MH8dN
kcBE/P6lm2bwlS6drS3QPpXgf23fJsZjoLC+4j/tndqStV38zDTFKyq7iD61a5l/
p0kA/tGmWKM6cX8ad6aBlLBGl5rp8pvOrSJTmP4J+vnscE4KaHw0GHea0LA06yQE
ZPRsBVhg6Qe3f0id8By0vGQ6jV7c/YhTUeRRqxh2SDwVCaeY/SU4pp9y4uCrLdG+
3XEeNs/SPHreH5WM5gwgGRuCZukKQcOzuLNJGAX+fxsgPwPUdqYvXXCTvVqmQ/we
JIiKtWgVFzb2EPYOG00Udm2lcp40TuevCWL+4JYetrqgy1VrnA6cxmK1nH8qAxZH
r1VabnFj2I7SrpRTdSsjLmmWrt5TMB4ZEjKSHASNANwxIVD28mkcOEt1NOjFVQId
EaMw2dd62rsy1z3B0LCEdlrc9/PTErB/P2jmEHdhJFYA0lWq4bY8mf5MuErTv0Nd
xa5+MEImnb2Xe3YR0r0l4ae6FFZooHKQWQtwvOBJgqcdUvlqyLaIn7oOX/yTSqWl
SHvTVLwYa5Gdyr6m51eZtr7sX3T2SY8mYxD2EjS2VMoyFK0K6Fot6Ju7Hq+Tg+35
tiZImEm3VU45YWEbq4gXBg8iaDliamOEErvmlIt7g8ejlckD77Z4Fy/fNmDmwCJg
bnzWTedq0sOTvzCgLzzuKXu/oasdjmWQL0SXr/FWByON5hqImgnUk209q/ZEWCqY
adZ61/PdWNdf+bTVHxnB+Ei5nnrPXBb7VD7fVXrI9mtV8FFjAiCIb8Q1U3gViKMy
+SQuedyJA5Nt0jR117HKbafWsylzeYE2GkqfLZZ0pGGSxeUU3NQpixhHIDC3gAv+
E6UjfKbv3mABUQfRQTy6Hu0TI28q6UalhzIq3JlChw5WFRADUqbLSoTyE7LUAiEq
/iO8rzIJV3OItGdEVOqfZhEZYqmdzubrHhonsanM3NPEcfRNWbIHJ6UxLBCpM423
LA8tyZOHox//1FTE9tZu88NcqzS5V2iopbsWrcTIAVKlJvwicMoW1V9MdtS1rplW
n41rgrC5Yf8b4NEBntY7tGuEjg7VEP8QROBPsYMjhiHPgK7bFR3zmmT/I7qX636L
HLRC8zLJpQmcxkZKTfqb4LYm8RP1B7surIgSbversLImg8plEmMrhQFNobLt0YvA
wGPNVTswuChLazkRh/eNtIC/KLI3jjn5eWrEqGk3BZjKWqEzZXMNS4bGjpsjkAFH
Yc6PC+M5gpi0Cz4iwphhZFG+CGX8epiTGCqy+jyssAUC95dLj3MXyeAvkU3hVP7M
yj46WgFu3ZJzLDBgfmUUA+ngpYn1k+iQzokqb6oSc+oR55IfoCD0R8VviUePqJyx
lFz9qEsrsQ+H4wYx+kYlDmj4ote5+4ZBB8XFRUu69xYCrwdsbEfdEWGzVbj7vCVl
Q1WuzBrdux47SjYwFHFAPZdtifWJ5YdD9y3d1dlqYqALEU8/W0+YYcZ+bvZ0YBx8
2o7Xl9SrUqcFpyoje0GtBKjPTOApNWu/dtSH8FB9oSJJTgl1E7ffwSidqMxRrbGc
RMR6f0GlTI+vYnonLhbqyRjts4FcVqr8UmmBDaImXEAn0TtyzivJokXpZIgUdS2V
THcTpMvx2ChSkHjYJtDKGTXFNB1qFOG6i3ouEUkdWPe5W74e4thI7sK2b/bYj/Oy
R+p2VwuO8NhhVU5Pa5P+RVmSYE6BbP4HOiI+ycBrh9Th+I0T9HbKNaheqzjnaRjx
Ua6C8b6IfCZKwJZ59tYlTsgKVgdT5pIKYqml16AnZgIZjM0L7T0kAjrs/GUQWJVK
XMcjUDQtemVzUHU1jNHhpY4d3u5IEwrmiXNMuXflT6THDvDHlOc9tqG1uyAr7R5r
e9vlQzvBf98fnVqFM3LEptqc8c+H5Zx5L5utvUANAjAk0TYyuX9qCTaRRadVQqwO
at57X7gXzyZNUFKnLwY5tw03Dy7dDHJzdr/+Bboej1ioR/wP5VNac3GnLh4foFlQ
oWbk0yybyERrWAq843UCE10Z5wIsbWMUztJn1wL4Y775O0cvIIOGUvxvQ7GdO/S4
X3n9zvZ1aU2Wjdx9BtzlBKtRnKMoDHmg5dSrWo5xLv+jwcuzAqjTAA4cfuZ689fV
jQeA8YLq0ANiUhEv1NMSYZH9wXudGcmkoU3cHQzQVxJBuGvwfoAelDeVGHDLBPcl
ENpKdJN2QinYzn7M/Fk6Wopt3mv05PRIGeyw/7BvGnKN5ZrzPAynp9ria0KlrtnB
KIuLwzuIFQIW568oga4sqWiMwnL+UnVfWCHD5iKAnUO8HjoCyBPIQuhju6EgJDTG
jMSAIUNxwFECBIV3dYeFD5dhc/0RlkRz1qyVrSpoSRdMLu7iDwfjkPav/xlk0YII
RI55nMlXcGPAS7mLDZoVa+P7sJu6A2fJWwUhTbtu9nzRCSWAFKGBXr4R22S5c3kC
cc80aYDePAVdCyqjEPjoun5ouACTIhjiPar22j2jIlxliB55WO9zks3Shcv2sx4b
p5QKjU3r598k9hqaROzlytWjhQEpKb5uW+OScWb4lhqa6tlyPDVjVSclbLD0ZYB7
XPqlCQ0gxUxsZldJEhgkPi/I6HpynxzJey3g6cNAdCsB1Iq1f4KSxJE/4yumPAlN
06d1+U05j5rwOSc5QvGTJHivXvwQZSybgHQSRIX2k+HK8DwFPkfCanbe50tDksc7
We/hb0OP9gs0Wbs3OyE/A5j/jLDoNQN6HnwStJWqsQgY7yf8wPVIwfkaVBkankb0
vagQFdg9OvusiuqyCSrzBYG1JgE11UMzsHixWkoxZLtmqsh8uX4d01Eru0oA3H6+
liMCauJbZQeTPHbmGVpSay//OeXaukAUHMEyt+wqDnaHI4kLWdLOE5dzM5fGMQic
PYQl8lCV1VusKCBLyRskCwcTJakEijfh2GoefAR8cNbjTCwPJ3bDu6UxJIBelRA9
s2IhUQozvYUVcPK35aOlpRGXlIsGJV9anTl4OexBNbJshRgHJEjDDENUkU5XTt8R
Y9gurXHr/i1HakNyFhRYy9hTwSQTzBKSX7/1HdEUFOtB4f+9W1xTfWc7VnoPETv/
AFRJxNKMOD6L2a2N2ZjfSq9Vg4SH14g5vCXt4pqXb9jLV6i8woY9kf/9SbuKbwtZ
wEZr3xMVLe7k351Cctzmh2dlnZxDqlW/Yef0KR0xhE95utJFfRJBb7xYyfqwqFgn
JlxEZFkJeq4hA7HfyAWY+wWdFHPS4sb3YfEmTubp2auvXXwlvDYIxDWYXXH/Tenj
gWtX46T/FWSArEpnvDZcKxTeoDhL1xh0zy30sEYltwAo2nxkvg3bPktJNWJZzCgY
QsPkbGa2110ceMX5AN8/pNGEAVPWQSjuFaxq28bkE9P/EBBRjARuP/Xize+aNST/
E4Q4lXNmvJrhCTHZKxyDtdqMwRO2jM1NnrIWJsJwo33PPL9iJwO0ju6HB/R4dHQ8
lw9GKcvZQo4OHnRFcBB4gOoljX/uBADSeOxW16FH2fQGneRPgVRSeMp1f1QSTQkq
nKxH9g8Ii9Ac5LiaGXKnURejqdEWPDC+NPZepbrKAQQLX6cy2sMyjgypj3XnWHk8
qGy/pRJTG0sYHIJOn6BGCxc15ZObbpNY6aJSkRqafvTY41hDdyzMBtlKZFjBfX/X
AOfijkzbr2or4JmfRkm2uhgorVN67c3kY7Kk2Bg1Rr8yri2ROlqnA3y8GlGTGWkq
tOs7e+jl7KYHq2XryG5tWvWFkel+KiXIKhXbWgTEaErpVfbBbprNPygLKklGetXg
Ys7Wuz0gRukt9Yh35I3bG9ozXVywFiUzJjYJfekQciS6D+04FgVEjuQa6gDNA87Q
Wa7VHqcnevHipZ5MzwUUtWOl5E7gw0/fk3ZXOPOIqWjLy3m9e06Ne5sECVdlnqSc
mwCnrMs9UPTvSyGezSJ9x7OxSfJ0Y+9DvBGgwx+OoLhG7z6vAgt7aENZ+YekHZXZ
Fr20E+1EvTLMlfXxljltOk6QblPiHnG9hnvQloxOUaZE9unBhTJeWpBFXMNnSztK
UYas0OArKUp5KxdrJmHU+Ag1GkhKwXpxkW2Y5+tcDPHnYHMduAWFUcqm4MBVdgHt
jOV4QKOEBfPfYDnuKQoFWIUqelS5Nyw+/rSSkb/NCR4d+hRDIdgluoMXRsBfNZo3
CmRYX+om+1Fe5OH758+BRsu22Ju6sc3BuZZEY3kMFGyfra1KrNj/rGCivK1Yjdiw
Tkq+YkVTUArAOyBKKeKXylpn2wak/yXhh88cXc8uHoFqgn25rlbrqP6UuPAyUjy0
GxkR30Ch8G+imMYSd2gPwQYdEYrlFfD+4QFD4Ta2hyaSs/I5IgQC1CCuJG6hTC7z
d6kBeIi/ec4UVUDM54oXDTTkbsR1DXQQ2oF7NsJdB0BPWDQozkdxOLYJZLcLvBaa
UPeusWMW06eYIIFVQFzDJL8PY4Z5yIxlk4+pS5zgtKT2D8I5AkIGt6B1QujLaBxM
sDaepePL7TbAC8KsMhA/1vGXsrTtrAP9jm/K16av1JE21dVDQuE87OQr7unl7NDg
2EtvINmKMZeZCZVXq/jzI0Q4S1xRH15NpajqoasTTxCVeaEmswqCreXJHyXDB98E
9m1TP4o3vN2Sw7TW9U6vGnjmK1hWmj00mzTTEN6X+33iVuJiXXctzNlVFzHY7SNt
wt2jQkJcl2ZIrMDRzP6LUs1wN8FfsdoKY/Z7P8qm+d5kijltTkblFjaNI4kAAi9y
P12qGtcrkDNyfGQgub1oxE+SLUwtLheMCGxCCDu2NZXCpG/5MdAw0VeRLartuLaQ
sihQHXRtDqUEhIz4jv89jCNla4r8jV7xWbLMHyShdI+SexOyWHYDuky7KRRC9cm+
+BR11Q/7C8sNvbXkgVPs+btQ8qGVtazVup+daepY3SIkOerqly7lnPV+7u0XFeMj
m73KVvj9o4TiISAW1u3IVJgn2Krr44KZJHG5koq+yDwylvqn+GMNfLcGNeQjq0lq
WtsQDkeQwS2ZBE9RXbFlearF37qnCVF9p6Lx4MLzaqrHw5ThrdPqriW4EghbLKnm
FQvPfoOvogaU+VzP8SDeDrZazV8I4nEzlcDRaBeOphFdhw2aOAfVmhKnDignyJu8
JoM6WrKapwUlsQHPI3OkcQrYOmd7Lb46qRrukwIm+BJ1W4zJxB9scFMYz2OOuTEQ
JlZcONYEfrcPYEoD2SYKIe107mcn/dBnAxCLlAly+lCvpTrlzBp32HDt70NLkMtO
QYUvrkEdZMa9fVI8eDJKfAdd/0l+T1pD6AlhHlIcQ1j021Z6auBurrGpeLuE2hCD
CbvsXrC/TiZKt/zxmhHek99U984YsjzpaN4UKjtLLq5TPUS5XUBLdeJL7w6JOYSE
G/rUs36GWk7D6Jg10T2zHHI7vKBZCqT8WC2YVKqcA5km+DClbrpBV1lmwtwsrRH9
fCZkxLZ3vcQtFwu7bBdISGRS7k+R6Ddwx0KxQXecRbxM/DmMf5h0Zuv9tSJPIDRm
6fNra2g8vshomyL0o/BFOFEeZdft+zjTiFESdIaGJy2UFXIMzH0B7jbgxBLLJt5/
qvmzzqAHyvOsHGoahw42xmBqCvbC7tqhDjU7YPD98Wl3lb1tAdWIbYRDSjyqXLi1
DP5T7S0TjzERPzMMjXEUQwp5PWkVIuXvuDhZ23wZ+MM6Kk8TW5rP12AX8H01xreS
`protect END_PROTECTED
