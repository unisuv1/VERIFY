`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o/9Ab2lwYgfiHM7YKsZhhSCRAbmgElWxSIfy6LUuT1rmAlKdXS3wD6M/JbjwBPtU
7x5LBwf5ky2l8Y+qzHxHU7q5vS76CUcDQ4LXHq+B1zTof+/UY2LnU3MM5SbHeW5y
CwtzN5GQaA1Lec2uHPjcCp2MRBvu9SCdRBnqGoA1h4w1niE4X+Vh2nc3gGO2KIwX
xtXITLcKdnXeznxwEB9ido1JNWaTdZv7GVh3l6NpcuhcO9hNcoRB5qG1B1juVAwi
q8KLnAbtg2aU8JOnfvPcq7YEGxWt42DdXaCmK2ga+twXafNBhjVsHUydk5a83Aol
OjFDivNCvTrp1x17OSCfeRYOpwYs3NuKiIqlby2iRMV/v3ZACZEDUao4Ss2k4NtB
S0WnAQhduH8IinPmkpMCsnbRTRcE/g9V9epOW/54ouylmWAtY0nU+lOpKUfyseFr
qPTmWx/dn9uUCxAdhOeG3jcSf8Fj5CRItRal852Y6T+gfzp9FZlpz4KG48vFrh37
7pzzQHYgb2P+fhiV8W4zouM1SUaO9sEVEg4taaspooYB+8PLCg7MiuE0KGix0Kl+
7IyQ55511OIhiN3mVYhVTyPtPU7b5fXpaIKKcK4M6ubMQUMJeYLkzvKsEMtoveEo
hih7ulgLDyBxt/smjf5tg3DjhSGvPVoemOj35DN1KxNPCsaRq6lVr5Ry7+frm5mO
ggwYG8zBprEUR81X38wh0u3v29SDjRquiJd0uQ0a76PZQNDuMREGjybkz/Es3+Uu
Izs0mCkBUUXD/aDSjCLRl8SXi+YVatXXeA6NB/nmQwvjQi2mZxc/t06yWsEm5rzF
1GsxcC3nkDbNOhsJ+MqvLOYDVrEeE+r9ZSkDlWF3v86zpLPZtITlkFOb8bkGhJzl
kK3EvmxTFKyPsfDy37vmfJ++BbfIDQZXwY8wmaLx46xJQLyBoOt+Xe0MlghcOKeT
/NybLiggR+xtli/3cJBz+Q+l+OQCf/+cxUiCkz9Zd0OL6o8PIKJLTpSyM/JMiIbB
cgykr+009VVjj4B0Q9nPaqOFQKaxly9RaVtYvdoVYQzC1OeGTCSihuj7OnHmcWtZ
D7NUngzldsQBaRYMx0YG7aMhVfoiBYSdcEnd3XXKHJgxdhYMGSJl0R9/ALDREQc1
7Z0aapW9nzUNveONQe0jb0npstEWGnFejgh7J6LsqGaBkwntkQTqEzgp9kUZr8M2
k+1RZKckREbz0eTqBcvWxxHWWPZ8B8Rg1lZayd/H3g2qILXELjxBD5oNMNUvydo2
e+25nrEOjakbHfg1yBXQxxT5L+G4wAMNXG2MuJTr5MoYQlIqiRW90DGvWvKqE+GJ
5IXddpJkeWGoz3x05kgKKWx/VpcRSlvE9gfZsrv6pJSQcYPk3LqKR9pPWKazlqga
R8PoVGZQ52rZkgjmI8FB0V+760WOzneNH+P+56WT59kzk3Yf8xttI1Kj7IuC4NG/
`protect END_PROTECTED
