`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
F0QHFAvKBaX9Yg7EMqYsVFBPP9QKePq8lpgvEqi5bkpfJytWUgBcjK1LqEY2l6sx
vz22Mho4dOmstr/ziZ6MtGSE1xqwuVkwZpZveewMjsvGNmQt9wBX6vCf7aceldbb
ywwdw20jQgs9jyWrHINswDGZyi0WJHcTUxScIEyq9mQO2Q4kRmCg4GIQ8AY0Dd0o
97m+bfMpzDLnpNtlJR5L1XXV/ifT780RdX7ztPR76x1Mch2VDsHAoHqfITO5WWR6
qYybqPwQmkabSCIClMbjiEGYRJCJaNjmX7NeaeHprqp/vLnL1wq0gyBzsZKn/eQ+
ePhQNeRLuNFi70YEUyf2U6fmvQJLITHv91R/IER3BUsMOYZ5D/Ts2ZRXibVpxDdT
2p2wmzP450BSpZHIeKHdR0ZO8YTWN6Zq61Qbefkj7XPyavOZlnFX1RDXtAflaTxJ
hZprvLCHYmsr9fDrAVxAc6GoTz6fwJ9nTSUyMZOPaQrpUrWLxom1gkfSLe39DelC
ac6IJyhH+jrPeKH1oj6yTFDID2GWyuVOg8MPV641S00j8MlT5OcnIc5OymhrrqXx
JL5M2v/L/YuWh+sFYPmVv+UWaiHGgZ261a6QYnnAlGagXwQLAdsywwDlsA/r/Ayt
wMz3g4GyAnrPN1FfakY7fBb1gB/xT01KqbGVTE42SIIj8AOyKKH21PC7jHfesE/W
sxG/I1Lutf+OnFeQovR/sHPXdVGHLbXJAzdJ3Ni3MAbsr/NCU0ZUQpNcFpcy1vQx
Isba+ocyLpGLTsZoOYp0dM/JycY9bHi05y6SmdUG/3LXcuSUGmvy+EmLJn7rWbLK
SA3X7nlmIa6h0lDPZzVnERNlBDfn58uqaiYihBpmIPquUxc/qtDzkRnC3c/35CDX
DMoCpeKzgkmGAaoaaRjfAwqlvyvPK6Bm7ed/IHO6VF5OIg9drPvt2+JZHr9mwFRu
DzyFBSs3Kovb2mGrdMFUpvH1jIkmg7ZvvzR6/a78iHJvM1vvyuyWW3VmMO/eWdWr
+isU0GBFtniH0bzKgz/LHucV/o6/NeVUsH9pTAdaaz1LOK9aVU+18kN+ez2ilTzG
o4BY+/XRV3ICBciC7U+yDVYjsCaN/oYPIQ6fKZpYGeoY2OSZzBh+cW6dUPfEVKBS
BQPwN7vqSkPdX9fxEA8JZW5U8ruqwGhkb+QcdXM1b7HKqJ1FFS5RiE9MDRJuPL3O
/1Z/nokGETRF7C/9XZfLb1fdLeG+rDZi0e9i6VPzrRbNhBKNKpsbQojdua59vfX2
KA2WAjF9SO1Q9UrHq1dnvkAwoIij7H+FgWZcj1tO6sTGmBNSsZodXJLg4uWpLJO5
R0Ge9SKnCeyYGTx9Lhg5A+e6NgM/cpmF7pNQ85vrfnRtA6NZkuNUe5btI2J49sYz
K8fnIwhfFX+KTzBZrtvKHzfJ4wulp6NwQBhEjHJ4Rex/S8WghFyq6L4GupPCNjAg
q07xRtoxXTSxbQfS1D/tpSXC0qNc3Hanu7dyeHWeH3HgxLlvXdePywDaCQaD4L/B
8J0Ec4teBYk3ircgx9tvdRW1cwOKA1prHy6W0oFOL4EKeaEr5klgTBwe01y+b9Tm
qpqBx/xEb3rj5STv7BDYQ/sJMnGV595uNecDYorahsbNOPomaQCB/TgHOQh85zmY
+6iyEaHpndLQO8m1Tjp2fgNZ/Icih16fCL3qx9/Fq9wqHY6/TSv4O7JhAaherRur
N4gH7nJKHxnLFeRaEhzqcJ/CgIPnCp8o1hkcjyjkMmOm5EfTr14PFLj61/yx3qE9
Q9NWcuUE+P5D5YkiiXpN6VG2FWh3qVxmWUG9UDbACjIV/qxWKJjDK3h9GYq2bdc6
E6nhOO4jvC2pq+77egqCx88E0PvkJ+sVGP2bL7UW0EGZm3Mr+hN1XdID0cZcLbrz
opyIPf6/3+M3nTB6Bu7WFvIdYoEMNbekG+u+VHFVCgT6GnW6qR60Rh2M1NEuQ1tV
U+mGBsY81Lobb7ViKVoFHQ+U5vqGVod07/WyTe0dlLL49tCyl0Drrw/HNRqGfJjT
fe/YQ0y3neEmq73wHmfwHQYc+b4EQYdGGfRHk8C1v8uWOijshknPPuBahlHwKIWI
d1L1OSikAGxle3dAsYt4bt0MruEpMOU9AElXcmNaKZ1tlM26RyVstOKgBykIKeG8
nICJYdYn7CyT5FwWK1XLklH96hGsX3xNyR+hjp/y2UUghF4mMz5W/jWJkivC9r/f
GYAIWFjM+JimiZIneZTXeoptqMoZrDbI3XPADQJQuVmxH15SjfOQVFpN7mP6U9//
79oXokOiBKdgpDbQyUz0CQWv9jupN26C1QC5ctfgX1o17a+/7TUlnY2rvqqGsP1u
LFSV4kP9y8nEUOHHqrshdw72clV+WOHTRDAhUsZz9/YRRMVoV+AllX1/Xj3Di7CO
yIf0A8gxdpM0NHYrG9QfgK5vzhfWZpnU6sh6j5Zxxzpc+TyAc7zNwzkrQaq9gZBh
+p9tc4OqrrfVXPjneMUVsWqHNW7icfTWWZ+Ido1k6gqxCe3qhTc5eOfnN7axGfl/
/KrtVjtcAcouxmGSjnnQh5PZcol0IQskstt3iwRKTlnYEVss2qqtbhAOgWPyj9x3
GqY/atCRLv2pnw9bmlFd96xXWWtiE9Obv2qt9IrnLzeFkN+Ow4TUa6SA7ihnHRsv
k7hLSYXEEuwCY7xNbgfHWny7MPhqOA33uv1NXF1/bclrZ7SnZIR/r/L3XUFC+hZs
RNEMuBdnRBpDMZi2ipRw5434XItFbeUUdwPD/2wRp3B0SFPAtuV/7tuAVRIjKdW3
pkk+EbsgV6jdOgthu40S/MOQfl0IpKs29W4qXfqpQ03FsECbvmRyKd/npOxBfUV1
G4XDf8Gu/1qvzlzlwH56fD7Pa0GHsV9yA2dSjOFS5tugr0N2SoyAEmf98ZDHeU1d
JEHqqT3M1YPzpW7fkGjZR8cEDvp24y6nCK2Ceco+n6s3MNQaIt03PwUA1daY9cyo
rV85sMRrVDD/tM5muwk8DeE9vxTaOPtyue6ul3iaJgxo6PmCQhD5kqxYDLUYv7C7
JakSK2gtl6K4Gw2RtsGfr1blZFTqKgWFsMkgktMr40cOThqqXttFUpUQoA2FJBG8
Yxj2jSCHIB8eV0PQfYXxXmnoUdRhR1IXTMufs7/rZPFIybJoygu4A6zIEKW9zMmj
2ON7GdnH8PqgHKxXEjVIGY73GXTl+gYr+eaOLDVnxCimMvisrKkOzkxPrfjUoW8j
iM/h6+5AHMSTjmRg20Ew1u7Io9xMfd/2zxBKK37WGXPQ6mdp0jR/gUOqBQLMylfY
C4dGd561A1d8FXrG8d4ZciV5zId2wyXOqCVlCq0Hg3WtOqnDgk7it28pVeqzShEl
5wBwtjOodWIYHgDM9Va6gLLnfHzRjR/Hdat5V2G9tke2+JewnN8R8hBFeQzbWWrl
Nsue4CMnFO0TM5eV6ToDEJOdi60kGp0F6ha4DgyEsjUesUkpkaN0oJPaMlgzIZ9b
CSaJA60eB4clvjr0HhPuovUErzYkrGKJq2JP2Rr4tWIiky3Mtl5DVKPXi147FT7U
PQnUaAdywZf7Xk4dIufbtFZ0gV4Y8mqtpeKSGgwe9F3XvYW1lROrRRATNWduQkID
3Gpn5510XmtaCqDHopnQFSPrtc4zce4HO32qbepjJPl4H73fHUbWiiIh0VaGwEdM
WxB1RYiW+MHkBAtTe+Uk0HI1pmkUDdWQhz/crTOrmAzte6v4EaIhI8HfTt5vVrZu
qzOJTxpM9MCfkaqw/P7ijsjwlvtjAWeu3f1s1Re0AiATDXPZo3msIDaXav4a409L
M3WgUVXsjgUVID6MaW/qWzTOtWsTCdOaQiUD6CPNfPscvx7Hr3rY73vp5lrwOmai
cBM0WP7kfRRgBNlzkbxVrYtGtwdbi8b3BuNALtqOh11tkkZZxtXInQg4sxHxqVuM
C1nNzrr3xaWeUjMelFgcJ/V4n+z35a+NYU5E9W46chdKGbD0RxBQDJGtU/fwD1/P
3utByexQCril8sYAs85rBxgh0ad5PyyQUF7XZqH1NrJAAKpHIA10qXKiFoOIDicr
/bUiPJAxga4InSwUIXGB9kTL8YFpWxqqYGMSAUOpIqcotEdZ5bv+UIbOFuI6G2Di
MKnvqyPTC9wt9/a82qQAn0q4GEAiDJDimoSaBztbAFcZvHaF7nGzMXT4YEattguU
w/15ELeWSDvHoo2h4qMlUsiR9ryQvznJlXtzl1evt2LK4JlD7XJR6ZGhWFFri/OA
JLYc1vs5IB/SE/5vrpP30Vs+XXUrMlcsbGikoJj+ztmbJ8QuenJKNLzkswfEIS12
e7O5swjsqW5jy+ibC0GpKEuBuwAM5o0YZR0nPk8sooWoi+wEYMctjpnFVEfU/YfC
ZPuJIuv06o/pexIVW0DXaU3Fq58zLoY330LqNFQMQxt1evl6O0ZjVv3JrgduzUQz
44rApVr5xHrqyr1DoJGzl6YBAkfFEaPGiVIif7iRA6vpmScZUTc9URWz5BLnFOPT
IjzIgCK4etRykBmcP9wnDjad1oZDf2aITmXRWcZitI3VFIWcLMh+rz21qdfTg4gh
M8nv30f+orzc/J0101Mcl/x/wZYB6ky1PRW8pqcQwIlXLos4b9AS3D1gS5lkg/xI
oRfg4Dt2SEsaaEtBlnKsYF5Gaa4J8s8yGE2DIxDbcx4qNYNpP0VL0AFFox/lu58J
BWhekx48+1mGOmJMlmT5yALTY22qLxuuMEya9lMwN6SATQWQ8jSca1mhsK9duOmJ
DVUUgbNxwKc78tgB1Jt0zi3ZC7eK+62DqsvVG1Z7p286uurLcRCEaUdudr7t6hiF
nEDiY2/iNmM8W167z+C3xawVF2a9wC5n8xpcW/jYVorodG706uiJRLzriUC1jlIG
Z4T+Z7c/svRaGUWEg5RvV8Lgzq6Qnsvr6pqY6AWrDytjSUwUojY2kNtIgxQJHQbO
9yLkLZFdBEfAlGuVR2nMSo4m6H7+TVv2F2WA8ZC+VnNxbfza5Pw4Nrr8uHtt0idi
kdx/7IZ8Pq4xZe7BdxWG8k5Nc8XDALjH1hcQXeydeVXYYMcFnJHOO6WmvNJJTrWN
d6+i+62Mu8aUwwKf65e3kEk8NO89NlGjUMNfEKEucURg2fARTlM5P0oJN1oVE3Bn
rTHqAFoYmVykQvKR0osmBK7dwWWk4FU4Cs5n9k2NXh7bMRhB7T+33oTK28OtpH6B
/5zz0f0u85Cek7k6yiD1zYpMLLnL8Rm6+n6TwvKe54GmsQgvz67q99TQ18d6Ru+Z
6qxDyPL+RbCa7rADwRKqj7PXeIyIuHwu4B1Hz6V3V85rtN+QxIi7xpKMPDexDf/u
EboFDHje0Y0qCXUrl2Vbt00CqExPce7i5Ki8zF9WdzZ9Nr+h/kLy9QyUZs5CkEzb
Q50YeCxefP5Xas0KEJhtvnLd4j5JgzpPHT6u7IzdIle4CrFkbQG2eq/Ern3lxMZg
vcz1rruyHC/24nel0uCcuimn0t5Gx++ob4L3msTITXkWMgwrSXC8PA66qJ5eWcdf
uYKOD8GRr4adFxuQCRA2aF7nttBAOaxb70YjgkU9afSa7TjG4GmQVgnDwQEDL4tI
RuNwqRMaUaGO7io9SsuLiO2Kkv03VfubhWGx4NU1jnxAVGRMGYRNFHor1dBqt2bL
CeAe9CbXsBVHfCYNNdOGzXIq1zd9xRb09+/WyaFUbZsNNqNYKDhX7RbXux7L0Z+x
ihC9TmesYg0t8kIMHHQ4w75rL8pQcjsBxwddofNVHehHldN1btST/Lk5ZHiwLnla
27AQN7t1ng+EQj8riwbMJAzV0juZb6yUH6W+oGQoMUkFVTvYVOaAri5H2f/d/haG
+uX2/MNIQ5c44ePKhWQ92mYph3NeosLG0zxNrOua4wFbo6aN6kzXSgcZtAaEBRUB
qdDEtqxMxXhHZ/p+VcpMX1lpNKBYuugkFWOTzcyfG5K5JE7iGJUJrvWdkkkUlTU6
lZWFGlNTXRS8w+1EsoLlqchwqr4/TjGhdL5L/s3y7phQtGaPyERZQvP/YWpZf8VO
IbNT2zdlsccSXjRTewGed6Ky+f5QovKaa+vY0ogLeOW9Md7NUC5v/xqbPQe5OL/S
16rlEgUWkLFpoGG8S1FdRKeVYxiOOvYgqNz820rLr0s/3/Q+eRMOek4L6mPG438t
BwPEFrMvEmFfUPwRBfm9z+1wXlZtJmqsQ7+P9p77ukwsc+i9SOwBu4XK8JInSV26
eJA2m6A8gSH9uSXqG3Swv0Vzj1FYoYHxteNw8mBWHiIvZ8py5WGMEEuCaOzJ3QXV
vbhDgr6KeY+KepC11U0XPhNi7G/lncwrU+gZqkpF0yISEokn8l/xVU/Jh7NWhuci
Cho9n2Xl6LeJj+nW433uZXwqQAOEv/Glb7IyShuBuhKL1ORweu5bOfQ454+ZkZQL
LzKiYHoCo2ze0sUlUzB2n8ktKlTDHOxalixu6oGPkP+slS+S7++BVIUbSlfaJkWu
Vc8FRjQSF1rRcL3OJ2Y9pEvFYWPwxIGhJ8WJCgQ1X0QiqqcaEfeVYqSGcZ0RNBQr
WwnpBFKsz+RWrSr7YcKD6B+8Au+uLbJUbHRF5EdjttdY7zIHpS/Lt6xARI8hA4IJ
XeBhDVORbUzV9YlXwPTVgHhHnVL6D7DsgZFM9ogMd+7CUqwphGIyCsPyzAcPgZTm
3OefSgxfieHdmbcryxtP7NgDhazRLlXiiPj+oNhriu/P07x23jwFxWxbXH5ilN4z
kxH+lwWCGNRMlHBefCMNVn/4LkO/5u7u7l421ppaAp2wyQEGtRRI0WAQ7yK5BDKU
aO0DaK8Er4RjDrAToRPwkniJJEmgTKQI3m6CCLfdnmreSy3Gaj8k8YfD1T2jZtzG
E0FN2Q1PA8ucs+/xpa5+nCGYw3THyugBvxsbo2RWGkqUkryTBb1Qaa7xYw74sW+S
rnMeq29g61S7axV45fF3c6yE93SQQgeMz/L/aOuDmuAbUgldIHZOzcpMNthckbWy
JkTIew4qH8vwc1A5LoXe7DkDG0BaNFHuOZZKrEQUm8bNPKLhsGntWyAuRGHmJswX
AkuxKFrG/rTRCFrecMC6VbO3leEyMFMCd9KOrU9M0j4brpwUohi7EruqXIqJ3Myv
AUTL4Sh9awF/6iDywNWrd8thur/GiumNhZQ4PoqzZTeXqR1w/HWC7xxP9+fdrT2n
aqXpkiDzSdYnWNP67j0+gOM286orqViVsTXskxuraQ4etkeBQ4rgiieS6KrqmmAb
zC0njqHKJpL7TKaJKucHlO1JDjtP156PTw6H1kwWrYYXHNS2E7FYlpbkoc+lPuBp
9dAUuinBYh9UUxGdh19QoVcTjtDMw9K40n1lvdnNV15oCC0C+mehhdOOD6mjRrNr
HC0k3aywS6FRhjyQxpg64+WvT/DaqbZtRt2Kuaa/SpE3KKMGEXFqnbqid+7S7uE5
2Dn2ET/JQq633rMzkib5mVGefVnVvwy9fZ6ewjScjvi3ceqSHGXLgdanEQ7mV8Si
5dYhUXZtGpvoGrtdpgDjsBy4dHFL6qQ9hbJ6gyBJK6yUxz0SxTzGP0SJ7r3gyUNG
HBRDsvOgjs65HvgyumXLcklQSFxB+GPO/yH9tdvlnPDm+umTth4vidPfuWWOkdz7
OW5ob32sjrlCv5NRaX2NxVe7wDlKtNUmbXEDsGk8RZsYOTJ2jtUG83RgwP6IKDxF
53aAEYJBHEjSicY2oknA58AQNjUOzbO5WKzBgO0IHO9mP6zEP3EJftPt7r8mjUMv
lvlNoFuhdzKmRjKtukbVl+9qh8TqwDK/FAe30tDMXepOzh4epY2VWEjeAIBWpwe7
XoYywf+yF9R0h1pV3ZDtrtHFOXreLJC39TBrOaN6Vill/efukVbUhVUo8iFmGyJa
PGlC3zRcfgLkWh/gtdl/hnKjykVb9VOv3cjeVKHwSYW4D6bfHlN5snp0HDEx6PjA
Z0MtvFsIHDO9ferKQdFFcFz+Skj7mQtPkJacPDKGYls5spawAKwDRrAh4NsnRiPV
uta9Wfb9A47WSbtWTCnOquhD9r7YVZrItj/NF282ucj3IOG873mB/aGdb3UO7Nky
iyjIidg9gINvSLT9JGA2nIjVyw2i330frtIDesv6x91F2Hyg1a43Y2+KmrICKdoN
3FsiNDwvR/EuVnlBPG3vjYD6F8ticHoFvaWgrknLrfsUhpVwmHtCBCEYcDBjp/3Q
G01WMXFD4I6BEKhd9UlauhMouur2WtvQ6IYoam3pmiSBL2njbc/qv5H2KyykBmg7
vQ0ZKbWRRea4n5W2JGKC6hpvsIxSvc00b94y+JsCo9iqZsq+ahaZ3vJZ4bm/97lG
ZeZA3Y+wEdQW4cGducg23NAPNxwhqyR8ChN0L2Wd6wzhi2sbE0plrrbjpzF7Vp/U
K/hB5Mi9ChFa1UnbkV2FHnKYwzGPSlWXr4dquYk4s+Oo6o9uCCbm1kUJvGPNfiBh
Fz7lyXxH92xFTDAj5FhJ8QT4eom1Hxx02yr/jdPDR/mCIPkrNpUAFqKDExbek0Dy
x7G37yfJWgMOKPVbEnrOUhTj/P7sINaVFquA2b6XgcpSNWHqMUrAy3LdSyHuPjY9
Hhx/RDBdJx9hkHmrxnQD07efykwZPlsGjy4tSmzyAs2gcMtmzPzWswYCr11VAx5A
xbBGWLLrPnQV0CKU+88Sb1waAzsmIi4GCh4AYIrFmBqrQKzlAo/s5JtFN2985Yo7
EUK/gy2M62OkYHx70QnpdoTuyaoYPxN2XZz55X7sa+svBMTJuiPU1shz+X0rialn
II8TbWzGR0rNF4xGKhw6q6YL9W3OxazyWfpZDvbDuBeuRXQkBfM33uGY+0KixAZg
D2ho3ECuElB+EQYUaZttVb0w4cNz9AMO2yEOJmrJJPjzKfoSpg1/ZnC3AYjI9zQN
s7ZQwVVCkNqR0vExtCwYZ/YhzVDuEqIwu274hO+9Q1ePsoDtKIpJ6XNl3D0lET/C
M/DtMROKBF0n4XHFC/sTC82+Zec/KwrcXJWvfUowXTwj9catoQ8oGN0dcUasyG9u
71wcm1Dm+9nGQQz0eaHRIxy0S/5OANtFHYSCtA5IdC22zxF/DPrd3hmJgObAhzjl
TVWHP+3e2icrzILvWcTfcIRwUA66Yj3ry/QnVyInYDbb2oNjkIRNbD8jS5qFoHmt
uPxfGTd83SbBhgz/GZsATfhoXTtvdyZQWtiPEIn9a4QrzLbNQB2vnfiDft9SB5TG
dbw3Xa2wd1fGWJN++GprALITQXdBRDpSChLd1IRtwyXSRQdcEWhBkqpvzLzhO3wv
rrerIajnmLh9JmSkn5+RWs38IhYwk7z0pRxPSboI0UK94rjUcsqpnEOCqyDKMl8w
tWquNWl97fvcJ0VHBpRuUTsn6N1Y1M/C2ccgXc+yjvSwRbefF43ZQ8tKXV/7MyVi
Im1tcaMp78yqiahT0V6EoV4l5vyczqQfgGjGK48abV9XmVEg24LzQ4Scz38w8kp8
sDw6vWox/mlL6uiS7T2E4FhoD8rhY/LH9kzG2MOFxjU4uU8VLlZ91aD5g+oec110
kCti23XM3kYFtp8LnLabHBvUKzUUmPBvkhBE/FJXgBCqSDETrs+tMKzMoa7ussum
T3xtn5g1bBnEka/GHqehAPakG1OcgppuIG7uKMrjTJU33AvIa/Zcxht2ZG/krZbi
LbuudvEhzX+Z+aQmL0Wh5jf8PSeaJihFmyt/+5Kd0Dal/dxpxsaBi2Eg1gXCkQak
BFL11Dfl2fsgNZzRUMTuyZ+YLCfOJ9IXFe7Gm1QS4vw+vKo/VdDG2iWXYNBNN7GC
VdIX1KIUZGZZf7mwcs0BU2ruDk2uwXTD7UKLi2UBZcd2GQ8gxSro7iv2nIDYCtts
zzTlsTVOyANgfmTrTXGs/0eFKo0VFbHdseqYsET7w22EvnBkoM7bEEt49+ofEt7d
ZSpkLwvRC4jILW2rS/j3tSe+fdPTNMB8PxUJOjIsJjdOeLjrF2hOi8FYlhULJweu
V3yHZwaBLauZOAcrToa1HOt9p+jwRkIK7T0JjVxVKSpOWBnMkPimF36ed0+19USo
SOVlWxn3ApocmANiK9MbIGo0ciYxH7EVXqH3loqF0zv+I8pGcyVpS46+hQKCayso
vx+KAzJmtqnJj0MR1H7+pvGuV7kgGfR1z//2R0jRBS8U5DDC1CQ5KGrv5rQ1lbxc
OaPpGIQJslF+8NU4vyNqMt6kaVHPPjYJtj7iTuUOb2l0MkQXqrLFGDWmlDJL1NmB
hQN/cr9fhVPfltgs3+Ldak91lcN8+mXa5HKf8GZXCPtjARarJAcAMobPur3VjR40
2+TKwmag7HzQvtaMF6y3RqKnwayXAFCM+hdCQLAKPXvtzc8b6+7mFf8bROWTDyc0
qNbC4AvkNFwFff/d6eJI5IkmFA4kqzC08/dPQKO3iHzQWzzRjNvfJtvqg5OPM4o3
lJpBJlS4uUh1AHXyjzXM+XT9V8o9KygAGWYs4LpgqKApr65yYXcBKr+U21qqeK7X
v8rljNL/wS+UYH4SH5j666rX6JXCkxXzfCE3aLZ+YTf2nwfp+inUDl5ePfRJa3Lf
xd/zFGmfaqnD+opEq5kzy1WrcI/wZvryUTPMIwub61VmXQ8ngYYWnG1w0FbR9yTV
eCEKgN7QhWabuESoGT36Ufn69LXqEDq4+v6ymVwdUajLAR4qMP5y1xf+7vlJFLi8
hiQE6SfGTAdG/FSiRA86i2a5ILGd8M+Ns7h2zJpTpBxo0T8dgdy+C1plpt3lK2Ip
OYi8oc2CtWyNLHMWd1HKQT25gA5GiRr8hhO2O6vEH1+xyOd+lcUnVunyOs+ZoC8V
r9/2qHioudKnrLhmv6DQ64CrXUryJATw7Y+m/2sTm1rf3VZu837KJH8HihrrlmYo
GgtHewAn9NmCI+IiWVAs9HTWxlI1AVF5eDORiCE3QNL+igbMovsPnk6HmR5BbaKg
qJQboo72ZdDTTBbWMjC4TNwv7Z+tMH51xBTB+pw7YnRp6bcpQQfLPNoO/CpLhMjT
gxH3KghSyzydLyIxSDGrOC3th7JVR00qEf9FzDJdJVE9lPF57OXzgs2RQemaGkwG
/VzCFwV1bML/0c8Hoer1ONfOza40W7FFTc3hRNNOXLHGEv6ovpagUFOhelkHaG8x
Ut/Yt11PJdPLVDtEcfHJpipeTK76WOWaio8CueRoHQurh7AeFT5X616xF/htBG8K
vjo5ttdDlt3Xh3WLlgSKaAxRcw+CdZUCZOPL+i9pmkHybu25OvzZa9guDwzyqMsC
TS8G7A8iLYCnItpeU5rW5oudm/MX1oB5VfiPyuh8CLh3LmAOg7VAkgG3a5UFJe1S
WNzOcdsFPrdbb+R58WyBkhWlMM0IgM2shnJylvgQTq+OQx2ArClvb4cPnkm5OqGU
ccIR6kAeD3ad2q/N0Ya1ITb0eYkpDomMOOgif+1w/Iri6cMof4jW/RlJLwmEI97+
+L6U+uDHzITMOOW00qOg11A7pfyJbzKEfBphMfeAGpkoBbAfgDJhv0OIHGv5Dw50
JUg03VOt5ek3aEbc2UStMGF2KY0Y9jVyPud8SypbpW0GU4F5uIKGPxqyLLnY9cBu
6JARQU6h9qWsEG0B/NJFyCATfB5E/8nztiAJZtUeUBzMXJhHGTH0mJaQLZjNsAXC
KjZqztXYTX5uG+Tj71QWModQ0X/1misdASm5WSSIRqPBKTpNG7WQx8lCJDN9ZHEj
6N6khAdIW73xQcP2B5i0Sad3huemJnDUA2x+kFGUokQJnTgF3Uv+myIpbiicr8Lo
bGuLNADmhOu7y7IAiA7cy72IRcW7C/M/7ZHXQzzhkMnHSUuCHsLcdQcxYW4n9avn
rLFVFq+gmUBgxRgtYkway9XBXfeUtDCBNKx0Fugo6M8TD6HFO2j1B2+a/o/puO6m
gi2GJoCDbPtBOYAEgKVKf8uOpeWJb5jUIC89Vihfyd1PkoWdVD5MWyy14QYDWqpg
7SogbDgICpTzsp+LIdw5IG/IFr3yAy+VKzOICn445MVA1Fokq1CZRGBrC1mhRqqy
/RNGtxtHSFTp/CZcmx60ySahiVSnzyTCQYT0U+hIl8+qypvR4azeoWaRtJc9H5dQ
6GExOrWn2KKlai0vrr0+T2HFTaJZ/0LlqK3X0zZLph3CxGfERc3xbGHQzv0Ek6Jo
pYp00MovL5/nvgBSvrU2NfbiUH9d/aMadOk9nfct4kOvGMqjRZnVoVFMvn/vnVGx
SWbWpZBWKAUcWIM9TenI2WExy7PzPh7CKMp6FVVdUdTSO05h7i9BBXr5jacuRnLK
4mqCyFuIAIB1Tleh9MPsT3GBNWz6cy+N3QV5ocgBJ6RjQURIbVYlfBj4z+2Y+4Rd
VYQNWar/WjjJYIylf5RZiMPxWNeP4F4kIyfXUGFGnffaHwWi+Ez5Al39GbdVF1nS
RM1EX5cH/Nv21/H8kFrZQbBAt3r4kza7S+A7pUEKSiRxE8n1dpzBd6W5ddHjXdQU
aeAT7LRUsa+pFbPYrIgvQwblgH0HsHHnNS+lniEgqJE5VTEDFcyRaYmkad6hx6W1
Xuy13Lf7t1v+daJOPR0vudfB4VjO23lZngax+WsMAvGG9ZKdAqkXQCLmQhNmHZbd
D/8pWzHt3ZTIPCtZu9NJqsEHtCelIxCaiiCic4UI2gNLkunu/fEWNLgnFF1J02UE
9CCBgA1ozIZ2C9RTqPwrTslltWlGeT9QQooi0PZmVXhiPY5nxLHzTtrJOdE6tjS5
NwJq1Wu+O1THo+Os6x4GcI+KssZ9hG0q7+wXyQ/IyiwO9qbOq0hm69DBrlPm/r68
ROLsDL+TdVolvYOkDiEoLPpV0izKiTR8EC7/ps9OYEpMC+8j4vHhm9oS8EqoYRJK
246WuQgVifTNazwb7S8E5pHxIt1QJ9k8O7V0c9ZvAAv7jbgrHvB7ceJTlSf7QUKr
KcpZmxMojpQfeAoAlkFCfv1lbT1EYM2GtgfCfVc+8TV65ERf6M8agDo9N/II21I3
SwK5YwOcMU+nd6eNV8eS7pJtqFZBjZcXEMf/C1gDuJok+udwYZUm8v8UpLL6uEhM
ETlRo99TaTvWZbplFwt0Oee5MROYbeK0EWc/Usm7lcOs+L4gadti4p2APfKC0nIC
4xW+1s57ysIUGnXr7fURlimY0XntaWVXE1n4RCI7tgsA+YGS7+32AGoBrpmw9aUl
R/eCTspO4K4Kg14BUeaiioi8uySIbuLV1MPRUdvrTUTgKhXHgyv9LscYFKpOC8VV
/au/ggPdoH/1br8jVAebiA==
`protect END_PROTECTED
