`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s55+bw2aQyspdPvT4c0tsQoOe8nF+NxpBzbbv7x6hHAlCzUPoOdK7h6HIsfbZ3bp
0s94HcJjBYmZTOkc1APqap7EfFC/FV4SoP3TJP6+PmPiNP2oy2eS90/m3Bv9y8mK
RPvYRCgE5fq+EJM0f9zZ/PNahCOlS96Zg1T7DCtLGkJILs2udOBszx2l78G0O0ie
kHa27LuRW9V8QArgkcw1Wg==
`protect END_PROTECTED
