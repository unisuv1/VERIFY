`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QjlNhNCQmoJyKk3heNr2bW6m6PegUOhN/AiaH4hJa1pfycumeoIEhvOs96QE5rT5
C/d5JEN28zLAcN3gR192GNxFZAWl8dbj0xjSQQ36UBaOdxNj3rVdzJwe+Hqf8Scj
S8MRLcvZgYIA6Enj4vCcmOd3vM2ZRzhoEHEYtMThGtd+r7zZ/tRW6PflhY8aXEOP
yUv+cbJAfQCDHM8eJcduYrBMUmoxAjopFnAKX8x44EhEbDmKh++HlE2sG1Ck3x12
YjqOLugKHb2FSoC6MQgOMKJxdhyXcB+ZNalt/yN0O4ZCUzp38titEjaHgevS9iYp
2H0vwQatuXdmtDYQgu5Yd/hGo++B/VvyIz2v/j5Tx6Uu04512JMgbkLTfNflRvWc
AWpgl6PrDl4SJTWrKN7jaC4Rz3fKPdg/pt5yUiJ+NLeDNbKh3OY2tF1oHuRovKM/
vhSWpx8rBGZfmuA6UFQ5uEJ7v+S5ecRuP3fSSkYFWmWxELUJc3zSzuaVDa5zOq1N
9CAdHvQ0cJKOe35pxYlGZDVn2hJZjR4OOniDQTrex63b7GqqdQ7Hicg/39CDx1wk
hhfZuNUaAp/cnAtfCQwpWaTCsERiZPY/00nb3BCBxGRznSciFEjTJG9Crubj4piU
V7aIeWOKBaFSuMwXAqOq8AlnVTq5ynmfiOyOsALEII4upTGBOpQn3+myzp2aPM3k
eb4E9LZapzRqLQCRxGxDtNYbCC9TxVe8wRFNTbUIBWBe8Iyo4dZyGGrNh/IOLeM3
LcYBF03ClN5uq+NA11IFtqbd708A3K18hV68lLUmYjb5LI4fc8q9FIm+Lz7fEKqZ
9xIuDdltsPSKQJYztlNcEa/604NJMyOE/1vX0z8FiHS6ytpXgQMWbvIkbxKSxnU2
pCWwEUYSK1MEx2ul/vxQfcy3UVvkjNWxkOR01aj9rXlTQevEHCHHozoLhBUtcIQg
JczeuGx83VVVVY4fuvbHGUhnUoGz3xwzXjPhc3ZL6CGS1Usn19mGjaF+Fmyig7p0
6SDZlfleXim7wqvhVaYvOtZQ5f2NHFDTHrWYWK25egKlSdhlSmkRLD6T1cIfeDw3
tbQtYMePYJ9UbNrOcVugX/YKDKgjUJwfuoYG5lfEwP90hMJ2lBxVjDuIKpjKQsnD
m2r7dI4pUs8eu9cbK++Xuy9W5X9PpWIAXST7Rx6DaqkJoAmZXcnCrFTAUIaUQjbI
FPPfX+POfpjfkrbCLScMVLKOjSX2WuyO/DXljJf8GR/9PlDxv7Y3TOCSlAgcvO7n
oWYTWTgoGeM5tjnyeAZzLzSeiaJ9k3KuZiVlyqI9tBmgLS1wXWjhGp24IYLtZvbw
E5MRlBnY0K9OeuJYW1/mTecCVFdZqQ9TSGh63z0qnkPqN7JGLZmJLaSFnaq+MQCY
UnwHJZClQZzKUpuH1ZL+o55p1wpjR02Ymz5I4NlfCy11FA6sj5PSaDnjMXaLXxhH
Zs4jr9SN2emY4kGUbrBfdIuWWzfIj3JMXEHw4Dp5a72npCr4TKPW4sgvXbqXSG+E
FETMKDMDjKYI19sCxAfoIqlI4H/OpRWqTSpZUdB8ufbt69ewPOyPgu4Ci3sO+/Z3
oWu3ht8u8s/egTeZnUl3j9i6aw5bPexJvXTpTRIjETGzlhqtAp5U+R4IWTkji6x0
0Gf5wB0j0x1X0wNzxKuGPST7+s3NawJYfX0o0an6s5USdW6lkreJXVYEoBYy5lk3
llIn3r/rfsJn5XTSxDKxruHQew4iHfvfim6BjvqN+mXieuBRxyXHmIxmhWWx0p+E
Q/qalqTWUgHNCgmzvmaklKxUv/JXxL98JqYNW8Ez/RtcQ6YF0Pt7yuM/IWonM1ki
zfLbJpJkLWcUk00xNdspocRDmHMKHDbd3qNbyDN5jk7uBNkwAYwyKhLfItVJVegx
STksQ/AKGbevsHoX0kHQRBijpa6e7Xz6a2Ggyewy/isZgHKbCXgw+RN/8qvGcZUT
/YMV3t4iMpSmuvDyQi0i1BjNTgA4/LBUkT3qOO9HcnqJSGRtTafpXujZW99+Yvuc
pBk0gzUxphVffcUOwpCo4O2j1JGC0NJVEDSfWGoSXywuLfnSg7afPHaO7L/pH+hd
mcW2nNqMo6kCQW2xdIXPXx/2B0k+JhWPPXaNaVI7zZJ4Nq4K9HYuS+pYw6vtI9Pw
QQ1NpAtyqPd2KWBcKJkC17f4D/qLRrg/4C4da0/HDhrj/MKgbKgootwzE41g3vad
hrcG7EOapyp0f8DMJgwZKgdS3aGFNKljr358nKNRBcEl2Eu9m6FXL5XJTEZJji1M
21GhX/eiRJw2GuARt8uW0sQXxhgHH8BSDd7FFhljqUqUJkT+YK07zAVdPPaArbD+
zvfriiOvA9G8/R7ruKpxSR8+f7Es35RdoC+bwOzLlHj5sTvbukk7Itg8G0To+lqz
mVpMOichBL47nkIJy9cr+1SXO1mZWE4A7g+CVHnj4P2ZHWEbWv2EWagb1K87CU53
KIDjL13CTz5iDFEUzq1BwkX8+//lR2JCjSFJ7u3kbKSWdAAHbmdtPFOh4SD0s+sY
6URUlEVqSBXW2LXA4rZOQryjKN+mDthAOOwrrjYflXIngDK+yOticeL7rpgVFtzq
Iuv6l5RutYzPiawrq++Ak8jA838YeERIynJwLpwWxOy22yTh+KwbMO+uZNaSwVKi
UrQ0+2r6N2o7mpBTI3J2vUkgRBR2rJl/FaE3BMgh023tBsQdi4SH33vMy7grDGyE
V9oXLNjsNE7CImJC4/aKi38/MK9bv0bydLlZ3CSoEWO4OzrmT1CFFYiwREovk7+m
LOSHXkuzTk6d/3tUjCj3LR/aAIboT2hFIiaEo5MEAS1Fl6CHtlwMf8/g4u+rZyDE
OJ43lfNlxlzwk7jRI0fqV5JowKkTh/umxDJJLhNQ/ViHd3dKdWRTOFRDL/XpAm1m
KKCplHBvHrznsJL03K20R6CBiIe2vRfm9FENhPrD5n9w5INsm4dm/qFujHEEuPfs
GbiFSMCGm3TOjQ4cpcVALA49EnHLEO5BhRqdf/ZVqQjKuxJfrYzHewOBJwYQyYfp
R5tIQBgO8zBdLDGlxF0UX6uNG6gUkolC6rW1oJ0vtn87GPgZUHVpA+ei92iNk5/8
jh2PxpILkIX3WjKOhcvAI3FqIYHnQhmWLYiTMQUKR9+GkYXKkU4aU7xBrrDDeOnO
bxRkJolf3uHvTljidw/eTOOkPIl0PhW+RubwkrN4E0Gm3QT1bXu9AxidbYF9PyO/
p2H7c7Nl9DkSWQfkyWYBH+taTlnJLRXsOF1Q3UR19Vm9e0NwJZG3eVJe19yCCwdT
0RgHEnJ9Mav4DAZ7mECj/Z0jQ1lXPGILkMr4GKlJ6Y5QZuqsp9imaFmaN+TogXE2
TO7F7xE3Zmr7U0Pki/pf0mb5EQtkLhL1PrIUlY13H7WWbiiyQ/2XM/iSfaX4lVKb
I4SS695GaS9H+dsWyP+5cNEtaYJ3mIiAppOXcwOfF/PbXVqTCTNZPqmKWpr1Dkgt
YSyP2HvxEq9EfhNraspjvA8QbbT7fw5jwvq5X2ud9ZwynPLqP7Ht7DTsGeEeRi3M
ydIhvPEtvrLxNOlgfOhtpmX9pxmMI8G2FTuhIFaYxAoEwOPxOnb4Sm8VxErer72J
V3Ka0OyIfiG09yD7N7DZvA==
`protect END_PROTECTED
