`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CnciDfxRVz9dTqfjOq+hoPII6TxwX6KTiJPiGMylcuE5tiwWaKRAc8ABLKQPyfvL
jy0QFOfUuKGSKjhqFKxL3LfZHyshNxQhwGGgqzCnbph3tMaSVMiAx1bXsbSswLWz
6hJ3irU/wRSX6ZEmbs/UJImH5S15mY5c+qsbHlYebFFS0YXrKM48ao143gV0J2QR
PG8Jkvpin/Am/vleeAZDAgaJKyuF0FhQZywtsylVKxdoOu5OQ/hEhBxB6QZ5kmYU
reboZQiJ8ki3Hu67kF8py2W/geHu6scqV7hqtCgai0jNrxYUGkzLcJH1RNnc+Am8
mGkf/SmyrPywNH+W7CDEqlPN9TFrlGej3E1rczhMHv/BJQI0yg5+4f0fcT+Mn2lU
fV9pAiMdF/WtWmC0xvZKAZS19g+qkTrCYNaBX/WYGGPzCK4yDSy4OEj0gyCg/AxE
+qhWtqeV2GM6lhQ6w9xbpG8JfGRvrxC6J6kztaUyibLI7HaGAGancBWTKQWdiGAJ
G8LRlNMEUQm2gLE4VNdMHq3v5fA8K+JUScWqgpN3ci9ThZQGcTl7ZASspGIHr+8j
Q7U1e51y8a8c9oR+kkxrLSqkgBzGXu1pAtNRxt5vAoT2JTYJd3YmM9pwQrxHFRtr
Jis5YWEn6jhz4d2b2CYI0PyRlX4V2RsKiaWXuitwAMfF1dDoZK4uR197+13cdB4v
CxExfvCM7TDwDBFTd+iLRAevx4PYlXvCoT0J4w52NTUtQc2/qnYbqGfmYLH1yU3k
Lp5zYnK5kc1haudK/Uxz1Q9GMEmIxdA1hW4Gh41LhySHoY4CjS4j6ynHdXHAB38t
mCx1LTVGokpk0y8tX8VDRq8i19MF74ncyGwL73vHoq2AZs1Fuc4LPfuI2pMQTCGS
EwkObSwBPQdBT6ytZE6tZK2+nvlq0Dv/u/ZidecBNxueNjSMrC+wVL/64K0tiMWT
dCDVcwjxB/DUbtYQMqnnV4uYFpYxHBfAulKC7RQEmGUW659xtZ5mUzItTeo4YNi7
KQRPAGAnb09aa2EKPKWj2VJB3M3OSdvVUvG97yg/7hzGHMlwvpFx3CZbZQfA3dJw
JejMOVn4SojIdnMmZp2WeNMRq7pwRqfPVg2JEqCz8ykr2eP5nvR0eU0Fu3jQsKH6
4S+rYOK+qv1EJEMyDN6LicQXw8CtZpr74h3uyfK4l+r1jHEXukV+XjZ5WKxvgsJx
an6MJf5MR5QcU2UBQzBVDEoo7UZpPcqi5o4vLC/qDlbdM9ZqxkUeDtTkr5/9GgBY
dNXTFeIkuUzk0SfaOZiQKotHrQpHnSeTyKajHoSqj0Cb6M1qXk4ME1XDkv3oTXmb
6CDWAIkiQ3slPlkNmvSMqn7425lJXVvU+9807sHXGBlODBxggI1wnJcrwvjFCOif
PW0InYirHs+LtM2UnwC61AiprfAk8piyzbjTIZp/OMJBU3S6CuZXWgsHEi3JQQdh
rq9kj+sil9oXfXh+f7fUT22l/j7oGa+hmChRylXprIJvcqOySZ81TNegJDoWGxid
ducT0DDQH4oRT4qNiR9zA0Am1Zog8hJmKhJmtkjwxeayF247YwlJrvokaLdCh+9A
2jeeaaRLIVOy5FniDaCmiTjLP0ZTrDbqL4c+joVrHbWOg3WkKlEI8dFwgSGJ+XQd
NRWCG9vcIdpO00aTbTt/MLp15X3Go968fZk02lRaIul7Uv55vlYHHQDJeOgkmEY9
IT/fOQbsLWeSXb6IbiWj8rGNCIaeQ4sbwms6zF4ADHWzWZ9a2Bl9c2tHd3pYItBO
XacE+j9Q9fMTpTwrq+mlTvtf1AVcSACYAffYdd6S6GjgOSNiO8jDYXiyDgAYyFtn
p2AWMNo0BIfT1rATtW/+LyJG///qreNZFXpZlDOBaNeQmKYJFvilm0hmxU2kTykS
uxmpCo30xTMTSV/WLaoEi3WOabbJU44uilItlrp9gyZ5nHcRroEuE3UYLH514oIG
uVsF8/oQlLww+H23sLNDltvDPFIqHsuZjCvs/qC6391FImnUSbHPyF+8oE/IZrW1
1RBC3hRW8TiJ2iOpeeyy1rFPHwE7wxv/5MevZTSKOXmpkwHsFoXZ/xiMF21AQFjf
e8EXAlg8F82uCkSlPpdduA==
`protect END_PROTECTED
