`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
RQyfiZN16c32RS9S88h6oE8HSAhEiqMGiNYIOau3VQL4KVgtTf2CkoAjCnOU2mKa
C/2pzeb/M7mK63a55vyTpgkBWHkHLbaYJ6Mx28LQEOYCfHEd9pDTG2d2skWVNJSR
cIOV29vbm7+nwV4k7lPeEgUDxklBbcg5JN6LHJbzPX7dNUMOADAzul37ZohN39eO
uRyw+Wp5fMC/pr1RMD/Ecw0o2ir/21AxQFfLjTihDlsyjwtAcBtT2ge4MFrhCoKw
v81wA/j5JpNXDSH4aCkzRwP8dNUrw9/jjtdXEXIGRcXm7Wpl6AumQ9s50lG/n3Fx
dG/pcn2aJOWNrsuCjmnGpFWFekSIfhJQxALSxeMRGUQ/AK3G/0Mwoma1Rwu88NM+
P+92PLutqTBXzoOa3zd1ZWxOs5rrWTZXp+761X0AvcmtqMzk0AyuWqlUELNqeMyW
`protect END_PROTECTED
