`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nCqJ9orcw93dnckDCwLD5cSz/ArcNIimEIdrsiZRxgh5itQRl6BC+GROrrddjp+r
w5e0VXGu3fM1vbrkGKBjlwAnnlFsgzby1fbwBXzhl5/etyD1hvPU4J6noFB/PCOK
FkIMmrV0CS1e87Xb3qgtvPJkBUWqAcdS7F7bdab/LYldy2gs54lIa6C9HLRJkSwK
vSA0DgYtceh1/OvP6GCaomy56IYAYoX43Gy/zjis4Y1TrkCdzxCL1Ejmie7AFSYA
so3VfpYtsQBsx9o6moxrfVJjbRc7f46Hf7JsdHxEawsfcom2fx5RsgzMcWjx0JK5
nCp02FYWhuZaPQdx++zbJaq4+bN4z0LzhycwigShIELFRihdaWHE28f/2gqyEWbV
qokVRMSHH0LqCmEKmR/wYVWAKW4FDhAjavBQPCgNkLRqYpupbpnzxtKtEqV+U5SP
IFKkZu8nkCh31a+WfBrcKlTnoosukmVktOpIvg/GrY7SvGAlpFzB8x4T8g5WAby6
sdDJqyWd/3OufhFsxF1XsS1zk2yY4Yd4SQB0aN2MZcsm7sr82hvSEYS78+21yTHa
N/+8H7q7H7CIMcRR0mz/NRFlcyrA1azeotTFCEdy1JoIF0YLhMVrIF6FS9PrF2/F
3PeUOo3EpR5ie2sn7FaUBPPutwhY6ugCFgyT0rndISmUwl18XhZOPBMOV2TeHB08
rUXSZRj3LyhuqMctnlJhkvG/6XFsl4GW0tUWxxRWvDTwbwfBvYjk3KV2qni43W9x
G5K8+BaeAzXBPpmJMvBNx1uRhiycoIslU5eLOsTDCT9Uo/NoTqlfBi4EK8RlG6jY
0nDOmDHktjCRzFtxu/Mxi3y1GyIvzVgCsgqo0Ex8rW/VRIWSQw1Ph+udFpp7IsIw
mlYQFwK47jmCCU1MoypZsRKhZFVcDu795RL8PRV4cdbM4qgDSi6HSmK8a5rxtLxZ
M/yu0u3B0rjVNypMKXqXer80nVD+W+lmRPJrTUe97ib48943NxSZR/EvR9LPRfvh
i5CDrdJOEjC+s6zn0CuZAHIvizIwOyFRh5W/wJpDo7h9wU2YgoIdepg7puWJu2CA
7/ldKz9m9ZscVwM/zdmiRoDXxL2VLxubQkrCigBkPuZZ6uosr6JYd8uey9G0k3dm
QNMSupH319t2mobq+DWAz+zix/AV4NhsJO5CpK2ca8jC9gOBvTOs06JUL5x0Eu+S
I1OleAaBfc0lk4h6+VIp8aVvE9ct8EpYn3f+hrSfTy0UoWiDZIo47W4VVXWzpyoX
Q6T2ZgmWnVyh+BX1l/MlCiXL4sbDrZtIG+WJsstsjBgdX7fcb36P3FxFvuDpgdCM
u1apSLVrDlIwT/lTVDo3YcPTDLZ894vu7OqTPMF8qXHVtiZfx6fR3t62X16AVNSO
348kmL+ZjRGUjsgm/FFF2F2G4XavhEP00ViOnCHuXLns0IYpIcacsLlfpLjNUVeK
xuRzcgAetdsEXBC/VcsA7RrdnyJOvnXrmRcMRqZdgas8GzJP3wnsWe0E/TVG33Bz
kKeyahExw+TWHZrl6DTdj39/qEa9gAa8CYKiYfHaiEc=
`protect END_PROTECTED
