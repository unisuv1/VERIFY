`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BkSyDt2Lcjm9VOGGSmOWPrY+HEyHBLV1RXqaUin0u7HHQOWi9Tu+QD7cXD42zlWw
SwOVruOD8fRJEhKnReOoAX23BOlAUJlE3nVBuGM95cHOMKo+IJU0eSuovURh7vH8
TPGFOy27ICf34fUmL5XsV22BZMiF82CmUhfu2fDlIn1oWpcCCMTYWahQbcvObfFu
bcLk5PNqkZGHJ++TnQ0fzJ1rwWuCiXBime0sRAeLGr09up0oXzgn0ObYREvxjovK
wRplYewLUeBaevVlqXQET9zvbCjwmkzSieQAHTELqqOvMN8lMVIJMHuKX4MruDUT
Lp7VDfeNYB2ZCB6y9sE7MNcuRrCPX5HkSBI+FosUMpvQQgCsnBiCuaTS9Ud1AJG2
cW8fhFjoMlXtI1Lh5g8VTJr8/trz18eLrK32muuavfekGD7dcvJ2tp9feKn/J2pF
mhlSkSo7VA2H2KMspKoKirG9SKuIb+FM2v7SJJDcaRQPO8Mfy66g8n72XFEzG4tD
lN9o24grKBK22pJZ5Wo1ZdR7NZsep+8u8s23CnXg4ADhKEGDNZJWTa/O3qk1Y/kQ
PblCG1v7DcDJzqolFaFMBmeXCO5lw0wQR54rOc0RN5Kbsm62pC+vN4HYtdKH1IZS
nexkhgrmKUsDEpjYN/ZhFgEg6VuBceWh1YRHMH8x62VvBTRLDUxnWeamAqINObl5
nD/vuK3jO1snBR+JtOiLce+llbY/NgKNzKJhjBiMdxcP6botgQn6ZII1f0x1uA9O
8QyMPfC7gHo8lydr4km8WsLhwYy0DfAGWK1IREmFW3kc8eVh7II52p9KraRi/PnP
UMcraqTci+sD06lj6Von6jXe+YRrZ7bcTdvPwTk0KznJgT1E2wdUJqolAB9/r7+G
z19EbQEMgpUbYE5fi+h2GayKh+GNHDS5SwDdk8VKdp+Kak6suoCYzMa7TOun9Tvx
beci3xcBmQ7TxFA+3h+SD3/LZcSSb7/ZoAlEjS5cZig41H4Q9DTeyMJyLQ9kc6oN
bv0yfd9yFsZaxlLXomUEUZVxraMFEu+jWwSu9cP/W1LzfUXTp2WJU+mfSvUU5lQH
RCkLRz5jrLN1PDaOnYnr21PQH4TQ9WEhHAbm6aZK4gZJD7ljFwDrfu+VCQ2z++kp
T+pP2KXDUyCXTOQ251tmLr0wMWo/JpB4HjRUMJdYPjsteQmdWyvvQ2FkRIfujYm2
zvh5QPsf0qTlVNLMjfNnYytqwUL2F4RdhyM6KQdPKIsAKf/8gPCKz+FyadqMC7LC
sHyNCRXhbmbMIckz9XyrQU7BHwLUZCP96MeOfffnDKQWEdvVspGqANaCKfNpswWW
d/cQMLOD2QUr4+9Bb1h+VF9fqzrTCbMv8ifV08KSSrc9I0EPTaehcOIQgpb4q1e+
XG218GZzUZKE9JYJV69MjjgS8ArhQ7sN2/l1Vg/scjOlBq4XnL+U16Y1s7E3TqS1
BiD8Az6Bfix5yEi0a1cNFnjr9vPmRaABGr6OiwrqjZ1WPsmhhoXahBrS1y+C/Afw
kH4Hw27Q18BeQV6SBKzBpl42YYcuVGXJvvBvKhSSuQM=
`protect END_PROTECTED
