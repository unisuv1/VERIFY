`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
nabmIfQVznOdIrl0lOfDN0FLBD3xAgXCF5TushOXzszWIEgtZCCFXH5J2geKI1zr
nTJHFt/nr7gMo/llVryUXtqGGtGCM63OZ0G+t/DYBUVmjRMeWvZxDIFP1SZhvErq
CU8eYGwZg4eSkXYfAAHCWXqSZfvLB4ono+DKocZ/sbzccIHh+n2c7e6JyGn8mcZG
Ezet283ZKH7O/ubfE6i/xKc/lYBBQ6Q5lNQWhOokvvoUYQoXYaT7rUmnEWFnFtob
KBH+mH439agXdLB5upQo86lFuivNT7+uZ0Eplaw34yOhHwK47AU898avztOvt3NA
o+vr1CFzM6zzlTidxb36KAsf2pKvFF2T0O1zIztplZLYFbaj1+lsOIxtaGtu5TpP
MIBQ60Et+P5EIPK5vKig98f5QYAVzamfkYZf7V5+hI75zABioT0Q/6njWHDsj4wn
gfDfTBvwmRyjmzHuFKtU32vPjz+1E8XY7CbrAh452H7FCuLCr9mLvRd7CVW+SEW8
7bJcjIwWCnuz+jPa+8Zx+gH+Pf3HnT/RQEteBaJ+HKVdYzbU4o6YhHBD0eHxt6Iw
J9LcuiiSskEMfOJxM7diM8TdfinPv1yWDzYGSRoYQh3fs8mok66DYgmcrM90/M1l
SPjs8wKAXHg7Fh4X+7dy910nQwD7lDJW/+8YvfD8z1mEjyaI8RqGtqa0IY9ymaGn
UqthfrjnU6DeYieas786N7//OjALVb1ZNGgPaUUNmmtq9owwtabUlL/uqNYUG2X+
w62GaCv6dMymJSwbeMsRtw0LKJAuE3ofRaemVRE47p7P2u9kQGWLLvvIX9ZvArV5
hv7z7whGbFSumI7unOIjMRtcUOmPLW/QHvNaLt3vqOIlRW77BzHHxTIODIn6ls7y
9gEjyWc54daGsLHJD2LVRYbWk+XfSm24yCeINO7nPzHw25xBBGkyjgfwcPZeXeRK
QXZrs79JLe9BuVpVvutjsxBGa1yuDL1YNucMdQ5N/exu4FsOHBfImgABG24svWdV
VPUmwib0OiVTpR57l/2HEsOrK5Kl7jLnezbH/N1V/pMCsYyDlDslSAAyVs4y14UR
1x3Ees5/bIxNcuxOfA/7KMIcDiVx+ztoSZ5fWHNbhfjvcjCt9wkfZFsLkoH2a1fD
bKWoEvGjM1ViHiBOXUj4M2Ijizwe7DuE2zkHmf/FhFKPGsjp3Zr7GfQHLs8d3afF
YVynT7ui1a3BS+2XI3f9zMma3h2jpO6fb6X7NjoI1b+SkDhJPnkHPgPk63iQhC0X
HyjkXBdgTjI8GrBieI2lFFOyvI1IcrOcZMMxxfSNtSdckY9wmTmwpIo/n22CUGOF
31Mhb6g/nHMKUukJJ60wELuLb+4m/T0s3kbxtHn3tAardM0Iz0n7F1qZrNVumC1B
Yz/WHfn+6+AkyFX2wQXzAQRQHT/qYhwmR13BR/x2kPcaGk6ed0mU2P0nq379hUPC
AnskDzqAeYm1wKK1+/tx+UT2XLICwduea0eAco7fKYjnu4cbLZVI+tcaH1lBWeId
nyP0qceI8aID6aZMECVLPjtqTvq90OW/mO8rNtvwefU=
`protect END_PROTECTED
