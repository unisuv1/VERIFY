`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4psQdQst0IHUP1cSlMiJsBAG+2mEncJ9oYOPxGQpOzjO/wwuLFkC6lY+pw6TQGcx
OKAIeHl/pbwql9hC0jOJEMH+ohaF+4wlAVs70EZb6zVRoNlvBE0VYQoG8JP2sx6+
vHn7uwcWmKZdwn7RPQT7wxQdND8Hhf0kxARlqWpTJCVa8j1ET6pXgpIN5cA6nE0Q
PGC2N0+DiJ2FMeS87j8uJmC5e8kygbXNY5L1cMHJlQLJD3C8hw4x03FsVFw7N/2f
JNTSzILnD88dQRNzwFfv3HM2s077V0I4HenyBSTWU5+ykRj15ATcdc8eHFX7NhNp
ts5h1Vd+jZTIuGaFPT2ju8dAVJ2SX4srTKoGzEgSH8v6s7XCSi5+E6kCHKZmcy5l
kGe/upl1mkHSU2n4zXtDrX6VF2IULoiDKsEU/YU7Ragg8/b+LAldsmW9NLooBVg9
cIbn/p/pP5pvOE/lRxqSJrCNgKlGgUE2TyTotjEQXzzP6nir6ussZj8pNghQojEG
h8tBpdwybCXJbS+RIDT+59JAaIFGmHac8p+3prghCMCClKlzeI0vzXdhiw4JdeJr
MISkYmc4HN1xrEh+NRxlqiPGbcSB3eT1mcPXF1mEVDRmKVtC72HtBvlrozp+UPJR
qGMhw6wR1MDiO8KxaUzk3EvP0RyfIQoHl7QakNVkvlPtpGzZZMwg+Fo/ewJV4gN4
SIFU695WR1XcyWs+VhsstKUOClGFS3DPRfQRctPFviwmwsY8Z1wCKYITs47EJ6yN
74OJwrFONR59J5ApmzKZzb6P0/kS0qEJZXsYKMnt4MSlP8sRTdQF94gHFsS8AGmA
ReTtfcYm0LSW1/Z06rAx1I2Fz5/OuCxsm6ANABra4awOONgIeLZuwsozG3Bcpap1
evI/deMH1/nUNJ10HZTS9X5x70JjtGbBU0S9AGO0KAi7U6rhU0C9hVl/fPsVtPtH
usbLVlEGeLZezkKGSLU7I2y8rqWgsmNFFtRUBkgxyWmiMkSdncDDdS/Up42uS3+Z
GDbPU67k+89qaRWeX8D3NvLZiNv79O44h1G88dBjm877he7EY21OTEDpAQQJw1S+
HElygLo5Y1V3g1zq36u43GZub2lk+RwmT/iqDiImUuUfoYa2+5zekVCa8meiWU2u
ImX0PAuICeNIJrSDNS9AU/ArGgUmdMnQ/UnpDbgtIBw2eDEa8oTBkXIIoJV5d0x4
Y/nGu1mfNppOSN1Rw3tud1AoAgAQE5K5W3MW87V3yvTwnXhqBW5vtpdEzhstTJNE
063omm3GvDY/9v7kj5n2Y+uDja/XK+TfDNeHlPnra90yFymG8IxMOHOfLu0HVmmO
f2XWR/FW4Utf2iQt9jBoZ+F1SCBV5MD/oddSfylXuVjeaZtME8cMQ8yWnPx38WGm
P63MnBNrwVYLiR+noagB/rPUFT53rUfvV9jyJzkZFnamhwdrgSPoxMpMOpdTbc5J
8NcE8g0WJzvIgycu+qICQ47IAsAkrv30GSsyf8+HWQ4FCCeDVthzWxw9pfwENc5J
vOyBcVmA56a1lG2rf7yhjx5gC0dl6Q+K4ME7DG+kDwn1JD2Ok4rr3vQYY45SZ6mO
gxWPa4/vtyltKdR/RdQXpOaXlkqhbIYfjOxH7Xv20WNanFa1ygv9iNZ/8XO/+OxP
7YOdixbqf2aXodrQwvH6PChdaTWrp5i2rHjgVuCj/yM2BLgWQ8Ix/CvQUJcnK9QM
JOc2jIPaH+Xc0cXQv/uNkJBSLzEN5YyuHSGEVamjjbCvH7CZ/AuOWHfQ1/HvDTuo
U2SBWUPvEIpmZ2QSi/Hnh7Kxoc8MwIijuI7l9217/dp9HVdSaedI7J9JJ+IHyJg8
jnRmvC9wYLRm3AshQqEsbdoKEFc4ZrzkwQPI6j099C5u+7TD+EglOi1ATtrEc7hV
7iTX5jX/9AY2kp7kdZCoS+bJwa2Cqe5cIImSJyJ6CSgYGg4x5l732JYwCvhQK43O
VUNrnistb6Jz75OPwGFHHVwpvHQuvjkgInBT2pD6xjZG7wTtVCQ27RVUgw+QjDf2
R01dWJAqXWvj0rhtOiAyNm5VrodyhFugpdsds3QAOgNsB/bU+H8eK7LxXJJQTMzd
7ViVLBG1JmFF480tG9/Fuvy6K3IqGe7TLWxmGeB2bv8OmoEPzTFQapkeR4AU/LXe
irgT72VIX80RmRFdtd7mquCt0SO7/2BP1+VfWBmfXl9sZEPuCnqy1HXt50DTIbwS
G7/rMEViujVs2XL5Do2Yg6oMl6oHBBcCaYov1nLKJ2QYYBm1LGnE3PzPMl/AICoy
a5cXSlPD6K1/8jrLrSGseL46foeMj4pEOt6JUUKr51ms3KVShfOBYOP3lOkp1bAM
Gt9Z9/QCWHhpAnZNBA/GN1mL5QZIDP+WS5zC0Zg+4z0UPdQAwO0bxXgikM0baDGx
rLoNMch1XYz07/gyr/ozv00BGAeorxQhQ/l37nVKyeK9tNZ8SWvUnK+0ff/dIXi4
O8iosBaASmuNqGHl1gQe+pYScQMDxv388H/GkDwf+wuj8BSwkAJcAP8pBZK8bzL5
u+XYXzPrKlaNG7otRszbnoJqA8eTK/cWya4U6OGLsMioopFtwYm1N3hoPMYjRY/J
pXxFYv8JSljFf+Ue+8JGlvLRRQ05P8xE3ekEhgqrpS8FufCkIFkDyb4037yaHIVv
5FhL3f+MEEE/+BWx1QBZxRZ3QK1/s7z3rRSyWSJPfxwV19WWXPN7agAJ4/OgH8iz
BbDIhX2Pwa/pW/zgqoqRZLHljQEd1F8AgdtmXfvlkSn3CiV12NYKNmNdTjZoDX+H
3x6kKhm2ok17rN4hui6UOgM2OMpVI+gc0Ti58P38a2Jxw/uEbG/VkUxjN1MXfhVF
tq4FpSbBeWubkbxxKe2uHMm7k1rcyIecMTFNQdlbmpGkfg5wDvgM2UcBWjv4quSF
5Y3XGQZ0Curyz+uGLtG6eX9V1Tbb4NCTg670Z5J7z20ZEBifYYuprxEdmGIqwd8e
91iiaLyTdgJ1WdCPn8DuneNcz8uSknrsOaAdxsCSoHliFdPW/6nlGbK3upQOl4l3
RUVX9wiV1cF9NblZmrWoJ7p6l3Qd0/BJ8xcrVk0EkhxJ66+0EX/Q2MTD2o57p437
GFmYFQQU7K1EQpoyrHwmGFgsRlrvePKogBHte+b4J6hoXysQ61+nGbRTYpTR1Rsd
rK09Zkmx1av8GSTepVnK1hHD6LvD7kZpwFaiiwdTqd0JKgdsdeCdYwkH/Euj7qil
hwC4VBOmeoM8i8XdCud3nLq0Ue0rMqamiaW4mKfBRQWkigtj7gw0KK2APDm2hIFJ
1+vZTT9MiOfr5Q6YGZzjMZcmq2fLkoZcQFwdamNRAtUYzxq61mZjlU0NNKwJqxza
Ncvi6qoNE7GP3vMxMFR2YiR/yTd/DKwoZz4nH2ggqOqmsLvgmACk4auwm/rpfrzu
/WP3u7MQnFIxevHrI8mpvMMEY7UBwFeESDFOeIzo6enr0UdaRUnf97NvWEXIwZlS
hZ6mLdHEAwkqcTC9zdzGFJPmC8dedAlEx0kEDIC8QjPXsJfBdVSQz2eiHWqCkaMO
DltZmuZiHlKMSQAQRkByxW/lAY4Z2GdLZkJXt1JIhruAVCmmOg0RZ15UVGnpJ7d/
Ymf0bR561GWG24nRbT+nfA10eNLngX8KAyhvpcZsOvmt6Zn7y708bJxyyOmX1cnE
2crX7H3/U7yBCaqsPqTtqQ==
`protect END_PROTECTED
