`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Wr9/PmVCvsOc03s6p7xZeYMCtRBoY0E9cBvMatUtWl9WWamhljg94DRT0s3FgES/
ZnqNtOVyJpcA/1NBV6Fiq6I17vwLssnoDIYjS/pz9MNfbQqiL/iQVVfwoHaIxiw1
2rKjGPms6Xf23gAKbgZpyrv7YYQ24BiOTVDaFASHbkpDH+XpgjQJgm0FbVyduZex
9G/BNRjoL4EdWzA4olScv58DJoiZJ2DivYSKtKWgviTdglUXnAwjJNESV8dJtewy
wFh9Gfb6CO9pKGmkXP7gAj7IdpUiMhu7w7qMmnbCdnqQfyhshbGtE8r4HtDPIGVh
7wdwwLIz7zVGY71xXV4iBGBS9/gbkYqwhXk1f9oWWjbnVEJ/y9KcQe6EryT62ms4
h9nrLhHyUZlKcaTpbH01JhXHH7RMU9ob1iaprj4DdERwTRpLGoGyrwZivEwL6XWv
+ZLLiQV4FKxDVzTgvP4Axg==
`protect END_PROTECTED
