`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gUEnTpk17/6+n2kS5ed+BPWPrmkT6z9BvYqAJqUskoxuiIViDlZhlnItgvShSBB2
sSt6m1WoxWn+8PKnTBzeRjtJqdPAqEOqBi7WU5NZwKgpNZvACAmKbrj6a113SBNF
FCp62ppFsubI9rLIYfVico4clYZCDBixqNESaA63XgzEi5SofhOfpOHJ0Yl8aGNF
Gml7VtWPgQw49ceTbRTS4ZcuKaoUjftfo+0z/etuT2N1Ld/Tpit5wYaXVcD6PoVp
k5IzxEnkqKV2wQ4Msq87E1CC+Rx4gp8pMJEkT3xkoe5MaKMHVVWichB9yruFvDMs
Pn48pMQaWs2F+RwCTNSFdGUzoT4HVbFlMXxUoMeYc7jgiTU8yWgw1oRM3eNwz07C
Ano/q9eZ+iYqDDtKZ/b1lbjxqP323Mgjpbzm/jvg8M71zWq122dWjhNhWXY5JFMR
v+WVBP7osj2N+Ndd9jUX0+jXuwRWUWgeNLKbd3gs+GUvNPKglkMEIqv9as3/EJ08
2Y6ta/AYZQ9pTV7ta3Ulo4LJ2WnouUigNNbT2eVXA6LQryEKJgk/DRaIReOvItkw
nN5LUKBSkErEz2xVuSDqNDFQL8q4i/GWe43B9jYabwe7NP9dV56BOFe+M0DxMFYs
HCvJh4dwzdDpTSMTLCAEGHOMqn3JFUHyqBtHsb6ow1NKeeSjvt9qm9S8LVr2gQ9V
+9HJguHb9Q/rykozHMEINnUjmcyI4GSAYIS8/1LPIeeGuOPpZEhpuIZ77DBm8+GY
6gk8lbTYpp7vi4l5vYdNA3Pl33BSP113CK7clp9Php3bwKy/wC8QX/u0NeGrss+1
iM/IBHMl2n0wv86A4tFLUTSNpuoUv+PY/R8e8s7kkum0cpuS9hk8Y9masmAeocHq
IIttTs3U69kQXx7wYcuewzBjLCIi3am8CWPA8HLZmM7s9DnSKEmpgk47nN/hGCUh
KDCfQmyZaSDO0/ijGRyinWIhRqrmIX1murkV/LFNZBrA4QEMF5scLYfVZoqZ9HlS
QnTeNbjnDF0915PS5VQoGzWUVycsV7hmVgmVL6cBdv43tHrHU8u6XECfrPH/iNxw
VEfAXxZp996MQS51tVfN88QskXYOIsfrmQkOQ/I63Q9fyAMzycy1H9Db9RBWN6En
hOVJ+fuHeZz6UpydhgR/CgChLMitSz3w7u0TyfviSdTQQxcg+4DP8DZzqMG7z3Lj
Gfuu2G1m2SmvVKGyLpZfmNC+kEkXWQzPk4glRY5GpjqdVMz9sUF//AGcj8CdEiLs
3xeAh8Jab5nGrrSCInpVG5UvB9TrctmJYvTN8HcfwAdGC5BRDsYjDy3kAur78OYn
MZDN4S6jnlnT4g7+v3cUY6alB5l26+ordbt3uYrvYjgfqFU9u66bk/UobFzAC62R
xfCJrLIeuSWrQMZLzb7BCPWaLGw/qcUX0YNZ1PNzDZJrGLuvqGhqIyh6vP91/IAF
3lhlVyQBvejVw5ekUtvPBNP0rnVE4Toj+oUxqWxy4t3Hib4/NuHJU0u7tNe+dV4w
5mHqqw22MyM1db/1hSJ0E0IL5goDndDG4IKptewiF1qRXzxLTjfxLIjg6LGk7nzJ
92+9Q+U9xeFN7cSHIdsDofqkcdaNmo/9Zf/qWd6VT3a1crH5Kwk3goyuvE9LaPht
uYgjdNvKnVpBltYP97cQKXmDk0r9iJTYMzNRjiAZL5Ot5hj/JZHfD7m2ACp9HhJy
Sz9x5p2/ieUkSxVNoVzLHBOmGUfu1bpUo8mMNtiM2ajIN7Wv90GkJhjH0bN0h45M
+sXklIDLLp2cfoITZvr2g62LeJWLpW/48tSEj0xmzZ74eLIVHOe/L4f7QTrCCXhn
5/Y5275JlBgiaki88XMlQZfSXa1W7UqCt49kz6SgKmRslPMxwlS+99OXrvl3nJnb
e8VbrxdPvAnOOxSvKQ9wacTG364QmqTP4TnrkcBos7wQSMmxKjyzjapOhtpRRMgt
e5a8zVHfKgaVtUhBQFxmS7Gquf2ex2qV1dUvsU0cF92Yff9Pqp+Q+hwhah1L/d4R
9pGUXTRkx6G7rhhxCiKSyi2TdQkEZLfG3TJLKZWRvfsgl3gwuV2595CPrCogpeAI
2cTi6tf1C6xSI7tqHohmSDAdCe8fys9k68fI/1VMHOq5la7YK4z2T/CO6wCqMtw7
I6OQPfaUQ7q5UI+z9lvVcKnYN9xgB3033uc5G2BQM3m8wUolxf4QtUSRMiYHgOLA
VfYj36Dig2m/i90sAUgsFMKVUFoyzvhqzY1JppPP0tEr0+2QxizsFraGPvH68Wnz
AOgrZ6MiuntRezDtnaL5S6Sar94cEvW9Qye/KJtZGh0SSAOr+D9aqYpOh8b/3Em2
Dib7f7KN+hMb+ep+dRE8fRQnVy7KJ5Irdl+coZWU8NhyVoQV6+mg1F3Qq1jG1Jo+
hnRz8HgMl2uQFlMKgiF7vrF74AbW6sM2u+jpxKF3wbiSRabIrhFLyRufxhtTTQjK
cBugrDEcPmQ3LBp+5BufmvjhtyYxLKgLVzEPZo+ZyUT+PYgJzlL7L60x0l7OTnH2
7NXmor0wepR7xw246rzHz2y19SEwYvrwUA6xyt4ZE7HlvUq3C2CwjEiZZumYO6fU
LDiWcyqpp5541z6Ck0J7NXSnIs0i1ekPZgsZhC7VO8+caKYs5BmD4Cj4ixe9ESkp
w9MmsZLJX6eALolPDd0vh62f8QQXRtJ0Fh/L3EQVUUDxpHFnE81y99L7PeIeeFgt
yo5kdQ5QQnzwgRMxLOTCWmghov4JTH2CfmnpCID6FNw61KdMkxNhhI6YRCyy9oha
SlCZu0awEpwqxSiMkyPAFTdLYj2t71kzaU+SfLWEoUFf46nNY8XsDIG6JJeDxIQB
0RrWCcAeORaCsmL+v2abks/CyoXIoc/G/9eH59e/vbjwFPwxe2KSBSbHy+IbKR52
pPAP3w1JK4Wxg1iuDcLoS+gplXSyQ6Iqsbu9l3rhUn6tbZE2d/e+UnISqCnkAGP/
1wEI/5jBYy4315nyz6EBOUnXBJR0dQaQABZ7oM1M+KQSHZw1uQ3uwWri4zfL5cFU
3dQzeV9cccpoZul5+AClEyxbpQBqLFaCW8RoVKZ+yPerweJmHyRofys4YXWJi0wR
JcVBhmDx4G1u5uHSe5ESDm+0TxBjqEtOEigq08BGTAE+jPOKqmQ63hn/H5EpxZui
eNSZEPBQ6a/BIwu1wVudsYzStiXbVB/TuZR+Ta++wJgDTntta7gGhB0+aJGRi+in
S4EItC0vFAGRpVCgKDWr/Ln5RacIlEuyooEZcy2hwpE0/pxOi94T3Zt8XoMqF79/
lPqsSsA/ybHvTUxVui1txXN3PIrd8QnwPE3a/agl/Mci4UA+aQUeK5EG173P2EfN
bbGw6sHWuqWFpAB2kY5+X00DpHBgNE2rN7LS2md06TmGodewGtFJqt3+uEweQkjx
B++Om4XwXIX4bnzyBGankkkNpuydiSdsIwnzNRv+HSwiaMZl3rXcXuJehowz2w3D
9M7EuyMbXvq20OQs6gh7KqXlifWspr4HxVO+AjJ2Sydw+AGAj55BGNFShHoyUEQg
TQtAQrKQURe3F8IG3DcyG5lnAOukAkZd1BprguTqhmLwLPMYNDV/h3YW6hoqtgqr
ZPYP95U9fvQF4xQ3OauZc/2bMq+GJ8pkKGGyx6QO0x9yGfFXcC0zBo2qw9BjdFPr
yIXqCNfHLdnk1GHoMaE0IA==
`protect END_PROTECTED
