`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z5QRzFXRCWORFiVxqo8OeUgm/pKoJFLx6dEQaMMiNqNlhp1h5lueIQGFibg1XOv0
tW6s0OsF6ZxKmzzdMOaCaSRx2tJvzXYoF+ufUsy7MxWhZ97werzyzNQmX0z1AAZn
YQkBfPo6lor6tfbOk9lDJ65vWGTHaXTKywlwGg7Ybk15T+bpxrQEapnIkPHjcXOH
mjzz7kitxo+kIZUZfPnK2Phe4dPsSbYWXqqswS/Mg2riUpNf3lkVyUE1qlXYxJTN
mSK64Y3wrUxQiNCYUjhG5VZiehHYJ41auv4ZJSq8wyIPBCJfViURzsyJMTTQ1Fa6
Cc0jcFGAQggLbS+3BfG9R6ipRxoWCBMGEaF0vw1uLfDTbOckao7+BpJC3pt5jFSk
K/sag7O2c91ihChG/JmB5eFw8Q63shIBKjgucP31kTwfusQlxGA4GkueOWcFdTwr
BDmjzjguR4h9tSNADCruq/c2ofkXSTkkF6BmWSygcwEyglADXTqEYNJwvqtfMfh/
pdbKJ1kJ2GGnQyX1WebsYScFfw6tVmKhA4Woezy2CtsokHLjPi50ey7IdPFYKxIK
y09iKBEFoouKwZDanq+9FFvOA7n08nPwwXNUu2m7O/Kv+DAU+Xe6SK/AWIHt+m/+
hbSohOLXh2y8dNAy+HoQc4y13f+YNbm1lxPZf3qa9u2T00RzDNzyFbroSe2zUuC4
jmc+vlnBtq0U6+5aNwgY6Cx6TiO3HItUAf6C7lq8JLEfxJ+L/DEw1D2lEg5Tx086
/aErPMB1BRXHbCs6FNu6sSNGYUwPe+O6yar9z+x2z24Na7QHGp4JthAkJiOHcGKL
5Fx31WFvdu0FS69hehUUjyemfJzmA9h/Nfg4V69czA0FxTnMuKz91v/5i+YEcAVB
M93vsK80oHENeuAYzRaiwR+EPUs+3fYDIRe0DxilU+LckMJF3weLgo6kgXZeUD2l
WgfRHyQFQsIdvHa1JM3M0BiciuvAeUSkCZlMUmt4Zw6+AIylxzZGTv5jp94mhXH6
6JZXydeyDMX2FhychfAgpio+MdmorIjPeS3xA4fSdWpkpff5w3/C4BREEQ4d8XkO
5hSMpYlhlCPYoQ5KPP0jN89uYGPp0FXudnLa2HZc8CO5fdcOVRZQ2RDzlLFHc2Sk
28OY16uagougBLwyKVAIKzrMHk5P0FQYzdCBby35kb56+8fGuMAfUCa4uZp/R3Qr
xO4Yv/NKHEWDksOmCnBYx+aFP5WxyIrX2HhVEDQ1MRYWrl+wyBaRgn5GMkxboxhJ
nqeqWzqNX5p9EgGgI71GBqeaKsSF5BT3Sp7sFNcfDCQZYb32b9Wu0qbDlgcmx+OR
YXkwCenSasazAopXNvDNBIdePPpaiamc+YaBK3x6Csl4a3wHTJkvDFwQoTeMl92z
W1ONzcW0pOSEgIWkU0cNTBtyOznoMQ48AEiEQ+VPbkziMd4z+9Z71IUKwveYqyQa
RoLwLE1AVXUrsK9ShQH5TzheQlE+0ABFczNIYojwC+ttokXhVJH/Gyg9VKnhucFB
Ubw4kWsnRDqAjCZ+Ko/ZGePi95YeIqu9KAsps0ggvegvXeqWQ5vRxuPze1MwcVU0
+PC38SpxQOPPt1w5zomykoESr/4zejubWgeWwL2aPYkP/Nsy6ptjhTMMgiVto6aG
Fcoip/6nWCYDzrQmpVT9M1HWVaZDKOvPTitJ9qnnTuBIrqDxmNpXri+T6cHlWilA
Y1IrpmZX7UcbQfWvOBUKlBAVXgUPyzJIu4YkJWbQCYFGKtJ03wEw60mGKkuE22Tm
WVXgRTOipoCy7A/1ExM0kuFPq0dIqXufPosM08xsKkDFYw4Bld1YCWsNESypcwdZ
UN7RNuPya7TlSIOOTY66gqupa8cLLkw+ZUyZIer9S14B3t5mE5/GpWO/HmnC688w
vVp4MtOrQZnB2N8PMgAKx/Y6T1jLti8kpuBS7q0N4u7N7y9KiH7vKm5+3Tt0y1B8
kv4HJehUoii6PwkUL6a2I7jX9snYr+blLdXN0lz9UQUmDnp5EGlnXbPQ/yIMSUfQ
Xr99s4qoPZWwFMitmYfw79+WeUBLNd3wl+qwXDNohRcfShjvPPwE2kY1n2HKIFEB
EyKQ8AHjjQzkYN7pcVpC0a5q3pVFrD/gac62SevXqSeS0awezogKUh+4A7QG2RWI
2tQjSlfU3It8aV4ARFAlNKriotYAJKMFxTa9/uL57pZBxAL3AXMcGj4CfKDjIl31
Tag7GWoFoqFbs5qsjP4T0m2Y0ssIl9XltTpnDghx8lsb4QZsMzMIPjfBIV0t+bHK
ffIH6eESMK/O9PJrtgicQJjF8/l35qRfKclGbkTdwjyTOAB7JXHxMamUwyn7Q4Zg
goEoU8HCyh+CS7mJkSt6/cPEydOuCaePvbbttQqPs+BgI5Avc6xDo8Rp46tPuhW8
GxdwMegtEUH+om7qzcVCYDnAmOCpibi0JI+RAiOi5TRCvBQP5llmsHGFd2PoalG/
fTep5R6v5/bltz+zpykUaXwXWnzD87gMkdNAU20Um+iKbs82iC4IpMIKBhzyyLCH
HWvGsTkLyd9PsJvjy7odYXJOfhjqk9NPTTGj9sdLFXXxTN+nqSmMhRueKU/s2k/k
now9/qmRriZCiqgSMKlI6ErNt6DFJNYCdAKUR6N+CTLzBxS8G9mb8XjBpY5f6FkF
4Xsm25ONMtGHC9BXZeOaY/x92cHUBUS+BF/eoykmwSuSSVC/RTlUXip7gXXju2DX
z0wds2DkdCy0E/qrBT4somfLcsI0s5WEW6yNZLmiqqjsQBVIgwtOVdvdvzGBQRyb
MSKpyzDx5/uK2TbFdbINvrfV/bxh7kD1kr2oBitXT/O+3lONPazYXSbuw6yFZjTM
mCtNlh9JRGPwVIJVbOvXtnhaDOHhmv+tGah89/DHf6roN76h+ga9J7XNwc6Pj9pC
tk+cpDNah2wQCz0cxGIZPAbPEouAB0Vxy5cXEO/goFV2NWtDB60e2T1IdUwm/pt6
91YTtC3WI/s4pMdfqT+UKEHLfY+EtojujW/jr08sa1paxijwbfTHd8c8ek+iGdow
Hi5nyQ0Ft0TfoPHrIxifK2AjP2X6BndN8Bg/6qZn/0GFOVi77QvJoStXAVnDlYDw
zL8XJ4f0/TjCCC61VBGy2cHOO2MiZzsjgKypFgqOPxSWRV1kPmGZORRuz9ZaIo8q
7X0ARyxKJyhV/ATGcRzdX8iIcjviA0yj7ML+qXSs+dpS+jVKhJDvvCJX1H8CQmbQ
WyG8kquD+kDfBpRsHUzw7ZnTAS9dCEbxkOyUiMnSeWNk/IKy81Ng4Jsk0NX0FfR+
gxECyF9muIBHkJay7IYiwcrpSNeOx34dVH0ECLPy2KauFahB3AjfR2wFXFulW5ZO
oyU8OM0+QrgGGeH7oyojZQUPnWWRDPDAspb5QqsFmEs91IwicB0/iwG3+ZMsaWUl
JIaYisDMhhaeq0RbW1V9n7jawZNhWg8nN5zsm60rm6QOhsT7sHfdiS7qsW4sS00u
a/O3e87SVptZq0EejtwGrHgumg7vblQ6JdirOT6qY2lmy9F8cG67xaElExnA0EzO
1X5xKGKX7BMY5MlcI52aSWcD9Akn1u7XI4x8L7W7GtMhvaEM7mZmVrmgnUnirNGh
1JMgzMe4gUISBfHZbGtQaDhqEPjy10BRwH/RqEcAOWx9hSJRJQ4ahXl+rn8KTOSv
Frqg/P3aeQ48GC4gMfkWxNdNi2/BdgCtQiOQsCy1Bbr+W+dTivSV3M29SAk/q/I+
Gzbl4R6emmdjpMuyeNuBGit1n8e3eRflxYBmq4mDzbF2PhdrK/npTSEsMc93PlWn
DXFILEG1ukawd+UT8U0WNwB3ODIds9HqSEn+wefl8yfQLec4C9wiA6RS2T2cQtRS
xQaJXaRgZZlxc00amb5GaRU22KI2hXb/U07+HEU5xHwB3jT8u5c688UN+SN020j/
gmcQPAHSHj6tyIldjg4wrhMPIUEiT4MQ+NBobLcrospzObXt0dG3ruBv5f0ZFomc
VA1z77HcMmGsd6KoZUwbLU0WhVHb/Tk+eNfXbfLZwa1cjC8IaIyE6ydOmBuv7yo2
v5zT3Ox+bMl3mNdkY1GNrTORlr+pbLMw3G/FtYbXDotmszi2E/yAeRFOBLS22PMq
1TCj2nUdUm/F183NiAFjpFcngVsbXewmJ97dshnjzzv74HuhMhoLXKKBOHiV0YS0
x6qS76ZmKwW6a3BBD/H+umRg4D3k+FZ1KHm0UXK9Co0HYnNMxIfbQ6QoWFHe6uVA
D9kYQ7WhA1kcOwiSG4Wtsyaiwx6IdwDvNKyrqXHK6DGY9ff3zUdEZVPYo7koRhr7
iSxvX+iNlsrCvJMO/XZu4gziOh6CytTIhmJLmYSLKae0vKoFtZsDfLgsi/xm5czV
VONXOMDTIgHavAxHuHY7gtdRn7tyNNdPNBeGGtJFtKJImQuhl8UMHWD8FUBzjkGJ
q1h15FmWlstBP4uOMLmk7jYPR3GfjtYKofZPOSJERcw1ng9WtFZq2UnL7IaCA/e2
eLaCJYY0nHrxiow07aLxPyyv76+XXRifYJrfJV7+ixcgndZert4YxJp9Chce++qc
6bbGOswLD+T/qLkkN0+wZowd5HUKfuNv8w2DuNHqaAGVfHXeQU5dHeQr8HCrcXCu
bbsnebbbXSSXNzokSPpFkTjzn7jed9Sk4satdFmdC8DTp5j3eipP4KjBXFNagw6z
Ibnc5nrXzpAYbzVCrmoUlRZdjxt5q98dmxzne0NwxsSZmtnSgwlnaO8IPy8LOHgT
q4mfz900DShDsP2EwNDsjZdQ0pgAma1ugIrAZ0BThwAvoik3ksTtPLNG4BFoUgZe
XLYnrVbvBGyPtIFT5PLASBRZDDlFBJJ4M54UPSDnx8D0UualtU7PvsCbbtrWJoTP
B23rJkZAQlXW31mmz/ABnwoW90zzLwSsGSqfbe4iXaUqJgiPH0FmPvhHCK1ScO7X
3BLxHh8sJF7r51czfCa7Zusrng8OXRhxcOY1a+Eom8ehiWX2NXMt3fPXoKoZBo6h
z5moZi5WRsHuDnUApGxLJ6Lfz3kCD/fi2fHdfEa5+aR0c7LiitYaChMqXbVMkqr4
Ll6LcFlvCsEYFUJwnN3+FPPOsxk/VKlallJz3/FejW3z6x5ETjKaV1SrmcFgjJhx
1/KNaI/lQEJOGm5dgDRhOTbGRbHZOoLR6nkXNq+5hiKQKSk04jT5dik09FGK/l9S
6UR6ElpPCMRl/nxypvcAIB+KKtfqx0J+CJmFLyZBdn6KwCRxmA3LIEON9FtJz9YS
nlSTqSU6A2kGe30erLFDnNGA6jRTX03XRvhJd/UUgxypq317OC+q8O+MMXE/Z3L4
blAIrDgx3F9SarIvaiPGw3RTlSJRwiE4n54qg0XSALRxtVXRhUaMB8xqQ4kA2+Yi
Xmfq9oYdDF1qM7lwejhvNqX5JP55WntHS3xc4Az0WwHesvuKmnDVl0ZFYpMx03Ki
jB31Js/soGut6TXq/yqyqzczthaJK5I1P8tgo0YsywcgJd6IqlNHhFCul/ycn5Y9
DssAIl9792iUhv392vd6+pzA+VXXn/HSGe6ETE3muleXe9SfDAWs5eh20s+KmBP3
tWYh4VUIkV0ebcC2gxaIcuvoDi9PcGhglRqccMxchyBCv7qaZusz3l1b2J8/xDbR
ojgNX1kd9VnHlnMj5+9YvTTvbKs0p+QXLNpGVfesB8id48NsOAktDpava+EBZtQQ
9sQwGhnM3e5RFgGTciqrIfmbfqVO238qPealnCWPc58rIA1uBhBzKkJvXq3/j67l
Wu7poVhu7Uj5+fi6cXqfxmPy2thfxAfCWwiW42oiRzwflzu2kIs7e9+nJAtmgG/X
xXVZO3ImntsTqT9MfxSu2F9/Odyr4DeokB3D4ZG8oCwsSO/Kt9pXZJX6geNmbkrq
JF+yyNjcFvtuB30vYBc5X2poWnvirhf3ubtlQSx4GQIFQAB4YzcOlqzA3aQPJ4g1
7OUs0vjtJ3kk/kROlq7imY1dg2cSXPhvy4ozUh5K0E+JGzMmOg/gLMAxDyWo5O9B
/GvDMVbknMZWIUXgdDDsfkziEgRVX+q95lXsenQd/88j/gM4GntRN92s+wLMdpG7
k0x/tRPC3ZPFo/xGZU7C/3bRR+aj+G1Vx7MVGkFFIQwvgHkpQ2v+QCjUf+pW//pu
jQus9qT6DmMVCkJ2w7UierxNAirfOjpuauCaraSXiSjRSHgr6fVXxRvSriTuZke/
JQd2PHbDX/f0blNG5FBP+JNAtpUVlo+8LXF9a4W432wZZGywr5kGfczxSJiIOiTO
DbHDyX9bKSXvQZ7KfBXCHjrsluAYAarWVHCjZVoJ8FdWM91RbhQAEN8fLQl0m5QX
qO8NuLWONJdJoTXCzNAZSZzuHEN4E4LjP6cdIso8korhVCOIq04CRmV0bjNx3RPl
dJ7VbLc/w/s8s4HI9Cj+Cz7fF+W0Lxd3G90e9uvYsil/O0msfK03kc4gpYoTe6No
88gu9kMr7Aiv51p9lAkyS2lnHGx4s1SwKKTDgnr+h90Pd3x2T+8HJYomdTNpnm9f
Ogd6+5HJt75BTsq+aUgFduu0UWXZ3L+SWoQ+Yjb1Tb6wBZIWKjldCOREoyJCB6C5
BSUsrVJOMry+nI1/o6IW0eBBirAtVJ7VniHNeCsGUBEsayJyGJd9f2zOJMqLtkd5
gRXBUIsFi3dhBXsde48R1Y1lB5J4/PPD7hmKjZPtziew1E68P14wYpRymTe53Tqu
Bk+FRFWEKE5yLGUn3nRIPXxV3b9HPtNTrAF6DsIgi5RuYYNap4QxTDBACu5+FI+2
0WsfHg21svzRpZGyADBWJFL1vT5osY/0MXf+GuG/MV0X0Ozk+t7vLkkdfbJUGKwD
E3sG68/0fhLDW56L6h83WTSPbsy2WEcpuFqvkj7hc/NbT+EbQkwSnylKY/+cEFcY
QdZbES20f/vpGiRrRZ3r/dyjM6bLXt/KE6OdbqvKCq1mQQt2ynkXr/yctDA+Hq4U
ntKI81XR69QFeJNTo2AN7I+OcOA7h3EQTx4xtDQVewI3JM/cptLV6Q1bfeX4lvlC
kZcZ7JCjjZ9EIkVoLnffc+8aIDd3Es0j89BkXtHl1B2UZr3uFELs+5K6prnHTFAY
aMOfHLN2ZelRIxzGuWnf2mOAnKb2BGeimikLWcEvpKLvPRgO6a9rI1d7GIDatoPN
TMJMzCyXNlTdmcYr+wwAhxN8VbbkEDawuchO2GJj9gg+JdlqtIx6/KO3hBsT6RQ+
S84PqgoobjRYhrztumn+JtD1kylAcuReSBki9cLrAsu4ntLUMqFl8cfHIe9SctwZ
N3oTO8VyyRlaG0bekg06r6N0srzHM+bI9WQo44iWz1lFhrAfyPv+Jg3h91h8R8SN
EETmSgo2yWNWOP+3W6UqBN9IA9XcVXkJf6B2fx4/Nd8RGxwf3l4nVxpxREoD4gj5
1G3ZGQYOwTV9ILzGSndxLcAeaNUmpgg+51hxi9gealm8NJXHaoKjB945nw77YaST
kUUI+ZCMvaI56o9xHOaQTN6FlWnS01cLNn4twCJ0UpW3T2HSim5D5yTeOPeakNqL
SKaHuzhAKb5DYBroJlIZ6LXEsKuU7W347VyhCYsyLNRqg68Q8OhzXZR4g/9ncl5A
QT50vrC3HYwON6JqrEQMhjsy9ImWyMSBWuJ2udUoTz6/T3SHc/a/SDJuBWU2fVkD
/FatC2dPWNfBmSd05R00Q4OEkiIaK4olZFnTxIR6OnhECDNEro1E/hgMNqhI6Bn0
2O/B6y4YG2i8M8BbBUsjyTzBIJFCWcoiSec+SdmTPad9EN9L2uStCHfen3ytF3rm
eKU7UXoCW/AS2lLBFnnXOql4RG5gRWlyNNYmkwN+zytwcC/bUEnm4lUBHWXaAk4a
vanzMkGfTs65jBy9sJgR/6hzodNkDZl1fWVHDRhOd6P/ghLjODOAg9y6ok5tXX0H
TFEC0C61MozyL4v1GvwUDunfbLri+3fZIQkYXxQRciHHqwhxt2M8LOXEiB2t2XCa
Cf/9RjgReNM0/bzoWz0xBgqRHHYPcTH/s04ynX5+Tv495jDH6lWQtLj6K8QTU0yg
HxM9xMQ/SQacDh3m41cLGTfGfQAe2g5MLTCx1xtaA2H1BGzQdNOFFGaEG4SQaeGO
zepAnmX6XebTCUdrVhd3539qZVQ41rT73cl/hbw0D8XcY5gbK1gqvuCZl74zrwQC
PpHEYyMDN9sUo+zkKiwnF8K1KSw/JypSCQOiSnj+6KMIiw2D3cAic3ZsdfzWsCDZ
BkpzJ56jd+ozFBJnob9CSOwSnhF3O0bWW96YbTDUtuAyGqhXzt2fGh/pzayGvS0x
LlIVYhmP0wJJuT173wCH3PB0LErVqpdm0H2uBGrI6cHr9qkDpX0bXo+DHhXgqCoJ
+ikccsNtzcB4qAyDV/Vr8wnmKvLC3p6xuSelemOl+HpK/S4m7owbKfyElbncUy0B
Vgf0anOuEDmXjLS3eeV5W7EQnkeuAUCSNVyK4o2f4a9yy4GXKQOPUaSUWhrZpaQy
heG3orvsn9D2LsQGglP9xsOZH58OURhKu2pCSOLr+sfFmG2ft1+YE9LE9wRQKtqJ
LH6tVLZOdL/4sFY4ePCbkn1L1VWhNG1h3skzcHSLG4OrGtWJpmklVaA64ViDZwTD
G7MBxbc5sTt0XEtFle1vdF6BViyCuNt+IKPAl39A5EQ/3TVymVYeAMDZdAResGNF
Z8YaqyLCmH0EI1O2weu7LBtdH7su+3ukWOL7GWOZ3K1/2eOoF4uT9ghNQIuJlLdT
oCDeBdQW6UNvhW8+/TCYG4RrAZDV/2YK2LHXD0HcnTqGM/aMyC/ksE9dO/JppB3o
neZA8m8uJPpi9ICRAAJEyLYCYoeoyP851ytsOgWFVxyPxGtevoxQTnYYT3eItkis
NK0/LO0JeUFEEVMcn1chogwKMt3sxN4qXjls0kkZlhx7nlfWgDmg9reZVlD014y+
FFxAIHPD+f5anrJHZYG+wO/SDHSCgd+VS3HDdWrZPkad0kJUP64UzBGSyk3B5kiX
onhusmMYZUn5lk+c0mAumRB2hpCosgB44QueFcmlAoUcnDhSqjJHatDioxzxdJ0t
Lciw3CXf1CJIN9RBdhjyfyrDQhjiTf+IdIeypoy/dYVHAdVe/qYJu2aqoxXhPwBS
4SbvrD58z/UyEr2Kl7J0wjOhZKjxX/AHvvm2/XeKck8N6Ca+38d89ZD7cdk8bv9R
A0V1GjURKhL+G1s+4OAQrR5e1AO0WHflZDKOGq02MWT/LTvXwrBrsUMp7QkrjUUp
ssUCXs2PKBG0vwaz5gS4CFNN7yiHAUjspy9YdmFd0uoJh9/a9p7ygrNj8zEAaOZJ
stOF3X2oTLod2RnVJpZTk9Tk4Pc0iDJ1WuIyKpvn5GOwYFO9bjgGfrxfoT9ULMr6
dykZ2yxyxXL1KBrXV9gh3hY9Zemtj4zpvcngoiPFUox0yOIhGyfQo23sZC5YBVAd
N62TP5bQfcpBjdWqjO3+FR7IjwSchF+bXwpg0yLB2Sba6iHgOHubU33ed/HG5lnL
0yH2suqattdj90gU9OXYVVYEfwUVs3L2sWXYK0P6ew29MVl2Yjp7DIcFemKGstRf
3PO4p34S7eLXvQpu2puzRU7MAGQ1LtNGHIb8zvqZ2UiubPlko48SYlpk6SxgcefJ
7FjojmQPkoRo1Pf8DKkDUMSCuGtVjcpjnJF7qnTwMEifpwme6oWK2jVfVHsH7pz/
UqOYKaYF9MBdt/LPOH3J9S0HLKV92cU6kR/A61RuEUfiGNCIBjB1vlakAZZzvx/t
6moeAn5FSaCoOyzFT592/RguMgJ39oq/qPVEW9S+OjupBZwc7G3x9d+j8jW2lc6n
ze5FoMoY+9EpqX07p2sPBKcwEoh1GMeAonnfaQDnqT4jx5fsga1VAvA09ZFfUC/c
JgV/6Ay9+WT/c6G3Lx0tQVYA+lZVx2fOq/0GALV/H5KQlr0+uCk/Mq32BatoMo1p
9XVkcGBC08GmPlri0O/BP7xs8q9zFD0kMnz86ovrPveA8G8BDYyvKa1exQQ6DpN9
KCPW1KJylZe/Cd05Y93IYCx7jpnE+jn1EmkopfgNBPSA11gNYFXRJQ6KcQuI8sq/
AWtPfu7FzzGuJRhOMGNfFPSX9CPZE7y7oHT5DQSMLhraeI6siN8zO6jldEVmgEdn
8aBqpjq23ymVTvWsCvwiqCn2tayJ0whlcc+PatvyyQ+iD0vo8dC017T4rVo97wP1
zjwXFyF/Gl/xbdFjVaV0W/UQGUxpZApO6FTVKnuS4mqJrmCLWmEicOmx2FOv3JAp
c1flwa12PGWdmgYXLPHHKLTpB37jxCWev+NT81lM2iF+5hDmokUSl7WFT6JReg7J
62IdxfUAxt39aTY/+Mv8qB9mF2ZZT4Tjzp0cTID6jV4EC0uQTvyYjBEjkV91MNbo
xhv03NzRfpEffb+x66akAg58ujialEKfU9fmUBqYcRemq8Claz3j0YlINROBg3aJ
l0PJ2BcH1EYt/1zi49g+yuoj2MQuufNuAv/DkYmEFfOnGi9Dh7Fc1ctBY91jstUv
Lrht/V3PfvjEYW6BSy1XLq+0Zf7OAWdjwXPwmIN4TS5R8RsZimrAx38sCCaBKPUG
vknXnvgnKjJsR5DAHZlawVWM0sZzs9VeIXT5gLrlPf3Rh619g0cq+T87eUPp92qh
Xtl9ZNopEewMzgtT2wLOg6opQm0y8md0zhubqqP4btmHIXTdjXYGNbcp3fGHH/45
+nXKOEl0o8mZ+Dhrlpd0Gamrj3YUouWoG9S4esxdd2oSxss7sk2EiX1GZ9BBHGw2
DVM0kUwh971DKbILmH6iC8+817kRgWngqGbIh3svo7iK/Xdyt6OGG3Z8q8hjTy+a
V8aiOSzOmnyMn7vXQpI9ixD7IXKo8lMj5lvITMM1KISFREl5xMhEH28bkHXK17WA
7fVdUj0OiWVFAHDGdbze4hT3y5i/aoFddOEFtd4Yu7fuz8jKlr3JvLJR2/LfCQAV
kMjIW6EG/8KkEqL1C4nsprooYxZajTrhYFx8iZ3ncqDTLyLayoM0CY52DLdsvJR2
/436gy/u2gYLlxz8inItTVRewMg2lxd/65JNImGQdiY8QiqYE1WPhJNXWmRcL91j
f3YANvP+KmBwfv76cyuMZ2iRqkynHrNWr4pkmOXWXfG4xZUiQHACBknRsy8gjT30
eFGAFZD+NYkAeWaCWpG3nd940vvo5QADbCIs6+xGu35OQrwGJ8st3xBdddwhy/qV
/d3/GtQVaKbtV6g/iFxibvnWV6l8o1UUpZMvKFCHakHIWehrXn/mhMkAXVANPHcu
U6H9M2HA11fAx559+1nrERT+FhD5LdsJNmqHfDEUcq2htrGYVZkCUc+rek3nNCDo
NU6t6D+4d1+pY6UKL82+C8Q4qjM1Pr98a2wlnMUoZA2Eji2qo0rUsgO0cbDkAWXL
i/FT9lgAYGnmLX/EmGKTQ3t58lLLA/pl40RRzSsMFN8fJ0VuMJYlxViQ73B4tTom
8XrPmvbGmhKd7vTpQRSNRckYuIajvCqMMR5xFf50ItiLyDurRR+cZf1NeYnH26FV
+2zxq3ktIi8zir5c9LKHHq7t9rAGyi5y3q45/RvB47AA6w6OUKJpl3OFTY0hYiBE
ZnOMXS6pHVfDPRWkUoqep/khsly6CnPM0Gc2dpI1OFkTLX4KePVpp6TsYD/GEHhO
VC57ptx3f7zxdTURjAVT3/k5CSaxYsubKuUp5RPyVpQtLz9q1FXNrFXQia6b5HgQ
Fnrocg6W1zXGg9Q1t4ZTF/rxlXksUJR0ptoXfKlmcdub6iQVbY9jF/FJwC3oSN4a
niKMunYUnrXVUXMsg/7q7gT2XNgWFFaArDOSuxseT8VNcG/kUnhZT7q19GCAxwRx
0Na8YgimLKkyOPhhMDt4o/JG/lv6pD8tqgUHRyluxMDThbnE0usgL1LRuUE7Hjmo
+wtJgVSdInX8CwBXrtq70SPsRujqQbbaU0c0UM2gEHMJAXlKIarcmNL2siJAxHyz
EGd4AhoSEOAGTyMtSc/zlN5qmBJuhqWp4Ywk3zXlYFVu7lkkKTkn04xGgrEKhcPr
FOY3QDIM2IIqby1gbqY1Shj5T1K23v2jsvicq6XpTg0FbkJFzPGgzWoYNpUrWYp5
wAdv1qswOa/YFnbLlimH5sFXHhki6U5MmEwq7jEnJkpTX2pxpqc9+q7pmqTgCjYf
QV1oHy4Vw+IL7oPvQmRRQfD2VWk0ThLE2ZjMd18kFOyA/w/Aj0uX1jFGRpA+H99j
FBBvyM55sG9lMus40+ZRZFXhkCZPWjDMspUOfjs9HbGhW4TjeHpK1heO0+UxvJHD
TZvJOhCSgLsr9YLamO0xys9cYVz+fWcqPUQdwmjp+cft13jSbaOTAtyE/zoiJSzP
kfilenTuliOTlF/+9/dBkvyIhqdAEru30ofZ3zkPK4sJWBgGyUxBpSC7jBosVGeM
k4UKpWK+xCM0rHKCphfJQTrUXkxoLTwd9I1pOEFkPQT/q6GtVccqoIzQfc+UAGIO
dYgoKeazAopScIrD3bgCTcQLTORbaaYzCkSTjH9u46uheg9m2NuBuScLDhegOjzO
+G2laZJB4J6N46EsA66X6SuIZVKcpS3Zm9NEcqNX0+eTFvkaZIWUG8J5e9HToH0x
RVoiolFE5WoQE2v2W6Hvw3IzgKjK1ElR4drZhsaSwNyT7rr6ZG740epiZSv6Wiag
GpLOFI6CG/c8iicG7eTwX18A2ZrxpJdZObo+TJiJvVrYIP/2jfhluWzQWDaYUWwN
G1gPio1o3hadkudrpNAk3sLtmqHnkLQBLnaddLOAk3X7yAgWRvINsJviTF0WybRY
dNW5PKFKHa5TKyBGWlGVcx+EDwroRZ2aIhxuSgFqwALJHgUNtkZTnR0yLTymLavw
Q7kqBYptZ4qYBg1wwdofTiREjHEdG2WFyd7eawsKKmyE+6LPISOtZtW45sLcdJvo
Ma0A1NV+F8CcXakyTKI9M9OqbPIR68F5Kxn0EaZTyRnCUaLLAZbUAjCqRhi9oqEL
EESdBNwvXAU1wq+YjXcWIFsTor34VEFd2MQ64PR7TxmEKvFVwAdLJkftfFLNciRO
gHL+vUXj7zXTNhprAg8XY0+2kGDItOK6KUVojbch0JNK46/Hv5N0VJO7V+8KuSib
heBAHPoaa5Q8dCMDNrezWfgs6QlpiKYIE9LCiZhNa9GoK/Df+K5qpFL2ZTXd5CWF
jqr4zPgRVj34ZY8pmXxAxaOpFXjhsFFJk9wgJfud2QDFW1qFkQDcr2BuJwpwIjcx
hsSbzBNcf81/qRqkCxa9DnAPPJorsYFv4IwNPcKhikhub+u9WTXXAd97qUE4mSsf
TAo/N0JL+RsSw0nrcJXOypnACTRb9Jy6XJPAbd3q3ycUtzrdJrpqVg7ElyBmaaO7
6xHKZL2Kr9HpyxMzsm64nzrkTCrfKhBwWNhiejqA2VIPE73KcUkmgILQay3hbYRL
TBYz6MlmivqlCFEfbms0/3zOj0CGh/buPpamGnID6xhTOhMKXazN0WXmnQTtVufD
uk52a4Nl9sltoIrT5BMeUTYvQNHbsx0RFiF+p6l6tJ+anFWLSEjGGogHZCmdaVbz
K/hYNn5JZJoOlUQlzm1+ZpRyrWEFSzC++4XT5a+rioAUaiKkUPIBxxRHToxSa/Ax
zZWfHyxOr1vvQZ37rOVmWzu267uO6QSwTrH2CPoJC/EKiFLn/Gd5jk46o4s9+qUF
dl6L1MXkruxTb3cRNKaPJYmKobe5trhXJb490UxXrduVUmEGkgeW+0U8iEUMtBDv
QsNk6/LdpXk11kCwtfTa9bfP24pm1eLQr4WhbFEVqrtxc++9mm6PKwfZRGq1LJx5
Nw4RtD7Z/xPK9EPBF1pT15W0Niibig2AXouE7M56IkIUu3jRJRCUAhs6xXbMQDoy
eALL77wa2SMWSjjzM+cSPryNjmrQS3jZUltRrZdUCwE/dtU4kL6lFwqGBnRLsORp
Eu263tnSillKwWvA62pvJrRMgHDF3UA/16SIoMPav/ZjDGwRGXXpv5DVUaxIcjS6
jZp3+J8nnPriWcXIFBh44jGvE3Je9DQVyHKPchv2jf3qfgxV/EYgPXurCf9E4DAi
g6O6h9hVzcK7zwBgn9tKUEEXjUeOzdhR5aAUZwd5hFrnAq/D3XuuB0mcauFVOUlv
0iDxG+ujlDrsO31jmXAxScF3XnZkomrKXU3VQuwfR+Ke94prNMHF1f/07LUMYGdL
vQw36h1FSJpqptiM63XUNV5dp/28Wno+tH3u7q4h1/cciNBPcl3tSO07ncXUy1Wo
hR4047GxcQQp2aPjrOVm6dSLdGymzPXEpy5d1ayszw830jpn7ogdBcGkaip8rQCo
bbsjzJqNhugWcxmMVhChyaQ/NwqOlGt9gkZRGOsheQDEAawu9bH6Jsl/RN1OHQNP
tXeopXxg12Sc99aKrSan9ztg8aWQqQsRbHOYJZAJLr1UAw7F8C4JrJL/Yv/dtOfg
hFbshhcRSg3P/ftTV/gTwTkHZzpcnFJQ2Tjog5mqLOuKGQiHDWbLIKKzpc/OJSEU
pUawfomlTlrTE9tknsLkMnc6cbuS6UHKoQ5y97TTcLjeDifvGzqvKktXI9pvynFR
0TVM5HAXzqcvLGg0bcEIFL2NG4bdCSvRCt9kfaa0p2P7Vb/101WjYtAjO+0a19AC
sMhctzkt7hsxiTvH2TzFDzlN0QesyeAmnPqbxugYhGgWOpoaRaaupOAFKbh/eYcA
dsaSLRWXO68yMcU2QOnjenNJg8ckCn/+eET+KUN1P4Yz9l81RCkwn6TvcSR6EQCy
gI3zoICB1gfH3fGfMnG9AaDBPE13mm6obR3xKffMfQWlaUq3UT9PrD4jcyYF+JLy
i9C7JmEGOW72a9l94OzmM0Juy1/pIVkeG7xXZlu8kRkRj+onHlJe071bLt04DCI2
akOcChw0l19Pu563Wng8nQXjYiXMljY4l4/BkGBxtIAiIHAib4LMZBXvwi3lAUnR
7sSiT1si3kC/+nwqJxYs47f+8z+zhNmZj7HUQcdpSKds+D/ccI7ylVCrrLFBCTmm
g32V0QEhuXbp1XWxDUMfr4s7F/xuIGpENZA4q+H2/1swECgq+bdZkFnRTT3lD/S+
z418ZUSouOp0ihXkwZDLvBi7Al6RxlROnrJFTjTV+Tx5nsV+O98SUQ08KYgjYcy6
vCg9lU8GQnRwP3dxncTNO/fuleoHd74ktGznHj9VV9yZ/Bs3QBaUcpBN/xSUjrEx
uSFLdryveyckfLjnudaL355s1lv13tWYETMk8DtfgKU/TpOY6eJqdNuKOmPL+1lB
dm1q4+gT7q9eFgILyEiKAG4VDZEj+0snZSPS4c9Acyjd68NNgxtwP5Gh+Bt5Adhx
02T72veoy0S+aFFtslq8JpAoHWbzmJq/0AVyQaA4+kaiwkgC5CyiCzl81ajC/N90
0oGI2sTDP/xhfj/jvpDT+As0gRnCWF9IGwyvcIibu+Ih8C/mm7pr+7tkjiuMfrEG
E5oCRy9wxHSFbdLzjk6ViIJp2tvJeUkyWhnlWW6RPDbJA25ksJX6dD0oosIiUPOC
AldtrXXYDqhu3OuuXbikM3Y1UuJ4d3ohsx8h6JZXvKUvBNVLvGSa03OKZGl5X3o7
4mmR6B0wQ4DYt6bL4KIQTjAXyRpibW3GsuCAAJCYWXXOJc5XUuLr0KINTemqFckR
wEw/3D4Kst0lQRtj8DJlgV/I+IEdSzK8o6H00sutEV6ezddhIkA6t3Q7INy7U6eO
qcO8gazJR4FtfKIOs7Of/ros/usnL67urufwzq3B4T4Ea8FkS3teij/uO4zsJC8s
riErTs+vEahG7YqIvpc81oxyJgV/QnbPqVIwSjubh/E0msl4eZpjk7GBSM/zNJfN
v2QoiUw24x7J16W36BuCoZlZje5alQonQqCdI7xuQdeNqA9C7UMz8Qe28dQOfxb8
ModJcvouSbGMUaisrfiatirCg640bnUzqPLoatAA0xMMY7w7I8xzS0D4t+Bm2x1F
YnuQlhE18B4s9N2UlHyDQWU4ut8GiGMgmMaUNNQ+Ges/COUrv3y/qjPHHtRSgOyk
ugbEZqmFSNkgwe+ffJHVUU1S1NZcBtzMTifnvvdpVbuxw8U3Thds/sUDpcEAQM1m
dgoNSwE4Jtl1rZkkcSaftomTsobytl5zlD5qfnLW8+fKakptME/G/xWwia4d4FYy
K5peDWjjepZ9rCvc+1CVXZU6ltHRU2yQAXUA7m/aurrBvU2hayMLqyoY045ioGXz
Q27+LAxk6fKqpaBSBsA+AlOQRDdm8qx3Mc2nGI/ou0Ymsb1sgo7bhMsKaJLvbDSM
MNfyT23VT/eu30WjUakDT1z0WXZotjlCKeKIeClcj3fb1Paqd2janbhRew9kEucN
20e+elqzZGRQ0gYhMgBvE8WCfSnWdaU/VHTecCE1qWK06DzGPmnKTjofwOdiur9j
c/+/yBM493GKrZT54Jze/w+H4zzyWPcOrKVKYgj5SEyaF6sT4BX8TVpZFnYJlN4y
Ac7glL++HOEmgEOdRPJnDTasc9MPaYM6uApZXwI/1I9IQz78aFrqrkyDbsmuh7m4
yhxVer4WGKwG7ZRYsqVWjydXcvafYY3OxTnhKDGBT/TBoH1v7UCgs8f6Xjf9mqda
uk8okO+emdd7SWsRRs7wHFgFd9JfMqvTA3Y4ZU/ncXr+HByhuRi3gXPzEDPF8kRg
R1JRznuCTJ/4gLjeQ+vm7lTzZYvrxqWDwWYweXAMtCs2o7nm1Fax1wkNI77kBfSC
P/UwYVsEQH9061Drl/6WQHMnUP0tjDCVZz/g2wSMY7Mr8QdXVddGitNAxtYH+R3A
UzSKHZWw7y2fLYWwg9xXuK+kJBhfECRalP4cP6OYMzOxweCygnRkQQvu/8jHtlkA
Pn2GsfwWk8DvZJlTss6uo2VO+2ihV6OMsY/OsA2Zp09P86rQafWhWBcXDImClG54
eGIamHDUQtiraWgTNICvaTMfkquZm/kAgfg/HTJ+EHcRyy1zUrl4G5pL76rJw9TW
mSAoqbnRwiFrbsiS+yIjeYNj2y3jIpFGEff5cGzhwWtFOo7Gyx1UJFmc/M34kynb
MC8oNDKFjSKqMbBwK436HNfnpVij3vBvN/0Az5f/5U+t057S68YIjWi3mARN7YEe
96ghpxHR4e61SpG7dH2WC82aUi2aX5slsC86eB2sb2xTvVORdAfibMnR2fnPN5WT
OCoKVD53lSPFk5ZgbpOCefK9Bpem4emtMO/CNWdixiaWsI3jXZ4jAWiXJfwGJimG
8YOHkId9zayJmPU8mT4hQe662wXPdftW33Trqf4UqZ8E5OXseGtt8NGn1yNsK6r+
snA1nAp9eUYTkxeIhrl7j7rFYVvoIjpYXTjUsc5RU81zVgN+dCI3jX710Lbtg9kV
YIZsnVR4VFKHUuXpLM73p/YGsC/x2TWr4RUfVAMMn4hazcMV4E2/+fwHw3fi+lRp
nZ9cVI0Ae0440+hvef8P8zsqp5tjH89v2rKqSy4dEzxwwPURMUG4nzikVC7EWe/o
f5/g5C09FXapz8/cMFGgoq1Q12PBESkkZdIw7v4KHiNzjLRfqdFiRLHc9r1qRwkz
xlntGsdDsthy3XS/tihnIqpqONK03TPCh4pdx69P9BYwazpIE6Kgfd6ZobRQLNJC
1tsk3ay4mP8UulOTSsf4mlgdX40hTAAi2Wh8lFvdzDHsByoevGmTkNUgNnTwy9qS
oLaOQUY1DU3g/F/aUFJjmmgbhnpj++adcMH2eTDfRDme4MUenhMS9DE+K4Er7FyT
PwTzM6wlNwWXJ58cLa2GX3HaqPsOmOxEaxwGjEq584X8ex1Frs2uKoI5BoMgwZtl
ImuShmJF2D44KJ3K25vkWgCYq7zogFmN4yUjYRSQdn7iGYlleDMPKA68O6GRnAGk
eKgdPHoDmz9UyOu02JJ3ls7RBZTcj4xCn/ClliuHSY3avKMwMGADRP5PXCwnxX7k
6GkCaDgoRXltjIYhon9m7ITwWWRFKXKnGQ0kUl26BqnsmquJQDXJcq8+ZrHpPkjK
CZgodRrlwtH/ZaWkxZNqMhuklIGRDKK7RMGskWw3XR6bw1mXJ7x5VHymFTFSfgti
JVCSgXzanB6qed8Mpr8Iw0tZx9V6bKTzUDXfsjVG/tT7gp72OTYgHmvvkPlHPQ28
0oO20YKCYPAOW3WxM4jGP9DFZlO1kzyJDZdB94P4yZKNo2ee74ZTdi+UEeXb1TJj
xqQAwFOZtKKN3Hk5F/C1LBBoOSSOrXjwq47y4xy7DQuJoFdL7IyuUirEcoEkeUTt
5md/3PWhuNFlQThUy2VLBmbE1Cr5UXMD4bRdbEEBstzUdJoTlvOyru4LjZJ5rhpH
QXbvFTf0V+PFcHywk8+ohSyMlVd7Q4JHaEgVrwtUXnYqtHxit1oeux5nUySQHWJ8
EuEDjBCWh0hfqcTBBfIAAh3DiRW7pMzCAmSLWX+CK21kDc/xIsh8kj6PAQphBq36
DJTHf5bDQUFBBFirWZHCTeR4LVNj4Ah8THg8Tekw3d0X4bx3daVUJ+V364EDhmGZ
VOy/ejLf/kypkI3BMzNhMp59z8EXBVUHovyvlv6O+/OEz0gcC63iQqAwgCxZg8NZ
dzzIsdFlxonFwc1fM6/at2l8bNaQy5SpzUmRm0fromnW+wA2WlWkKGpuQxehCI45
1NvFu0G6i3GxBohi1PqgZHPCz4eTDpwnJzi0CsHz+BCkGqnjCwnSAeQg1WcerSC4
QCQ94mgZohw+pYgPo7HrzC//acXD36rjziKNiJhdH7NlQJNIBVzcsHcLdPw+Y34m
A5icOYdOP2Hh2pEHc1y6jqbvFFBhIayzc8y/97oq6u0ZqPsOjUZKXj0wWT5vfvxk
KQtGBm8967emRx6F4FiQ6FPMeUyxLiPGKMW0JQsIsf7z4/byr5islfF1JccG6iMu
ouY9fxNQSTHCBHH8emTDtoRm2y3a59sYR3KQLziqO660WRtq8rZXcHTWzkQX7lFm
X8rtee6dfG/gf6enYtSmbLx+FDHgyFUQUp9bqZ9FTt6QFZ0qhZz5Tfk+ZbvtQSMY
MihpLntvOdY9sGubia+zt202NhLHE4DsM0BBP6hAy4rGZr98BqHm/0ylFam4uZKo
hU6PNid+yj3CElpyVo6zhyyIEpgoeoIx4eqRNubSktgD8aWyX0xet/zkrxwfyZwA
9SqoZBFC6BJ/lk3ObtXSpzmDMtsyQm3jRoeKQJ6wGsVbZjDIV0f6Uc+FmhCnOMM0
ZObk/EaJPxRSm1cFeigx9/yLjBLONvNGlKa+6W2XrpQ7N8QPeCG+JxmdZYTQBAiq
8kkIVCrviXHjC3fExb/gSc4JoKTMcGsVOryWZ/j3VrNrdRlCs5aiHFRYpMerx9ko
86MvUg5WpQN7DFAYIGKOW+oMzVDyAyf1BH9p2qySPiYaVpndgX+ZwK+8khxrqBer
wtJwt25SmE8xqEQvmHSB5lLIUAoqgPlVR51hGrlFbfN7Br8CeTvhv8zL8YHGPbrt
IqzQXcDniT/0Gc83tJg7LCkZVqkEQH/9Z9KAP7f8zEcaUBdluI1r49T1cmV7lrLj
JUkvBrf6xcjMkGafOxKxNuxQJ+Z05GtoGVm58lU56FVdUH7Uf20qEVz0qDXeZbkV
G0whcRnD9RuqcqE+spMKCn9Spxusi+TnRGv0RShkOp3po+wUPto4/aLLW/8+cBis
a2cx4kwpRBcwb7WaFUYc8Ghh0GVkxeDJ96rKe1ooq86y1nTNchRB8Z1HMSakCT7p
TtmRoP8PMCo474uvHrlDGq4dQLcZY9kEmDT61XqvcR4RtJG1UGv+0cUEU6wrMFFE
gOSNiiD7j3DPAW/g2zHf6IlbgEKsK1J1Jhp2rpLLixoIcPnc4pBmCAdp8D/mvzh+
6qQzga7L8+rv/LrjY2ldtnicJQ1uPth80YFHSBvMyUh8r8m1aOa3aeqvwiTZOQ4c
VhJLoe94hUrzHgWEUcDV147QE771qsF1iEgAfD88qqV9119FrTpE/XStxI9H3O2v
KYAh44AtdB5w30beXLnFmphWvzjeE2EaPpUHIdXDbYLAlYeRlS7NNHftxmRnLgGS
irWCBff5l9KY5S/EzUP/ZaVRzIEg2ObyVC7/9eFX6vLKILN8FNN3K0u1eRhpgLVB
46Ys1g+tFH1qbFD+kjpEloA7YajggEVKSaVUuV35SQ1Zg1aKt98nMw8vkO2HH7Hj
fF6yEloqBW7GByHzdzTPthROZ6ctV3HeORVTcOhBvyGTVT3U8AbvG6E1bkeE3tO8
VUlDWjLixuwf/aIRqDKR7hBd4Oz3APKTxqBvXbrHc3EZ0EXvFw7NSwpggiiOyhAo
rK2m5wKsRDa8gKhwpcXaNBwA+DEPoYJZhvo4UH75NXAPJWZUHtQmM1I9yaONq0vc
k3Qqu9mQnEzZwOP3Z1RUd7uT/hQQHKJlbxx9PVLxMlKDNVOSxk9costNwxpid4HA
Lcru5HE3R1/jhkRhvA5qVKso314g2TOvnz2qxX5IO4EKQySoz7NHfYPoqoGRjf4T
u7vNoPfnLzeJPqDdCS8Y0kYg51nzXDLaCbX7YyGTKbdTzc/yvZH8DZFBozChjrnw
zCswyUwiSYab/BZqHZ0wpXCTF46JmtpblHoZLSfVoPCqrmX5vrur+fK2rNtDSImq
et54tJehWDaql3MQZXPuELuCA+CMP1fRefr4JoUUZNgShFtHUhIce1Gbh1UlUv7w
5vIaH8cGkcQrSfSOtDcB/G5EGBr5g1K9f1t3yDy/qyoz0Hqnxr9q316j6j6kFwwp
yU1MiwkUFXxyJl0VBlshHZNQhM7w+9/Vp6WdjZQNhpq8RpCl/nH4T4D1nAwGhahC
2KKZjAasCs5hq0sUMR2LBUZYOII79zo+v8CfeXOPJOBxQTdxYrarS+OVWHGfKmNU
rMbhPtMcXs4jfALrnzpoeVU2w/xwhS/6oAcQN9ymYBusPZ4604vhiYwWTI3usMML
/AgF1w3t6V8beDoZG21FF666gyHsOSTYC/8ccurY6qE3WH0XrKHuUAbr6w7D4DLV
rfXGE9tS29BIq7KUM2uk5QdTr7IIqDhG3d/Vvo5WHtsD1UepO0TKgp1xuGFIiRj1
tLRrOC4qOOvBdzX/p7m9NyDEozqA6sf2QmPAS7b3SqJ4GjF8NYkjb5NZ4i2Maant
c0ViBBU42ovGaoV5RXLJIaYP5p3fJBj/T9hRAL93aFZA+ZoQaJflWKVqaSfZ+hIl
mTA8PCG8BycFtms1H+4J18xiDTv+4AnniZ+pMclcEDX+NZwKNAmtB4Gwfs1vVVO4
k+YSkv6wLQZmMa+83Zv5qhSxC0pMaealfDXst1N7c4y+scNLvTV/vs9uWUi4qCff
4cNSQ5VfGqdA+Pgawk2pEwm4SMcRczCStZfIE+6K2trN2DoYWFcPyLyy2yBovz/p
F56SgagvoV9tfy1QDTkFJQNEbaBiXs/eCcV0BbeW8nSg77ug3kI99i70BANYN+CY
obLyopK+zAb0LOhArAYXhqpdlqBkkdpodoV+7xhBVZq+kDivgdtJnoe1Uhw+xJVv
S56qrTikWK7N7AhANX4YaV+nsbtyryMa9XPivtXIox88y7RNJssCdIotv+zFs4Z7
DtIfWpKyJ8KEbz0WseVReLk8C41XuGi72ElFCLDJVzTEqzfW7p+pHjNLs5ZEyVTP
qUBDAov5WJxEc3ZS40affa7LWQIt4i8Wc39wr3uTytOEGeBg338iivzljGBjf49h
JKN5fUaHgYKlOt+0O+kYeLB+KYuJoGsswBU4uX0ARTugVtIw6F+kBJQleDkV1wvd
2bPZdKpzMMNB5EpRxI3qvomCE3Kbi8fx9TwymaQfOa15dTs2cP63y8Xn9vvqItZl
d0cieMFech30NJS5NCC/6N66UHoL7W5qbXS+M6GZPjEhDIB4aGrxLB/XMDYQG+GU
Og7BQ2dAo3ki6M5ylT6AQ2S2YFrp2hhXMiemoQH2HZ2ejlyvmPYX8YBjj9TLVg61
4JS9UgHv/MWRJiLTPO3nHNMOn3nL60LYGthhgzsyDiMvY7h4HqLbW+gfMtFDHasK
jswLEKaZpkbwgaIh3TiOwk3Agapc2hfmmYLvOstZkvMRZAEvMSPQ6FN70YLHrO5m
CFRtVXDksRDcItkq1DHNOsZc+r9arb1qgLZY1Mhpef9/j1trQqOiO+FbM6GjPuai
zZIA0SEpg/7fba1Jhacec1yq2kSlGJ0Y4VSoiaWIKLHbebxV0GzaPqvSRyXhZY+1
EF9EilttWDGid9mquOGYc6EdRcbE+IRka040RHUqubAOtU2SR4k4AgNDfTqaN7pJ
gsghNz189TegVUGCE4573qF7q/rO9t2iVZFoMozeJ9SzFOzD2SJpzb4qph0AXVLr
UKyIuKIZzQBOtYhC0kva/kHPy9DjhnMrcuyFK8Xth1k7nF9kRsQoL8fCse/KSwWy
dTLgoMTRd94fpb6n1pxdk/6bdEhqcuVBJ4tg8umzmylNx9tOiRt0G30Y8ODRN3pK
2HphAz7N1B1ObWlPtn0Oca4WMLQOkkAysNy+COJduSOB2xamdwFEUZTBbd44VDIv
LScRCk/9ITmtd8kCY18VE9+hMBTwg6Ztz3Ua3G8+P+gwf9IIlNDNnyAcJXpo1IuA
BxCsQcEuSp1hXzPNR/8JKefUyCnS+GUJm7NjI0Abj2bSXU5ylZ54xX1/mzqyqWI4
yUOrRNuVBBI0GU7gvq5DCp8pNGLu0EiTDxTKa48iFgXmWN7kFh3WPCoqdoA7gzD9
ilVFKj7H7vbg4dH40mzEa+nIKw4H0Mse0joQqJBnYXqgKeKscVM2JAGu+XaGj5sJ
WZza4t9mO9hUzHVgYKf4OfZMm2YpzK4onn6J5QNvqvl77bGS/JWYKwRnHq01pyu5
EPeuOmhGpOBgIsI+q2+TKPvYMVn9AgLJXC+as91S/6i7Vu9c5HZxKOFVxwqFFhyp
eB9IFlmQnqpgr+cf/5m3JGsA6PKmr5kCaMfAiE2GKG3wuFepPuqhmOAZ0yk/GP4J
/k5ugL9wMq96ILuFhcYhooGiFb4POLIfAOa0CZ8tQhnM9FhYiiNM2LKBIvD9RRyt
aMpk5x/FLA/3Nz1eBgwBKv69QyWduu2mURrlStaan29/qSVcRBytdeTBHOjG71Xd
i+CPGHMEYKWyP4eObhr7cYxbZZh8jnTcJbVMCTIsYIPZiiI9h9WvdmmHpLL33ztp
46NpR61+8K3JCbFW7M499aYkP8Si4OblCE/WUgdP1xgQ9DpHjFvkGtg2X3AKjFFn
VywgCiaHrIgczuKDRZXbAQZ+8ho5DBEg55/8e7NzBzWVpHf7jtJSsvDwgFLWmb8R
CfjpL3EVTsPPmDUCr35JKoe1FOoxk4iDh86Dsr7NPs0M0/RvU5bGKUrIxgFW+AFa
DwcQ5jpbSEp21yB6ladJlq/OF+90hA9tGyAbcqQEQrz7u8JESJ1c6C+MCzxyQvj+
+rEx7+Gy2WJHS2gm2AttS0WOb8j0knJrTwC+EqxPDBC4fcoAUi3IMiH3b86D+NRg
I/izFYLR9FJihJCA4p2H/59PwRnxKVnsVf/XLPv7NdCKtC7L68M/NJ0N62p749Zf
hAlNT1QfvLwhWuoyfjGtiaZl1Hpz0s8lPfV+EfrVa1wGQbapo0pr/aSULlirnBn0
X9oU7H5xi0dCWcBqeiLMHY60hWsN7vZ6EijQLMivKcA8vn9Aay/KFTXVFa3++Vi8
Al1zZtSRoQdP0WXfn/uAiP/m4TIk5AYmE6w4/BrSy/VY02UKR0IIosbsxH0bUCH1
3kqTOWHu3FQcA1DTxhggoxvohwUuE4cI/w/htA0EFIbsrRHEb3w1D5udFiK2bF4l
2u0QyuP3LG27TNkTee3uxbnboFgPwtcqiWk/WLNsbMK+bFL1NF2b3PZ3VHPPkacp
OWMjx7YTI229ndMlyfQeJDiE65BSb1wId86GRdu8xZrkYdnCDa4ZpyTfU6Q9uO+H
lAKwwncoJThDdvvCfFrDEckESDTjFOHqrD1JKR62PLZlS+qPuekAGS49tMJA7STT
2RmTyNErLT46PsdhAUZBSjvHbwDom7dW5H48lRmyC52y7xEHHNhOYQABJhkr2+D+
AMdgVqjoOQuY9wgsyHiIamqoduZlptBfVX0LbTO0K3Ecf0PIe+VOk2YUd05wzk8d
EI4rKqon+0K667nBrVcUVm+ImYfjFkVXwDLIV00keLf+FClUUj7qagzPJd+VGkvM
CTyg8mrjj9SVzA0oM7rNYGk2uH9z+EoAI8+jdbX8Nqm75r23VYqBZtE6PMavhj7u
hdv29WqQOlcCHoDaw0c5om7tv2ayxpkp0B6RA0B8W9gEv5ig7NhRpJ0y5IETc5S1
bu62zzwZHR0sIbVOBkMfXcpA7AsHUc4RWyzTxkbGXSwaWbTNDBlHyyGJLfD1SPBk
ewtszx2Ys063tDYm+GECAMafNlQtGREVxyH0Qyj+ZQVSTxzMtzA0p8wmhI/Z3cIm
mB0k/9+zuVFMWpJeuEtw6CnPdBsZiv4rDByJLS6qfVPo7jq5ChT1fXWLMFzVbrfF
dG83gAL5akDGVHWwzztbHguoriOfFOQMQXE7KroXpOqmDBe8nhY3t3FqGj4WHahB
6mGis6mYWq00rD2bLn9Fzu9/c3u/HIZi4n2x/Z8VmDQ2UtusGaAjfgnnDBrMONL8
HNyszGoKu5XF6DxSuguFuD3B9Z/QE5++EUDiSOkSqUe5EwkDU3458DUR0p6rTF1e
fjdjCF+9ua5ZdwpQLsyEoBjMMgUsv82oUp4Z+1lDuFEKzWAbEbhGpA29Cmj/1KOh
U8cNcyw9+ntXvcCwjNzqC59EBezmpSSWKT0smD+8Mb1eU2KzuFV54j6jlczMofJ+
M0DYzQ+kn1nVop6Ikn0cEgYwb2Rz6gReuH0XM2bXaBtsRVPXSQp0+SSe64BvVAix
Aa3I0HyMbttQE1qSKr817DmGkClYxTxG7HhopWaGYnTVswP9BrxT1IFKWrcOUBNb
bm4CWozHjuoPO9lPMpoTP+g33RY6l164QpLisCNSz4eEaXJjabZQkf/kjAJIhC/Z
A5I1nZRTh1Obu7ddQscbG6As7vaG+Ox61FVYenUSpwO3PLg/sfpCpvhKmS6fYm5m
729GNYk9xWzeRBP45bl1Dwl6lUsc8E5b5UrJIiygyiC9MQylMaHw+ctK+1KVKZyT
KbhY0iNS9FeSCoNOA/qGtm+XhQVeOsbUv7UeGe45Wpv/K3uVjmd+/xsJkU4sLvG6
lcEIAvG/UerDCunxgh+dlody+JdX3Cpf5r/qqglpF06T9SJI5zr1cqPAZbwoBP7p
RlFG2fVLeVOqJrVLUzWRPuFCkmOqhfk1E2pEaAiIJOcKQQnn/XAhetw6nIU9V2a2
sv534WVNaN/epGidRz85fP5jW9yBUByzKPPPoCLXriQ+xg9NRyXBCZ88DXCxroLr
egbg9FO/DnZk7N7ksigOlPlvmKhkLaGu3zQRArEnkHE2wrvTHJEEqnTl9xK6b4Rf
pFlupo3QIoxzAark1Dv1fkYqO3xQ4sGZoArX0yDrtSyrBV+HDVtlbbD8IAKmAmgx
ZHqFMY27TTSxPGBoDQxlbe1SJsnBmEr/op1wg1ys4r+2sfYRLOFYpPguHMl7ATUe
PjoAWFpcKxZgXuiXfUeoj5V2snOqAAZbz/gkbtIZ2hyhkMw8qBFOTI9T5dn5o4Iy
bi30SsbxTLe2u+CI8x02vrMKJW7S0eKNc3wwYIRJ66LPAyU/AAJp9dk/xFmsjkuv
YhkYs3NLpJIZbDCTRQbms2PpdtLdEkUdOguqULBbTgRzUCi1VMHpYTT+Mu8ZVoLu
ytTV5BeDEZDVfbLkI/cbfYoYAmQNW6LGpQBpLpus56r/FliTiYwMjLTmmZ/axlIJ
1nSYDERBy4YhMsbMysrA6LoiTks7LJmRgIO+jkw34jW9YQ8cXli3f/yeuscIgB6I
cvZgZQ/dPfp1TCHtHZLcNiKO8/rw7ZmvQwza4brewsAqAJeDFMaWRbKqouU8jePB
JmptGUZXd3HWYnJu6KRxcqFUIp22uC3HBS5BI9z2kttqmsOIwiDt0uT7cvO+Ihzl
xzEmyhFn955qZX4n+m8bVy3d+TFV5TBh+xbiHjMH09GsSMUpN6t0V3x5hQ63xSZs
t0cSFAENjo6zlAVML9o9Ycrii3ZL4PdnAZead+QPfDbLEA1w2rdps0kSz1zz2jYK
s8krEPO0dBhzQB1D8ZcfHX8so1E4YxAdLKjftISkZmf4BS9NNsejKuBuRbyEpE0K
sWqqzrLjaBjPexTwatPDfH8JKp/fvMbTp5+NAU70Cof0HL4MkQuxvFEzRUc9/Ikz
I/02kPWB+Gz7P6lMb9U+B6ahudtA2QSKNTNnQym9RX5Ifplss5uTszn444TO7mNj
/QXB80CvJki+h0FKWiTKf3wZPHh2raddgN31jgU5U+eGUBFEYkndH9S2YWyGz+wm
D6ceQc7KrwWBM2gDr/Yox5i2IICyUefZgwowfe9cN7VCuSWckjk3XOa4A/xpR545
vGsfC18MOIklOSmypRoz04tGup0e+1a5Rr4In4LbCJnvn4f7fu+A0nMogSghfpLF
dMAyjvhfGGG+HPs4ahVCQsbwZbiMKH3EsFNsVYZjqwEM5kcQ4fCkTC7ZYzaL82+R
kipi+kuX0Ue1abGCT4Dvvx2l4El0CSnFfgwwOc5qVU51yw7SPgcI7miLevXAflR9
MatvFcEVhtRyvSasq4tA5GTbV33QHGu41MIbCMkbs6iwv2qUJNuy13X6zv5UQgSY
YCP9ZF+0PvITNeCMddeGg7A24B6MyiR3id9vvbNY0nIC60WyErv4s1eZxfAmUeJ3
HKc1W/tRqxkihg/D/cRkRKqZXKy2DCLmuJr/0mbjizQQKVdw9NsMVcz/EqUI7/Ji
LySFg92IoFtl0HTqTQMIdeMYPy5KFwhIDbB6zkyViT78f1vM/gOEHsoa2rhlSq4N
V8dz9HWCVl5CdbrsYZhUNSCZWECiey9BwxkrQdo9zf9+jFdRsjKiwSP0vwAsOFoD
X8ouukAmWpfYg108sRHUunZwjDmhpWCHwoqnrtnbh+SRi3FZ/LWv2IRJ9A/pP1Pi
L9/yXs4rY2YC433/Ge5JE1vtSMKRu73aUUcy6B6I0M7goD/xfOPA0UQtLlbDTbZZ
3odUX5unX1RyMFZPXzOxCQoHFrd34Dmhq81Dy8xOxOWeplTMT6y/KwjGBPf5BSHw
xWZZD2BWym475Ky3EZY8jBnN1f2XVbZT/KfIOOUCeaMGJzUlr3l6u2Nq2l0tbmKU
/Lq5C1KPp4d0sP5MZnnTJRsbUi2OZKHRtYPBmKMrbVMc0oJSDsD2SvVMqqBq+o5T
xNwmWAbN6ewdZOxZi7Wck0gWzaVhQX5j9thjd8aUXLboVzbgmPGI4oDsZQeIehpP
JHKgkKga29Ra5yJTVa6KkvMXKk7snXP50awJWDFwcOg7DS+a6nhyURMLv77COsZU
7S8D0McnXjfmNq5WjefiSBBs6aRlc37a7aZBP0zM9N75qoWyo6PH3uBLrMHFMiHW
gt0mrBN+Q0v+e5Qd5AnXgvMrBFvKPNKSr/7hn/l7FWHbOTP885YgsMjNbAoDHDA7
xWXCuGABZoS7ZltLvJz70CRKqTAOlYwU7IeteeYgoyE0pMk/BZ79GliX791rtP/L
oHhdmU0ii+dcTRHQiqoJQ/mRMZWrHX+vMt/lVinmVYXy4dgJzji50gGbEP9TsBuh
3ci9jNcvOHtt2CX2pGJy1bBDYAtu7ArkGvhvAgQwNgAC4U7hTeKKS6YErfNjaovh
rBI9fhDujwSfJta2M1FNpmVbj2ppy3gHcERJ2gs3HwF4a0oGU5q3qsJBq/K61k5e
BFmGVmuJskfYJAhJSAZ4lyGYlVcJUwwO7vq1yKiNzsoONkU9s1JkZuiGoWYoUg2N
teQlumqqN7KeLDkot/mSR2h491zKLDFBvfF1TxXXdCGqz1WBSOi/uy9DoRn3iFfD
niqIaNi12wbsJ7HixpMJg94KftSFIQJswMBR32tYdcmIsNKjvQsQa3Ecmj7+LdyY
tWKVr7vtwnJ2m8y7BnO1p614TFeqPGrlRHwoxVx/x6I/+qlro0Iv+ECzP0Ozw0P8
FuOQ8+kONgkA6ZC77hnqmfKfEZLZK3hpDOrBcWaf3lQ/7Yuy3FPXEoX5WouHSZA5
1ueFTpTO3B6LaPqc4LHUfH6UVM6RtyaXmlZB5NuKwFV2bH52MGt5eGfcW2tmZZMB
D4ypHZGmQFrRnIHrkVIqJQSPibwAKUqdWyx7Qf7Pj4eagtboFM3QlpRV4kQfwzpt
46EbPlFFbpC+/DmsTbhZD1mZF4VfCmfhcl1K8z5SdPeCdGIbeEWbPBILkinjYSbD
KpsLvM7wQShfxT5KeseMJIEDxrx+mCQczBvQVpFYmyr2Y7+94D5mrRm15fecXOZw
b0s2br5qiZdsrpcd+BmE4zRSjCjYravGecLe6NMfCIxw7lPFJ+UzbJ11v2e5FVq0
JUdzSf8+Seh87l1JJ/EL8jEvI4Hh94VK2lqoEecBXDvJnkpb7IfWKf6Kb4AvOE3A
rWej5cGX0qduOdPIvcHMKyiwyALpDwHhFc6OGqBTBmRUjhRN3EYglrE8VoWavn6U
Fp3lL6opjxxdiNyCPx5pde8wOV/CuLg8e9Gm5Qq4eS0J48nyxbPUYKycNSXlqr85
oXwhr7uoD9hC63mh5nabb8LMk8QGWSbDKkSinNqarHnyRFL1+jN/IzdhRf9SnK/l
+SRAz9aUnLSKvSaEKhZwNlF3j2RBI2vlSip7OF03WcefoQF+/AP1QJ4r3Z+soW0I
Y9G5gKXQpLkhPNGKhCLt0LzXlbuiGgGuP/R6J+2mcnN6H2+LlaZzeoO01dIeYwF6
UrsXQ/S8sljSkKQeZ5+Um5uRCK+tGcnNe+vr9mxDZ8tkoJGlfxziTT04BiO7/XZi
+fWnC+xaZ6OpKd0CVKXlQOd2Dar5u3/MXtnTC+ffkglcSlEyRTOV0qX0vwSeXNkT
E3RSxW1G2VNxdiEgxVCSoKXn5kwbX+xWm9jFdU4omsoiNQ0Tj++XfizHTl3PpvtN
zNn1ugNMefBWf3QC/9wt00x51/14e+h3N9wDMXotxMCZvbjDAg3kXkgFdW3lvN/K
VNwkRwW5Tirvs13NGNVMsXH+pLy9V01o21/QEXVDdsR0oMYyX7NZ+HRq/H72UiHT
AHSOVMYt1MFRY6QVnY9kDMC5WjHQ5MmsomO7PGeYvLHeo7tfDwCqAybPsEm/7yTH
iBFQ9eNP665Y6onwdxUMZeuKRjW/rWiKfQxPiC5zfzUgjYdLAiJP/e9NAc3HfHuA
6bn1y6KsHFsbveZbgz/GLyh5eE4AvkFv7DqY6Pu0vsvlL+67jGAhVPGrrV5/VKF5
mgvcTi1x4RGIO23V52qmtPGwQIJjCk8b1RBxTL2PMLY57SkJUZ3MLdLMPfkO5DoY
eaEeciuyS1Y9eqP/F+FeIazTut008fTVDOHSHUpgXJIdRU0SLs3d+UHK4BFy2sY6
rbyi7tSvlx0FWFTcZgl7WaAXzMTk1ifI99M+L+d0VxgZvWW9ui4qKH1aMyH7EOel
jyvDwo5eeNo7/5bx8uB8pbnOWdas4ks5ZwoBY6lSZ5ixgpnKaRtSaZTBbry79/BV
G4hrT/BZB1btBWHNppI1TGi6mwieZuanUaUt7qM/X+88J4NTYNkkXjStLhMd/0ai
2vvqKMx5pE0mZQZr/oSlzoMoAsHVIV2OjhpHC4ZDnvlQazAo98INQS6fDyHwbkw9
yY+TFOCDmgXsx1I3G7Xx3QA1uTqpdyV7hF96BgCazPjvR9d2gNSr+J2kgSLZjWrp
sxLFjw6MgjymlZTScjzFMPZ1ByKUsmFKDWXfBAVFoNN7J8YVOlEJ1ScsyvfOOobw
9VMVqr50eDfkGSBbh01+3cQ9EVh+YYPzujD5QKqS0mffcRErxFDFnMKwHw2E2QhB
OuGmDGFv9s76xS6M6YgTEwaVErKqv6WR4qGZWiFZBwvMIXfZfIDS6dcAdaIVkysi
L0v875dJKC3KKIJsZxjEhh6uYvDyuveoWOk4N5ee9bkiVdBET3jvrP7Oxf3CtIuK
nTnVWx6i8PpkjB9VGGvSVkwhVD6s774nvHUdpMpSLpXtAvJUs+nG3oyplQDe0KJU
m7jr7l7nECtcm15Sce6c0ALirfEx60n+pfA2Fw6flsFJVKtTdjl+XIeL3HLlPRzL
XLDyWwwgqLqlMuuIvX2McjjlaZrSzEquqPXKgFLPS86sn87pPUPndS3nW9Pie52a
YzBbgUswVM1Rj7075hVzNlE8NQ84bIDSKEVjLXp6B2GoNY8o2uq7GlTulKB1kb/f
mtuBo9Wr8F0/pBKwU2u/fshxvonnJ+PZ9+FlzexcSN9+kBIS5wQy2HUbFUJpOe6x
if33UY8l9LkTi0+H2EvST5fvJ/KmJ8DjwMkDsB7w+f247aA5mnHXfkHAAZprdr2s
yUiI9nrv8bpB5WDOxtvxkaP4vobHjC3YBgmTOXApXgtt+FUD1hek8Ee/uZ3rgcIL
IV2Pb/VFOwvt03j9eEyFrgn4XKTOCsa4Cup0yJsayLFVR5H7Nut6FrNQn8U6goAv
jbRSNTECRcALzJi97nEPMEh8h8oLcbz5wQt+qwuHONcikVQtAhoz6zPXbfMnFSe8
vdQoRz2mU2FQyyjjf6N7h7Gr+4rU5DfbZZbOY5MPHWTtE0ebSi29pT3dCdES/P5Z
9dyK1Lpdahr3SC0WFyXaQER1mOG8FeF0kJlYdDHm/51gRZKm1DZVzxnzHr260AVZ
3NZDPaEOJ4oRYLDAAGZzln+JaecqSXedBlVxypSBuZQgTrqrXt8TQuLud/9eENrH
Wa9jOhnB4Uk3LAaQa2UIeRmNRT/3W4mi30WRVuUf85NbtA0SILjHxMc7kz9ctMvQ
AP/CozxQ64Ytc2dMWUJsGCvmuqG4f5G42sSTHEQuVWKBBd9Ox4B8QTYfR8JUSH4N
x8L9LYw6t9WxDbGaAUL0h1BBvBD9n14pcXiQE1gTcE2Tv8Prb//+vFWl6yxbIvgv
020f6DmsQSMesR9N1mDGM6PZQSYirp/uOkt3fS50HIy8ms7cd/A/R169qzUkR7i2
T3ksZIn/ElS2lp4nLrid3B+LY/vSUIGHqnyomxj6VQQPO9I0likB7meNwWgBPFeP
HS/H+DxiP5fwV4FJ8cMkI3tnZDLeY3OfpKOBLHbcAEyaYW/Quw8a17RajihJ5KXM
wTB1la274WYUabDrC/L/1Grc/t62fmiIq1Jr5Z6FD3i2ycHfvtzUbLsY53L2fQoG
hStWIYef6XDLguZusTOBOheDngj1UDl410xjd+/O30sMyp+WqjGGJt8daNCwgbYE
jw/dqSSt/8PdPZrtuD77vriaF8MFIqMtioFVWezEKjfkBEKjabunIdQQqC23mkyL
lt6A7jIrz7Mjt8vGd3JJMAUQl2GImHltFdtLT37TBBg/VxI+3da7tMZa50Fwfedc
Ar8gvm7kcGIJcGgkjKCH6+hSflhEtEkJ0ctQI2U+u51jGXkRsXmHlLi22R4NcJJ0
Qu7lzmwAXGyawCr5UWZ+BoWyTIZRLgr3UElu+hu2sv3cWlC9sEtgUK61K/iJVRIA
dmkU5EC4YSztCXvHtrvOMoLaTp7WbIROI3iyn53hh6Qe8r3/3fLCZFs/BoBlaU8Y
YJy0V2uC3yUb6YPfbriN6pfEgHwPJbqoEC2+l+LuR4zWOfcV9djIjRsU7ENF88sT
jyNsz78gewqPTgEVEqbyi0AknEyduYXSxyXRseqlEndxADPthjxWpt+TmKLvp7qv
nKqWqA73Zz8GbD3xh40nTKu/nENyCu+nmADQGmnjhHTb3gdgaDcR3/8JFrkm5S1x
cx4xHwlEeX2nMqF3Yl/HNZ3eLtcKPTVfiK38ImtVlV9m1h7KK2PzpyvOhS0FhuY2
FgR4fFUyQe+rdw2WafNAd64seCr49emJ3ZwEblUf0mQKvyJWEC7IWOh81uQTMa0B
oQ/J5dNJyOWnIG2NSAkpj73kVB1xcIOEa5aP072dELWEfrshPmaaFoU+EKCKvv12
8wttAontUCVlTVSSDVJBRo6NP8/2Lc+3poi3HgWXLwKcnijPYxAeuFlIqkyq8TrD
PdTcVmMUAsXc6WqBR7I2YpoengSkUj+vne4E0RY5NljxTEPMSENltKQpsLUpvO5v
8H587m4NpT+KiWJyUUg1GW7W4sGCCTPTuiUC73TEJHO/FjTvJ+GtqTUJVOORiY6v
Alqcm2ySv5ZfU3PMgmNZXquV17m4ckzl8b5wPep9TxQGH27zxJbZ0oZu5nXi3FlR
uaaMILjYh84VOkmzMOZdG+BqHUsivTyud9G2FHfQBeF44PBgZMb6xhEJUoCfNZNv
GlwyxsA6+HKb7re214xyDETu0NoMTfMQMMoxdLK0EvCz3Vy3fXrtunpTocs5UeiJ
b1WbLwel4mCW6TmOH0cPKNxdYNxe9iDi4gyxN6MHZu41BTRpxueJ5AXZmiVuuey2
OBE3eguGFboFeUF0o3N8JLwbDicJ62ZBMzhTMwPYdqxMsBmoGgSKFOlZbLtfkjSz
dHxFkvLsZ3o9nU/3ZbVKkHMNgqgJIyGomfiCCpNr6CZ4ngYx5Owq3Ae+pMahovLq
SoyLIYU5y2NHjTOX6dQYjJZ2ghRa23GBp5eA2Xz9pt0elJ1UvQxyxuJG9jxT7KWx
n/sE77ghMwCwfU1t9vcVKWE28DlCe3QN65aUDqrj6XyNWxtkRCqDeeZ5Umm8NFsh
eJ8ZlyBQ7IlDDoc2K5+ZHieKEa1Zevj1bGPtXWsUDJsbdeR0HtWteHoPJbcQWh91
8wKqtg9JW+sGZxzFv6jYXyY1dqWJO7/fZSBF4423zVnRr2LpbIy8IML9Xntm4HXp
o8JQHKJA5YaIIbnjT5fyRbI1/0KpQGpwaVps+i2HjN7hpeYX81pa4EVHDrVtoW/9
n6s9M34dwaE3ysUpjV+qlcaW1WY6ikBhf+x605jKVDNZtqPBeTBnqFpFIeoUJhdw
FpYXRDl4GrnlY4hW/Lb02heoefstfA1+dDWk1oZ1ypbtOrfcqL6OuvicfXmuRLO1
ICPtOrIBnhMUD46CXMs0EIJSxCF2/zqZel5CvE/T3Z5X+rzD0KixJCBUXuzcv0r7
fHkgZPqXB+M05lpIpQVMK9+jDh+lykSOmcYXMbfA8yLVTx3CRyaNWw1b+XNQljRC
ozcIYT13gFbkigtrqetHAwtbtjoiOpEKQTr7+8+/IgOayCATNVhGgqr64b5DJgUi
wgALCBwP+LByDtKYBvvE9cq1ar+gpI2gFzO6MTvXlCs7jkMK/W38R4TU6orb+G2K
bt794G4iyOhHz9rp6MNnekzUAyymOXCqsmQGAqYmCyXMKqsP+UATMOzteAM6XOVf
bcxpA+IpXRKb6i4/Vdw/iAhlE2+KQswMhe0bmp9y80Cv27gIAVlDXNCBhwCPsbwt
iMJ9P1ZGTjd90ByGJiYi7FDJqhNU9VZ3xQoihMZw45dw2zxrlEIweZlGM/PiX+0u
1xU74ayXGDWT9ADG/b4nTT6thn8HbwayH0GUjpkbmYsxiLuPsVdmgcQIX8uq4yKx
qWWjdTvB0uRomDBpIpBo8jszmo4DJoDR25NfvxVHo2ulNnIQhLTujrsq5jHQKZm0
cqOXTc4VIs4AWCWqwKdjV0e3H5aZdD0Rwjp4hJ2wCGFoXPLfNcIQ9CR2zdZL+0nL
smMZKDSkzf4BYOuU0o9XTanItyKZriVcNnRqdVAvB++u2wzqn/bHYq6kvDypHWZY
EEqjTpgZdeBhJIOrz0X3evdd0+5Ws9C6vcPpnwZZVkVqOn3Dv6p/8vDdN++6A5AF
TkCQdDo5hz7szLTF3Y/Gt88FlaFTP9ixQ/0qsqEFCXj6CAIy4AJ2R3hUTm85H+oM
zvEXvSpCtF8auHFH0jPuKo4JAFDSASG/cJAi7IHnG3Q3+jiPKHTLKpXsvsjKpsc1
X0geos8AW/pD9YtckHMafn9vbbhqjAkTMlyug8cGhACQ/B5yRrRzsxxbe5yLWCfx
qn6ZNEBKBcniIkX9B9VLY9FFM3u++vqFeEdBgwThO9ARrCX1PdMGeVJaFP4/cgV2
CNpU1r3I4vStoxg1tY/+CznKc2F3EXpDSn1nQlWXyAwWOnXiSqk7IhRVLCQx5I97
4hxUMsTvaqFYM9Yw2bobkxDGYlBs7dnDg4xTg64j9/N6vgpm63GtCBAEfK/HfO0e
ZQWj30gLrmeAk1ueB6HlU8Re2uDrXxMdjMds3/93G1I96hPIkO4ad5qYidAbl4yB
Kv6MDb/eis5wqvFaA8a/s0xlzEyuir9ZLOvVKOJrvfIm4POUjuEAQKCZa7/sBfAT
dOFxx9tFw6QLq59sN7oay+sjXn0UzOFhyVyuPiCQLd1qqBY0HO7vGVqxRAJaDmBq
2xuy2GbKHf+LHEEeUxOvtoi5aHp2oPWH4XNCfdqwybxZIr63S60DyJf7VgC78Ton
7LMSP3A/q4Ab38+ea1LDFXoc2vDjcEMDvc+W9eV/7D82e5BfEwQh0t5RO66YSftK
sTUbsZuyEAjpq/bjQ51hszjTpRKflAXwnIzEW/pNPbvFLSotzMy7rS5WQ9gyCBk1
+o4B0HGQ4R9O3379oBZYCtgcDtqrtPI2V2/Ka/z60142qV9NS0HsuqAmEsSCGv4X
kpa8js+Bhp/bR5EdfyMaNXpyalzz11QPp9c9ZSZxx40hPF3xDOkOXiuIEDBgDfCn
33g8al6JWRMlOPVHvqf0S9k6e7cNP4LqanCGQPVGZlBYjVas/B7Zu9RwFL6wJU6z
RvR1Tn0f3VTo1vJ2VsfISCOgh8CgHjX9+VKC98NTABq78/MJKSNsuZQa4ZTb/RRI
PHGAARXv/BorZsZPoNeRq/mzJsRrR3fsP5PcfpQogoMHOka8pbbvOjxHnNDjTkVh
mkPBnYh4ogqygvQsFewvbR0GJxsoQyh0Pjx7rb7N8/x9WrzEtURgk8O3TK5V/Ioa
iPqVeAnOiqGA8klJi60X8SBux15beDRGxVhd5KuOJqEhTiX+BuriA1otst1FYcxF
KbqQd7nuJ3jecjltJx9djq6AeJYvPZ4kob0NlzHm5XnSB+7XhjrmrVNycx00pe64
0XgdDUEveESV3CGs1VkT0I+WbGuTNDBmPmacf0MiKJpS2vObImlfmbJvrRshqON1
LhF1qMbCyDy5ifeSUJSL4EIBHnb27wo+hCEwZfHjzYopexee7w9ZZyMYx04E2EbH
Ww0gZZRUgVbeidHNucM5G5E4pY5mO62I1yNg9/UTGeVd4GKfIHYjZDVChK3FPqr7
zw7gtxe+kg0mVwTj085PJ+YYKJLjvyzzfjuNemYQVP3a5T5dy/Hv6GVN5mTT/dHI
2IAaFQsUPeVibC2XvBFQQ3wk/D3rE3zUV1+FiyEeRAaClPYZhFrEDKEKS7QBT1iR
7EtumUB1pAX2Hr+W/tU5lNw8pFbLi3rUi28KpBoJFCNSeOLJyP2eFPJVleKvdsWF
7xIgshNnfO+WlMp8/izIn9mtJs9Yy6qlWsYG1PSJI49tnDQVkeWHScpfjVmapApb
svF1VuK7QRsJ6REh0RLLeUz3rksu9eZkMJXaZWlteIU++jDNItZEMBzlE6k5CR4D
s/2MQh8h+o594rKY0iIPmgzHKHyOk2V+VMHoagB+nj1iqRGEfur1c94EnFnebCpT
3rS67NknmaFS+v7BvRSKWd3bA2EnaelRu5AK9qq9YUxzNTJN7ysR2hdbsqzqF+rU
cP4ZKXq0yMGPkNgMGORhl3xxBLsrA6VIDR/ZMxYWMzPA9jizfebm6jH0isHrtHju
gtY+LGkkOdg/RSk8Deus1N/79aL52g8uzGxgpMCCnO0zkjMLYUwZCgUY93h9Vsww
J3n0SJelFeYUDml0AVsDGqJnqGVShUeEAQ5fha0SEP2F+qNkMbmGdC7ETX++CRM8
LZhJp7mErBK2r8MXY+qDLtfBj//ghI5yh411wrdMn5z/lFSwwzm+3KqGsamlmwpW
droNFj0hxndmDW47FDBdMusuM/bZsnoA4XZScVlZNQcJJBCu4Oa6te/XZV5Ywz+G
m6Jh2DXFkaFnNwyEQczIJ3ha6fYyRctlsQIJNE63rCPoe2LEZSmRvTTFockNUFuE
nA9QX9+ft3HpOFs7KwEy8nKzw5UqlxegWfbeIPt66d7UDxC+BEmr2mvksApUdfDg
oQ74v864f7pT4+d/k4VLOxbt/v/0QoPuYEqGN4R95xbrcRaetqceC5q6xR+sWBNa
1lDU0DnP3eNsRgCGT1UNl0BftcoDXbZnS4Gk0bsddgt0UtKL5maWL3uUJwQgV7kG
CiW+HZ1dtj1ou+zROOdpAhpuj0eQ0COCIGLDjBvQknkHaehU3DnrFD+3ItucmW+3
YBwUneJZ6xqRHUZCLAOPU7xTo1T1/rdgLGtO2ut1T/HZEsi5EGfCRqtU7kA/2drU
WIP/FGCNiiD+yLybMzN14rk8YVwHmUHa/ma9L7sJ8e+XwHIyQMzoTng+nUhh/Z8u
DwezvZToA0sEN6rdegjnyOD3xanJM066dF1pa5Y2N7pvP4nHO6ZY04/iB2Csu43e
Gf5+KrtKO2v+nI0ZZZfrSa8a2s+sJvYRsXe7HHrVn0lbE6WvxSDE+WeAXA/y51ou
8COAuGmIb3c9/iPKIlORT/XePqrI+8xpGpm/sSaNT49pfZaeT0lMKvGzD5TTTh9L
rxpZfdj2EArJfUznNvCiclpDAM2WAIJFq2paPVZSZLb7rMx8pFQl8ApLz4scZITD
Zza2UKilaqH99G/r4dK+CZ2Wy7TUCocq8b+ODvHn/ibFttAV3vEY9o3BDnmJRpH3
NCaCvdmmpEIQt79gkkJZgsmjJIpR2xO5UdoBnc0nsPvoxh3Z5ULdPDQbGf/dS7mU
4U0Nzuu7EDurKBAiGg4Eu8hu8zQR2oqo/gMzKsY6ofObh6k/PE7gK/6DBtyfeu5Y
SoWWlM8WkdXcqv6vapx4xL6VEDr0Y4oYo9LgTZY1/gM0sdVdN2ra+qQEZ3YQbVZc
HVPGVDV3GS4l97BDshhcT0rspWGGh3CpzFUZ+s2EUAYwJ/UDTZhp5/mxUuvFRsFb
fuIvZBjFHcpIzFjDziqoWYXVAQI4CTakzj7/8DxBpfQDZBaNJhfbnndPJOP8qZYH
Fdfg2p2OpPLLtk9k9gz7bsqwDA9anngi2k45NCqXCpxgQbdNUUs1YfHrEcXd+jfe
g0hUJh4E9do3IJgubnZExMB2n8fXw5UnHN8qlURLPprfuCq+yyU7dXHqIOsHPqBT
wXQ3nSIRzC1TkhHRJgLjO6Ed++ZxyRCZUR22pU16vsuygJyzRqYsE4j4WSKkhClA
3YYPrio+XHOUJeOFcQ7jcHrabXJyOBd6aHkGuJZQTbT3bMkb1og7x4uCILdKiX0u
8fRxo3t2fC+BE7JsBzSvLNO0D6F60OHTnF88VevNc+JhuXke5pBXf/Yw9qFc7nPR
vM1i2peh3N3yvRj+d7WKJ2FeebGQi9Q6028hSwGvCSWoeEP8cYs60axV4FBmCuTN
1N/i+P6OGPbz+TTPgzn7D7Eapur3MDkhuAKdHG32Gf9+CAH2+mlpXsxDT8MqgYHc
OvUp35c7NZhabFaxoHzaAniBjqkYgJHbJQvzoQaQlYV8sXCPnEgk4lyVaeQPPN7J
KcNi/OecXxF5+i/lQoijj8Mk0lUAzG67n86A33G50polebWkAGeW15L5oVp7o89f
vkxGqN2seBYqYxgq6OZXlC/ZRGxpPV9bIWHRa9a0CEv+RjX5yUjfBuJyzV3T1Xpj
sOWhrwHHcYqY+H8SWSwCmgnVryBaSurqs+n46qT6egtK20BtXm/Jm+X+7DpGheF9
RHVGUKtuCzwef9xi3p9mLDZS/9sf/M+CjMrwUGmz7b/5yPqY9Cx60NIfW5IKohYT
zy/L1e/5dbAmbN8L8f5Qr+PWLUSXHE2Y7IMBOKCVifP87H7CtMWbfEEU6AwmsA6h
2+I+eRLWVgP4PpJViv7jz9QwpSfC2sBLIDqZJZKPckK6zPHzKCKZxkkcJuQNVpht
mUcdmtQ9h2r6ntlJMJUBemfDSMPyT0LIGbtLBd8E3lUyd5AQyEg6IDUPTTiw4Llo
EJjovmySPpgn0wF4lNoY+IV2iyP4ypkDW/2xsN1uJEojlJ07Jd4Up88iR94ubY0B
IU4CMg0SIBb7fkdkKLgJVGeWUL5BWQkySFw7C4dT8k35T2RPpl5Xf3+Yg87X3ORB
7Xk0oMUmEwaml1snJSdbmwg3lm+wG0VEvqNeFHuJWWL6PraO3VzRQGQj1QuHuvHy
Qx/eA0gzbZURIEe4Q3/ZG2B27LXbBusOQH1cLiYcW7SAeOzb418lQIN4g0v1A9+0
xnpcAQvNdsbQPWAfltVrciSuP8kE9Bf5RjeuxqI77xMQwJZY1rIMVFG7hxGts4nm
Yf45JfB+SN/dVBz2vjkJKLmOniyNIj5rFMMHNsbHrIlkbTduTPYWFb/c8R25lrAU
xSqT61TC2ERFfIiBashDoL+WLx9eeemUTL3TVTblQ8tZb3qZd5oHKVKzltm+ZilI
2G+qQTPndVulExbacI5iX7SFGa6mmIDBYFwpePKBWi+JaUu3PU82JQ+h33zNYi3u
FdvQfwVXQOtR4yxpQYLaBaZVKCWd6raN1BmQeypT5oZoII4sHUOTqPLnG7X8Uy+t
rJqjI814G4Clbi2RWaiq8+wuhI6iY6ksIhSwo4aQaUWK7gFJcOwL2a82Qqzz07/H
gz0S1uvfryncjpR+9m/C1olBhSwbvef20fXFef1huOZ5QDMo7XZhj2cX8K724pSk
iaqANreWtPPGkd6Z5ODlsZutAfoBw48Au5bqDfQn9zwCyGX7OKlwVWbMNQFLLlPK
52UkbH3rvOipesA3fd3C9+DysxZ4I69CwQP5DQHwiWG2gQRueHm08M52KN5WzwDT
rcgM7gir3Odc3Utok4UBMXnL0TSTBUX/aqQdDSibHZArIrIsTm001yOGztZ91Mox
eke2YxO3EMSHJFDGlKfur/s8C4L6qWLDu8Sbi2ZRf5e057ohaYNqQcox66DD/Ryj
2rxZxVkRHhUMwl6IOJ03DRBZHRNaUzFnxi6NA38SqDVUBVtcZoEsSURAz9d06Q7F
pqgRoMsbK1w68b7XzNuxQO16VXVKSFK8z2rLeFVfJMkxfVRyeOjrBq2uP2+PQuSz
IyrFTCpBh/shkX3ZPfb8gGPtFUBMc+zPKXOGydE0mcXjDCNyGkdZQD0e02IWKC4M
hZsGZF8iACnhQeTVqbRWKuWKmUU5CCczW+fQXS+OQsTWGgMMPZDKAb83WeyDuGuZ
+o+wPyop8VPgtVmiU6xipu5b+IsCdINy3uosJtGuekN57DwKdicXNA5jmkuVkjBb
Aqiap4cJnfkIc4gweCs5l8to70N676UDzISmbu19nzmuZHo7K+fnYrXQSYRhTfZ4
G4f+ieNEFY6ofJS3REzCjAYT9fgy3cPM0R5obGn4kXVU/IwFcvSdG+Fmmr9SgDHn
jLwr3D8fR3mWWPTkfc/HpjAEtAP0vipeZkqVxRjrZ9ugoM+k9MHLi587c12nSETW
HwATXc/HcuorbiJQFRTJwbhl15PiavPIBfV7hdBRbb3J7tTqu4RBGMl5q0tEMBNo
ibm9unDS/t8YXZE7rIDv1e3qyEDf6m9xCUeyruGSeECmgrEzbxy2jxd+frjcTUhl
9+aK14uyjW6g0a1VIJopT7suP7SGd0hQOJbVnvOP3cYylezCswSzLD8oaAX8ynVs
5leViU0stz+qo1oa4bVxcfxM4P/CEADSkJFtNElYc+7l3SBxn2R6M+5jr4uledmz
15fxrRF3IAm0ay80xOHa9RRYgN5//7gfPCDQPXlaOpgIIhFfVvbolGe2oDoPvuep
WLZQUrrWTW8K0PhH+GeFcUB4RQr5rNGylO8fKiyktMzBVzc6mqq60yruQ1tldpZS
nWwVUv5DKuL70TmTCU7lzGXVNop+ikiBhzsa8Us30xZ/o7ghyxC2x7QRDljd9xgG
UpLSczSYLPEvil0vzon37BFTHd8gP2T5iOwd1zaMrCt/GrwUtMRP20zAlDDKckKF
V6wWygjcWDHmDEXq3wdN3KaB67VFxdcQbW/4DMGbMQcHyAFdyxdbPsfXudVK3lHd
I+fWDoO3RuQEPkNnvJi7jNTlrchH9VPmwQbpXJDrxO83Rk8YPDfIqiUTg0Gwf3Sq
5PMtR8js22qijMmo0n1p1OSXo61Q8ti/hKna4Yr7wXYEmd88hJ6bkfZLI+4YquB/
PJanGFuf7VJ55EeFgryM6pTKch1EbuUw/aGKyiS4AdOzvg0Dv6BFluJojE2AHBYx
jWKGHSNFgb2Y9b+QCWsiFMJoPt3sbaxF/Y1iG1DbbbKXrOKunl38ML8q/MKgjAtM
H2u8Y05UWMvCdUFw2J8sRc+kSV61/sXpaipOl3HI9PKGRC4jUOecv9yHWlqoFAAJ
RzLdsjpO3PAxg2urK3fpDUTb9vcXyUyjPE4bmNhxYoIfS6Bg3QQWakv//I1rc18X
R4f5VSCS+Rfj+88Wb8AcpbzIbd1JtqLPDL+msZsVTyEKlnIIs2FkdwvFVvu6H0jP
7YOGcEkxNeKPdtYRBWTO4iXCA9UZ1z3PSwgLTcSTE5v30quPAMoWyvAdUggEIZ8z
UuONtpmI80NFfDs6v8WFCLksUyGlmAkJeIJIlJh8SGpKItrh20ZfFCXWyRy1VBBM
N1u2+mvotaovPFwpFA5m6SWVuOGHk3ju4gl3Tqv1iNkGRUP9FpyrCFQ2oFLOx/md
LJHF/vjMmDDp6inUPdjrH5qmnUnP22tLm15NBbpNrMTZHLjGrtU2wzPGbV9hd9eA
PkCErhiqGDlOv1+DRAUMAOAe5UMqrA3EpqPmRZT4iAOAoIR54100rZZ+veShlNhO
pZnbN2Wkw89IFOiYlL2UZ+OYzSFIDVj+MqcbrU/BUqQ3F2KrRf53pY+0qeHeYgOs
RZkyJe085wCJhxh9SBmTieQeWyTjDZuObz+K26R+qP030dmeHKAlkk66tcDOe96s
uYEQOJyWQHUscXIBQQxEVJJwRcCQcfY0NDULcR+K++gmjRoQWORUwYvJQ9bJE386
3TbSzFKA2jX988X8ENJxC/wCdvp7hjmQ03H9hMnH4M77vS0wobbrX/rNr5pbtWV0
QYL2QToOqg3+rWUzYc1pK0x0WZsutEguJB3kZglvTeSr2sex6753xKXXx/S3QPEe
F5G+fHEIASww18EIplMhu50JAUxxMDcPqS9sN6QRm8RinCMn5VFZCp84fK5B9sTq
pVcr7WW+iR9O+awfemcinLiRgJC6YJ6v6zTqd8+Zfd+vHqGS326G3OmxauiifIRW
Bq4kr/W5GaCZI145GzurAAw7XwgQuRdkNjOntfzikZXiskB1hLNIYRIYaOu+rm2b
gtWvCjBVxFmaU1a3ywVBofgx+mMm61/7EvahTr5qsGc7vO0dHlJzO0IRJqBEBydR
+7L1yJS/S228tmiF36zXZUaqmnx/VXR9b/SZrKl7Jpx3Zqmcvzz1FJcYIgp9HFFh
MKfZ7V7CDfd2idWgYhGFZVCsC/0Nyu/BBbmJ5v/J7TcvSaUs+ClaJh7QPLX/FUaI
g39i6PJUPReBMIgG478jh3wTbEKuPQXyZ163rZbx71lkSWYFIvJ8P/rRlvCpFh+m
jan1FPrc5DvKFvpkAYVqlBtW6qr62aPI1bEx5d07gZL6r66iTSaJOY8SJTGdgyFX
fHB/GthM6jEQ1ba6Bl+qVnbzsCXAmbn51yakC0DrlKopmAUMPMQzofevssdwnrdr
x5ukVZAfsv9NpupSusoUhAtkO11K0yi/8P3bfU7J+IYBbEEUVCFXsQHNME2UJpgy
Eyuug1353SVyqDQn7xc8iVnXwmGaYEUSWdpauUmvzc9aztdtS3ndg5bkM+wiFg4K
1K8+AlxjGbR4nHASxD3PEbkTkWwqKvR0TtTaS4yGw5zHKtrEMGhtOnK+pSol/Kuz
otKinNoZ+ope6zhSyScmKjtGQpK1mK2RjZbsTNyQMv8QLAnP2NonGy8WcVL/wtCX
gF6adDqqRokSFujNOeYl0UA21YA5EdcXifUqmUncUnJfjwWpidqnGQbSNRTgkUGO
XpjukXoAIF94ZNEtncUrgVFgHWRbK63dFnTjouuYS70FQ8JLhdggFaggs0Soy3qu
fHakcyj/WON6023JNJrBFLKMjD0h6JpehRGPGesLGqaThdUY0PwiIWwE7hOVwg94
E2Bks7GCgAN5LON0pgYlOBmo4NKJvqMDDFH+yudqmknmMqIkcu818sn62jh1VTvu
dKm07ItsctBXv0tYaXXOmJf32Jdl+4Y/E28az5zmUethHKzn6fn9Ym5QUFj5OwlC
sr8DsIRl1z+lgeS+BgcUeDYEuss5CPON6RlejGoW7qJIFLx0D3o/VPCCBpydQSf/
HW7zb1WARcjxL737l4CYm8S2H01is7+9YwO9tdftg1wWU5P844z28luKVD1LrnDb
WHqscLvjsWKCwUyaLh1fAwNVkWjSnLqLNsJJXvauHl6z8A9yzVecBtnDA/oyqAOY
Iclp+MQFTMhwoBHmLeMBvIg2cHCqEgvA3FQv4xzzLFyserwRHis0CU+75J+SXgS/
zOHgsU4qD0HzegSC/RXiOfIpyuPqtqXZo8y9YFHxny4wOQeBRvSPaiL32VBCXfV6
k1D30/8LgaRRcgYdILVVlgYBqRatne5SwLUFnB6g4ovR+8DtjcnTWhqL4mUkCwh6
ALwY36DutOx+yX2fxoCTLIHQUR8tOXlywwKs7UUplYcdVLN6Gk6kd4sE7kdGIPgs
EWGrLa4naSToeRBxfjT9PDmmx0Fxz03prPDzPdCcE8HdY9NZCnZKSFJQKeG5T+3w
qMN7t8dqf9bM4p8sFz4213r/t/Eekmk74A4d+W76Hp8ZecUMxMia8xlSflAbH6wJ
xlN1bc2k1YyPj/aoh9Qcdau1pYLTckkj6n2YaREqy5JGbM+HDiua8YCAg5FiyKAu
/LEciTkSds5sY/bEfVOb1LAs/ikrAQLCy9QROFllIfB44AGY9u67bX2AAHopcyKe
j6y4FJx3pbh/0uarrU2917b5SBUfr1ZBwiqTf/5gEUqYTXBuWPjy5noQHA9F3Za6
4zgYeKjULkPp7tvN8vDKn6yDQuJ8Pd1GsnFem7xOESTU2D1voKPaVbnJG4ZI9Lit
IJk9j1uoe0qhnEDib3kZKHKykZ7q0gCt3khALIwgw3G/1XPgRCzxyH100sBkj2jH
hziZlszo+B2qpWceoCFe+xLSp6Y6rtutAvJ+pracVJyNX8nHnm+HkNjTWKIEFg1g
8KvdFB9uP0xIpTmk9w+ypxjlFhG1eIZDL+W9PYDTEwAZLRh/Dgqh8xKfHqZwNwdT
CX+g9bTmDhaZq2N2tfN4n9XsrK3wTGCSe6lXdRn8dO9IrPJ0ZsHO8YGmQ31rIOK7
W6xPgq7HvfEISWaAlHbWDXDK9otgE+Go40yZH1xAdaoX8j13ZxlXnUTxTwTaYPf/
owujPYhOBNYIbAIcNr97yJfUl+LeTZLS9/ClovE+d525jvAUTth+aej8/RAiGEK8
NlAzfeSHOABhSzcQTmyhECD12Y0zS0d8uEZNmeN9j5CRO5u3clP8jjlrNai373Lu
jXuqXksCT8QZ3tL2s4whRq/NDkBBopvI1DHzMyti9u8eXBnEEVAqQC2tqXrqlVCa
fWrpDsVfUUzi5EGSj0w+s6Fy5StxrSh4pQDFgSSq21WeEgTpPuU0S90A9bJ9ytiu
urJprDndUznacU7dExrJLC3x19oMJY0O3lj7oE6mZ4upbT/C9YPXDhK55pC4zop8
9eDV51fyrJg8AuEQtGiKgo42DkmKDw7cFi7c2Hrl3F3TTvRBscHLvWDVfGd27ViE
7qj93CaApalt02COXPrjmoN1Fq9kgX0Pme4xZcdKr/IETBzK2LzQllLhImtaJZxW
do0unSAW+hyLZVfPgY1Qa6h04XNbx90p3sQppVUQeI1ScHt/TwBzi6RlwK824rsU
wsSFP0qor79CWcnVsEV/wVw1pP/LHOPIcICAsE+Q9c8qa247wbRzxRU+TWKUce1L
fsWiNvrGJZGPDw39PoEYDBRjDD8kmW9TFvacHkuTSjGujxkQIUG8DLNF4P1JrkG6
/zmiazgBatUjwv25bj7BiBfvE5VAewyV8MVn66A+4tthI2/6MAkkZC+Ua6u6kJJK
VM1Bec1Gczb96CbxaHClFIOXZ0GbZL6RoK2SK9zIlo8pyxNmYMXN3wH03gbTMo1G
6aqOBc/CSBTJ2j0xysQspCqcGQ182O52rCDRi3zbfg9Ft8O8HDSn0bobB67E1EYu
TwPc1FB3YAEEUMW6rlhny2OuyuJDV5PHGqV/DjkZvi5sKeWUP9JNtQCEmepYDn+H
Ea0ini/ld5Mj76A74OIlue80GBR5jhLdh9ILzJS4hjB8YPo9g8OWuzJV0T9mGA64
OEDLooes34S+bOmbOX2TrLAmXGAbq3MbgLL+pES84m4GnE6svFJNp1z5V7IBhlUB
Klwv4LjPz3Mnzf9rAdA51ER7bvrJHBed+3jti+2fHOMbWVY88apeBY4e8mN052Ll
y/Xc7X11L7vOb18ET4uSN2Oh1k/6BtAPTL9sTTSqv0YZ5vEOfbiJeqqiA+x8drFq
zM4jjoYIAkZsKi0pZEqRVVM1wxqJOBX3GSOh1wXKiJUuhKc8lJiPsdwUKgQdDgJx
CQ3kZ6VK2STCbadztdD4wyfPR36eQS52+5uWLuHIwJ6xE+rfAT071QzYRrMvwqsd
wbV9AdgG8HaBk9BsVTzNtXOdRjKaI+Okmcs5R3bHw0+6c2twcFDu3UBPEBBtDxZX
dflylSnrC/A4UawJ3n2emWou4Sd0lVlbXkW7qTAQkZXcXOKJ/tt7Eer8UPA7YF7t
FtiztHk4ELqeRUuUR9keTrSOtcaod1OviCRBwCdU6YW9ULt/p3lmA/3Svx32tX1k
5d7XOCWoHGSfDUm+uDSYVn3Nqb7IiKk9295X/DgLfoe/udlcPxjbVLQBiCfIN6r6
8Xk9P1ZlTAuMfuycO/gBoe6Hncw7ftXiIgR0E0/zZT+DpJwVdAtixDa7LQtqDKs/
gmC2eeZ9UBwBRoqHlqpdH4YDQlmU7tfXwCMy+rDNBR8cAqQv/ra9Fq/vLrLLhab/
UD5Mng3WrXowJIUNpRuNe2DqFO8USapWfup+dq1e3UbpzAJFuowIWIaXXFx+ze+h
LOEXc5I56iWI7/ZzAy6sHhX7lnYDu7eWlyyr5RGl+Z4e/Jc1UjzT6TE1TYgh9yaT
3eu+v8Hf8yGjxjzLbHBayYl6zbtrJ7PpLwBFAYOIMkm0LOfz5a2Jbdk/V8yIrPcA
UNyim0gqHviFxe6aRw3yIkZsALSWcOMj0TGMrwh1Bki+TeYZfQXjSS0o4et7rVMa
IZ8Deqv70RIkdvsTADhZMH+7C5S9BVZvz5nQzp7WCnX3DkzESHrDraTtpfrEdpFz
inTQ+NM/+KKo+xh+457mTp9DXl3S4tgzqJy79j5Y14NvUteN3jyOXP2kodv2JlUT
X8zrjOm//I9Y+m/zfmixGxrhurnzCEe1W7QuKqIXIavpSArGMF+qD7dgE0J/6VAq
QmJCNHzmajseh6STUYJyiPIEGNWY9wJs8F4oOR8aWdslNh4+u7LpPYs9xE42qa97
NKi7Hh74RKoLa1iRs0p/xeLdJot3H/4I+iHNw4yfs60btVPjDPbvWx8KODpy6k/E
N9Tjh8wWSJ01hDwxvfEsBfFdcqjKD2G1d4AGGqHAk/hIWmdhwDIjyravih1+e0Po
u6yQDQ10W6Mbz1q2Rh3h4gpqcNX0CFutHGDEGgid8HF6T6+fgdfJ185vKxrf+Bc7
Ez4vDosqbDQkfkHHjjCMDqLvZPIUficgAsCFDMw1L/qYviRENRHL0+fdTAW+Jm9D
6nBejm4y47zsrGM0Y4zyUDpB93+LrmMEl+Pu/0AGHGZ5WvO1FwwYV/XjUZwqO2Wl
RGCCehmKwkZRgejgj8LXb7vNxQ75B1YXtWbhwozyUfsd4uZmpIBYtrlPBeImi6o0
xHKphRXXOtWiJbf6z1DU3cAyioAwisiMHepau2Z3nPYhaYU70cz9v0Ev4Y+sqHsY
dKC60ouUcRwIsopBNJPcE98gdFTvbSGmyJdBB4yzkBE7k8EC8BRlKQrsq3ajDFNv
KUndxM2D9CoKtPDD5fqjAzHRJDQfMsyFj4Bge6xgtOrcnuBNjXtLgc6itbInSATN
REcl919z4oCm0W9xMUO+cNCeVI5JWuswvn4fr9rO1vFVOx/uix9ere6JVHQ64W2W
ldIH/pgA09RzZUi1wAtDkXNZd2HSDw0NhhvoW8JONUbn257ACAJjr2b/xqv0VcDm
D1gfCSz44+LnmcHhJxRtvwGh5L8ss419XXx8RJIkPdmjiJiRghhJzYMqkYOe5k9W
eONeLUokfMCxUV8ieY3bJKjUzqMhVz87NRUbBi1PHDAJwbwxTLYhIhjDaPQcMQ4R
3oERn+fLSZ5ozHEQ/9dDji2Zrq2QbRiIi6EWTfHRqJ5jlz8CcPDKVTwzwaTl77/j
DK8B5As1cp03JCA0i5XCToOUFbTKyIJtNQ6QUqBATXqSzgYvCy7rYjDIz0oz1lGx
24TzvNUlBErLadFdCNcM+wto88YoBiPwjInd3Z79oh5KgdpZWTOE85znrXpVouNR
3nGAzFaka7g+ZFxTwwVoJ6p9UG1f9y0pbz7BRBxD1p/CunPwyLuBB1wUFx4Y4NWa
kkbCpHUwJM/BSXm05WVJ9tv5KUWK1PpuZUVP+qNTfL8O4T5RmZER1NueUhZo59Pc
t2HZcSoosPlJOWFRPZhy0CVtp5AQfzhPDdfWlkHacX0S9tE1QY7amub765vsvmUl
Kd2QjWWXNKdP4imtizxB2lvgFUe+ye+EFTEllsFAiZm0nnsp/j6YjXBl7Rcy3ncj
/mcuEqkQL46fykMOsJWCoGDykxHWcY1czB6yhoa70/UBxVA8d+FaFHRkrv0xZTvz
BzBIepE6sjSx6OyxeHVPjpSiY9Fpr9cIsT0ZEjuSPGS3ovQpBle+kqRf/mxsWY2h
wdNFDP5yMtPq/m8Y+VFiuRxCjlYuCPd7HDhHSztgp+H95mvhc8q2Tm6BkIsKpFXA
hMRFqhe8OHth5JplxRso46x/e6S3GPJTumwWTa/kKQQ/GLQXWtP+uRrkGkV7BPfW
sAYihzUxrO10oV2BxMhUcQ4jU+kRZOgMEPVW7q1F0Uf63nHVs8Yfy2yqKjUHPIEb
DgQ1dmEs2CtxhA81ai77xX1qJdvUnh87G1o8DA2zd5fZKWcRsPjMiJWCJt/Lz5k3
mpONhp+RzWoUye0p4PlVkB5Bwn+v8dyOPUF3i2CeDThPVFALPpiaw996yByCcs/I
cQCX4IQMhLbbz5ceb3GNlBSt/+dO9CDo/h5SRdx2ryg2BTuQ62c9aaJPc1apdQUF
EMHMTL+GaT2TrhTU8ey++RwrsZPgiepDDlyKGRP+gjxaNJzoZrjylCPtrSYqzvYh
La8Aah4ufwdlH9mzW2NtTj2QfXilRTynh/7uHrP3ivkzA3Q/0X6WEMiPM1IzMThw
rXOprBJXZGnpbKhozxYbY+n9uzhwPI6xsOUBIRyuMS2nBW2k5ak9Reve/IpwfDYf
/ih+GPjzCJ1aT14vG9BSlr3UI66DVFQ4jtnvx3ghZgj7jOy7k/WY9l4+5dodaBz0
kIXBGY5KQmhReD87i5Kyq/lq1CqDb8WAjUjPM9STIrylLHoycLq+sKxu5SxWLJUd
STANkjIT20jFauyhZr7ULfA3eaul/u/3icHzZi/GD8xn/nX0KaDGLa3dCHFGLIbu
BhNlYOOQPB2O+3NTDRKAlH6ETUr6j+dZpcY8nk3Hnmb2KPGXyxmGGV0LOWcqN2uI
z0SfarKzh2E6pHCuO2/aXaoufr3/YBhzG3I6+sK8YwNHhTvXQyzWz+5VJh9CGMuE
THpDZXh6XVXH+WhZR/2bDfKJ+9HVpKXQ2K8y6P8OQ3RRiBjSZpO3gGZE8wQyUtAy
tZjFxsVPUxr55bBHDo/GBDntRUTlZVd63xvI/LPLdBCbz1hpxrJmAbn4S6qa6izA
c9Fy28gLgEH2VP3lWIZhE09t7PFxpkWwMHvwulDDzAUxNsQuYCsnppJRCFLPhPx2
7XJH0HfKVfHSlOsiBaQJC6lmLln8tETJvYsIIdgoPFYlLCBtXhw8oUOur/3GsRYY
BrKitzGpHx7HFMKrMX6BEhdVJWMgSnrM9AIBKNqpdjfL+ENclisQdmJnRd99BsZ1
V+i7iaWURE8uJz3SCpXi6bWpotyCNcOpkLiVr/DTiFfeTALQRxNFLJx7/c3cKE4X
AcVBWQmpkavLC/4yFbnctn2KB7Q1tOv9j0ZfMK8PvVqg2xBK/M8iyzz16Eon7IIB
ycyRAo1cj5DqtyzNlEXHRi9zaZ+ISgibpiUBI0afDP9Jj4hKUTY/BjiKJRDf7O6o
HERdGA1Y9kI2wmXlMcqaVVhLZSPIbuJWexZRYh6azc6j4elEtjPtGIL/B1plTTtw
pXBAH2BZfzDurbTC5t4NHJkXyjmmQN37Mak+8Cz04wf1OnRpTGofwNZ0GGfPsc1P
Mo3LXosRCVHHMEfqblRhksbFSDmGUk1A4aUjXwYuSkrT8CyxgofKs4YCW2gVKQOU
bjiy1ZercP7sr+1bCyxwlYVLBRF7IxMCg4pv77kKAQ8TSkg6ZoYeS2EZFmuRm2vj
X8ozGCtsMNSJpi7y9EEbsGzNQHEwneL5YPJ2yUHAJXrsl7InVylzX8qKJC1bpvII
Hdeh5jf+k+oE8fzaPc1aTEW8kWq8KlRnrgpKNC3cFs9ZZ9S4XWn0rpFts0vqZe5p
fv54P3DoojsJ3tx2KOhXuvhgR0Ulzyxm9X0yyKkRdYB9Y5n2AEwZ3CLOjQWoIv2W
PmcUt4DzM11skNtIznTt1rJrr1mMmz/ZlEwh+8l8WVvjcMzHtkEtBV5QU7SAQGx5
JVuudDPXLuLyZPfMhltU4ocPp3ZnuV5yNgH57/wYzBRenixyUMopD9cDHlLN9MWT
AAcF1hpluCcmv4iPnX6RdZp3zpL2O7x5LVSwTEYG+mCTMxQbOFapyRkApSyFjKpC
ieWjifP4PTM+T9OCstRsi4ppQH1IJm4mZkOeSY2DR2/bX6Tb6uFhcRcXnp4lHLDO
viZCjax86ae3S/Hei6nApzEWFZKPeSYYGe5WwyT5QOAUr3andYGgxZi+tGdvYysy
bTBnV0wyX5chbJT/DHC13/gFF1uigiMC+7C16BYvN6f2RCJwppu8f3+73PCLeNxz
F4bWshiKWG6cDY8293RXHmeQsfEniYEoC8sa9dAz2nQfXdXGvWuerUdDJ7evBRIt
9ykRo/hyVCn7mS4Y+JeUF/eEJ44SonQ0fOBmG2f2Pz4aDIIlapjbsMGzWPjRvMQh
EcdQqwVDRXc5FzSLbeXT6r6E4TlAja6NXuucGsyuctOSvNxyBK7Too8MBG2LQ4mk
bMC2yakWhQXJZCENDqXKQXS7c8/CpyEhP/9r7AMfEEEeWdQwONvH/r5tNeJrG5Wl
HeH5wwY5B+UR9ALKniGOK6dp6VBZA+vn9gPuaELGFCHStZ5m4sulfHuKr1I89qSL
5wIzGaewa0BFjWzMu02yeBiR0yBP0aEbMoMmDO6rmoDvLgYfhT2lRcxhxjVNvOGu
f+y/8PobeuWVoflsNvJ4T5bgiAVczKdm1lxs+chPNGoeg32NqLZZVESFjZKZ4aRx
pQ1Rg1lMvMOJH40L4jhYFvd+cfbsRKYnhOidIIu2ByVJ19Fo49zDTG+2U37/zHDK
TFXnKadzFeZWIs2PZxEScNSQTgJxj5sY9qPw8/XcIrYEU6yysly6TAcJkVUXR3im
jC2mbr84xCYt05K9I/AwE1N+ACUIuCtcqKo62PyDNjFLoGyZyrfXnSZV80mglMMC
yfyoA0mH7GLSeUXTLFNlF6G2Twu5DytHFu2FmDskNuDNw9Yk9FP4iEKeFa7PFkJs
X1CaxgtS2OK9PywqM4rU+VnWicFOutMBmuPHHOoZFrB8oZaKUxjaRgkrJ1WOQueS
OhcoC71AAcL+LLiFeOpJ6bQEDfG/DJYaKWizP+sWXebxH4P9QAGjqnKbLQC7t3gw
CH7r1moO55JiQJ/8lqDVKIHfwciOMYZIToUj3kz6kVHzRTR1nj6vgHCfUexqjDNU
Q59QEqwIn2P/IoxvOm128Z7vsV3/Ztzpe33nQWpCEVycwkyb2iHFekV+cjxteWWV
8ov52sstVo8veFH5yHNA6cArVoB2HUoSCL2PrvA2CEy5EAmKOO7qOo2xOhex0sV3
y+yFhMp+TB9Hjnh2exwNzr/CO0ru8FV9GI+k5kIEMRffgfZHx1pPdE/AwnQapXj6
cz+ZmEy1Nr29tdQZLpZXgD7RT1kWNEAQyr5vq0pRGd1c5IMOHWn0wqYDLmca2VuN
YbGOh4sNzCtbDFQyvFH8mlO8tLp+yIPakF73A9HsHDjPBeCfdpsC0Ix3dUKXs2wx
AsbY1KkNZINr67f/xsG1N3bG34NvY2kcdioxCmvnUXapzUhoLnFeF0+b6hzlSIbD
y1Pq+Y51NujklvwR9/IWhNRrmGKVKEW/cYeKcS5WvgrBuLH1hrInrXRFRjvOPJZf
pAqItIgdY/fJAaXWtEsUOavGuVbMLANemzJ2t9jNwBy3lWb8m2lZTmGroZguqxi6
NVAtOh8Y7P7hFUsMbyEnOt/cbcJmBgUvBPhNNB0/BDJq13AcQcWLapKb7aoCJmMx
z0xO3XwYmqVT7plxjveOUym7Scdv2SFza5OrJEgWOubZyL0gqnBALbGlyPuA5M16
Eeu9q3EMDg6/S01IsUN7d5VwLtbYunFDq4mzXeT9MWPMxKISEFKYA56N2mbStDQI
7DOUId7MQLSS3lrBQgkvgbx7AWQdDWe2QPAWMObimCkBf/nv6bVavaFcPLWAy0/p
1g4dzYlMsnDvbFYG+Gw16DjYoDSBrP7Z1wAEMGTaya64JuTVz3O6HyDEqn4TyqS5
sruGSXGKLjLDBBR3AmYjP7hzN2uKF0F/G59zmfYFPly2P2kUFcIzLIUfa/SiTqdv
v89MQWqtAJ553fcdsU5hoA1kYAgaSwqJHBCDAtpLNQPcw2uUZqqwID44ulxm0bDe
kpK6cwtnYRVwol31DAAeTX08+yvPtH+E3ZdSNva9G2y1icjFFy6mZtgLLJsSLaOy
SFXZUhdql1STHhFK2oMwdaxActAVew7EI0ZpGOsFdK408DEqQhq51hVZHK0WnYeS
c4tGn1ns73Zbo1wbD/2Fvfrzg6Hdyg2e26844CgR0ppByz2Xlzjqh5AXarnQx7Iu
Vd935mOm2h0H7CvX765i8ljmalxjnpMYjRnbk7FelmTVnIPy+PN2jEtnNAJ1vRnE
TyXgVDqe7QqC02N6LDJ/Zpm/n6AATeOL3i48htzpikWHkFd2e3Gmd2Ro9fYUGWAr
ft8i1mHgnoaOpvBmoPNVYX/vOI3lWIBb3tu9Qtzj6LtdempnF3QT1Qe0Bho5uhQ2
f+lUUoZuWOEMXkISngA53KqD1grMGJRBpZHS4BNAJRqgwkXUlBy8MTHz1n/w/xLp
rnebeGOnc0eZWBuARSSnFfo/PJd2QIgZuCteMsgssmzPGgX337vXDpeECBAGuDYq
GVO9M25wlkGi3D51/poTaKF0UcitBg6T50JVYKBMYnsnuQKrEqqWmx4wgDG5ZLtb
6fQAPlFd0p3/wfdK9So0r5K4G09wPVRktVG0IVXsAzOG/8h0487lxPq6MYFjuADj
0lmQ5pQClJ1xV2f2vsMQ7GZL/3e9SnkFg6VcExHeFPvFUUqwX+tDjB5ODnN1yhLS
sawMp3YRTsFmLQzZ/sHaGOpi9MLPjnjjJyUikg6p0H7RnJc9E7XoaWTT9I5agcMG
4WpCbeZEoht6wBsXtJieX27KO0frfE6iCNdrQvarapJhy+DRjRjZ0gy/jCJs0Um1
plumkfR32hjd0XoEMrGs1Visajfoy8c2wd2rPvdW5EdfmancVkO49d3zWeabcR47
n0wffCrYmmIIEmBURpuWHtGHejw89Dh3RQ9jo/WNNf/JAWeF3OwoKRAARaAgb6ty
MJB6Jy5c+SyrAeAVoLW82A25plKxwYLRYur1ElGCMSWd3AEP8QJuEmrma33pfu2r
xiKlL7uTkRD4q+U7Z/4Kh7cW52ylH7kStofvvD8Sk9QyBCemXA3PsztCt8RFPlyk
uAFdPueU7GAiuMjX63L0WSMappx0PfL57eiV2BIj5CocCzyoDCGHGxtfkyjtAdiT
+NGxJqH0g9Istz6kbsvf2bYdY1DSh7jq1Rvn1InLqnn1cMRFMmQhyFqNzNW7H0Vm
uvujobG37+t7D2kQtvyR3hEZ5SgF8EgoL7z9nQgQ7r98X9ObgW3wkpY2AQ39FSCs
Wq1rhoFW1fxsK3Tgs9vfSgnXBuXwpI6bTCweMGtYObO4HUKJWJ2Mgt6KUgKGFv7m
ukrT7gCFl8BX9H15rbS2hdyvkZ//Ig8oACzeo/4qMj673vtUxq4qH3ZPMvj+GVRj
RKPTB+rMUZ9D+y5AXEoJChjzxq5i9rxkwxwl/+Jf2bUG55Dr9sXR5h/rQbUxGGOo
4MAzDnKReeaXUu9jHv8Jrg+EZiT/UzMelftw0o3EdxizqIG1i8LUGlv+2anMisRx
NuPFtBoSPNnzZaYyISR7JnUWjzSYvthVeZXhFZ3HlPWE8PwgiMA7BWFfwedyjO39
TK4E2QEs9antmeu2RoAfboO9B53NWqrIHozY6n5Tbdmaas0ER9jNwfC4rS/YDtdo
dpVkPtgCZVSqFbN8tZhUxB0SyvJJCSiNd7hBcbz47Ip6gqvZK3AaWiDMzJuURR/0
XDh+aacimXXCFILv8jrrEays/F9q9p24kQXNW9AxZqaZlUMuRglHtBMJcwDRDjyp
tuEgqawhpexkYnko5ZMD/Kvr/RBJDdELWVU9I0PWpgtAUAUf7es+3ftrlHHn27VN
xcGEEJbxnHiIfxOeY08sHGGI1ljD8/SdfGg80SbCkQz21+yzMuLr9rkp6DsD+PvM
dvhlAwhQs6ZRweqZH15YrxWjKtr1i+WCI3V/6+Y9YLwsQhrx1OOXlGVcds5yQxlO
Zrln67PyA3iKSmypGAsXiChXEfZuSUcyRou4XiP3n+CplKD96wQxysSlTZIwvFSE
NJYtUuWmoiGb5xgZIkcWcFJuK8nFUW5IjkasWItRsYo9BT09XMRWEiJWZsSJ7Dco
RLTCva4ZHE2t+1WFO/qvivbzH1v/Z9wp9debidGXwrgML10rNZuVj9aUEvsJyL75
gXevwXRptgq8Jxk6wDQIujpak5dzsEQc03M8l7z+wt1qtscabYWluBgFCAVn+9pw
cB31F4zEo3tXu++87llaK3SxgA8bjhKEU+BbwM42p1NEgKVI1Fc8AROEZiOEjsRB
mSoNa5RKZ+hu2vnTrKcFFpweg9ripdxIDv9D4rT3VDTTzRUFhG5AcnvxncN4L4f/
hSeG6elzcO6WcxEbju7Glh7dLK95eLFngj4gdkGInXYXJHkrPfx2NrGkZ+bgiIRG
NowYPuo4oywAs5pBK/jQuYSasVu6ll8L/Re8VNxCb40BlmTvupXF+gkupQd0U4E5
TkX7yqMNq/xi5MpF95rqK6t2oKXONKdDYNBgjoiBThp5TuLAijUU7hq2oix2uX5Z
HWsCdxf/q+xZ0+KmQb8xrVffT4jMPLExPiiMMwruH7gAnpYeDpw/mUSpOM1sbw+b
UqjyG2bfMankFlNIShCPwgicCEgqpWHoD7MpW3Fw1dGhxwHZCZ9teZKtbMMDsXMv
DpagFflbkQFWYzQkXPeZezeQJNPQ6dUlrzKUgdZj5YSjCVZHKBNNkh8YYRVbI0Cw
omg8raLS1TWJ3gJkJKpmLEy0CV0+w5QbXjwYEltVT2cJ1LGxW1rAlEpBc0n7Mt7O
zdpyo7QvPVOSnsllCBdwVcnyKbnTToYC1yzWanBMKp8/PYwdM7d6Hrd5theSFptB
Fio3P4MFJN0yBJbivbzjyTxSkFkxnLe+70XUx+BFbWuLlsFUHNolUDbfpvoLAVre
+Hj3EcTHVzLbuaKdqbN6xJJjDayRsqva6o/Dv9VvEzZXl5/NKvLQs1u/I5cX/aL9
KGbL+frPJlsuFLMKKtVODB3eUUUOwDWRXwKzXWGSZUpl8iZdNYUakfgJNC5/tetm
kk9/kJMagb2qbmVi3HKlh2Fk9hizHz2HUPCp74wGygxnua7ZUXtBCo0XV7tNezBt
+AQv1LqmhBo1RRcv4c5/YW6C+B2fVBcVMCXbzJwv51ZC6q6OChdkFoHVS5Kvs8nj
W7vDFyB3DqfMlECXUDaVEzimacmvuHaYIZL+YwC3qeDLshcCR2oNF83Sl9WmiQgG
E/ibny3jJHKUxGWN/vMkdAFTevPIm5OKk9kCykpP+Or7rkCDi5ux3LG3D+5uVE4c
9YXc0TPyARyZyP7pgPYyQzkHRDobTrMyTcVhCLwTFLi52gn+WPDsWpZg4WGSeMbb
xOKAwx0rIWIiiDjqJFgHJUDyeLbi9E+k2C1BjYhphjU33u9NM17zhUl2AC8J+xlD
YHD9KxScqsmUXS1PgFxscWk3633AfLuf/a6V5lhoJHdEaavhPkFyJ9+RMqgy6m9s
e/ZZtw/PO3sRGVeusyiTzNNXEX80JCCTMff8D3QnLv+XRBujmpMwercVMEudn5HA
z4q0qbLAyuv8rC1kYt9nfoBg5tt/9B2j4zhO8N0V3dfjX3dBNzEI17ykSHrd1ukm
jnk2JLyDLHDoFVVqfswvJ+reGpiGDIFjNxSIC2ur60jzsa47gjks/v5VJi5b6a6o
oc+E6nHn5nwt2tlJQbkZTJS/WLCTGQUjyabzbC6SlEBx/x+wGcQRVpb/j79A75kU
y4JztHvmrrsSVgLS9lPu9g/xj3LqLEVztplAGHlmNJKLbzVmT2mettutZ9VivYt6
91iFxsntkzJ1ySz8H42Q6HyhW7rBRp+rRs5J1x9w/4SE+GipB5Ain635iBxrNNB1
YBlCiDJx7+5HK3yDyc/Orx7Cmg9ZIIebBUFAKefNgibjo9Q8Ws568Q3lQaLcm1JM
O1tVPrJX4vumCzGmSLFcvqCmglvt6nLrJhYMB8a6KNkjoN3ESGaQNLdlgf8+4Ljw
URcw8sbimH0X5d1iXmDB1BzbGRI3/UChnQ6FDsxwWPBIoyjGbsO8MbgqYy/buu7c
2zMCLRhkgBveljmBe+H1CTNQXICuFSQGBdQH8IsfmYIsFIP00oLgKFgw7165IEoV
+ao7nbUuxI3GpecAKFH1InKQx1xBxHLIMjH5VttGE65DjVEkI2e/63C86hm0T0Mv
SyCptPvDD1QIIcJBcIEWVPAv7/0qjmAkE1qin+rbExVSt2Dum4KH5sp1HRWvA8c8
jvHgfmj3vW/kx879/uaSkDdqVf8RX1DqS6Clj9fLha+3AoVDm25qQbX0Z4KmlhoU
TwpEUEbUVDNS8v70BuhtDMEC96n9+bNHCGqOR41jbMXTEubtyBC4x6ert/V5vyKU
nE9wfZGm1l/2yYS09ds/wsUeAPSWqMgEC0rblt/dbhTzjJPvQRemU5nT4PfAnxF2
pEMHa4Wt4IxgCBUN8VG/1n1OsDEFp3roUnZ37wH7lsJ1l+ia3kGCko7YMkTnI+mG
T19JpS1cFVFCuYCu+H1THQCUUJU/HxiLD6/ryB/yRYDAFioVi0xIJqtNo2US/Esk
Pd9b/R122lS29S1GkYgYZMbfoS87jBB3PjmfUup4T5k69HPwqFAa19eHs9SDhBhs
3/rQ5FPawU0/I2fwTjoE9/vETZVYUPBlfUWM3XfhUGoOXjZlzBqnjQDPDq2w0mZk
AbYhWaEGWDJE3ApJgmLJywLAD8RuGdrAjGzzhqT169NJI1UT5144eNjV71Q4v6XV
UAaXaMm1l+t8Qg/j/kIFyZXcTJkk4IqrL2z/aC0eUGL4jadniDvL/k456/Xdwoto
WsxWFa59jl3dk3OaD5nebZT4T+eaiiHIkPsLdBRGhKNPnp4dIRp2SsIqFts18gZh
bk9WEnrgEkOtj83LKfGprOU89nQI1b9tUJQBSO/HRDa7dMXVgYDSroemuciwRAjg
6tJikrmWON2ZV1LG3Hq3SZgPj03Wgox6aWzcJS2BfLfxI5Ul1QTy5q+WolN5I/+h
7klGCWsWAKDniAIUzjDZMv+AXQujGELOM8+DD2J/jg3WH3DkDTsFLLEfIZ8pWIXo
uUacM+QreabI8FLhvPzXryPYnXXV/BrfDWol+yBo+klSXps0mLzAB7LbqntFsZtm
Ttr4EzVNf4t9MgGl0IBzWFdcNlRfU/r8ECTHbICM9hjUTq/GgCsuGtCILjZNGZxX
FJCOXnep/+9RIddXDqrzj4XSqD2dvXMGaIk3I2FpoiuhYCEllMP+cDbR5o8FHIVK
yg3KNmRtt4NuRp5MeruVShk6I5kNWzDvn+2vZRdAtw+TyaZnBrKTR6zCyXdeNTfO
7vYqwbpRofBEGcc2iqn3ZFfxqCHfq6t49ItQ9IaePdwyIPH/PFB635/EI3ie/R9i
eIsWxgA2drmKMiEfweFFBmEFGGq4r0lbmVW6aUWdHavXKryxreNOm8X/jIlzIjtc
d6894d4IszjV7RHWErCfWoW6Ljp1Lqvkq1ild1J5okkZ2j3h4Xdtcfts4y2NT39U
xnkq/SS4RT+0K6U93vhzYZNt3gA52PbUSSY+/6q3zCdFhoM2PXzK4VtKVmPYhQiG
n9amEERqiUPSDSa1eMeo/zj6LpouNQarEstDx5pqiLkQzJJThyYBAA0xV4YTI6u2
s/+rsWpT0lyIzkM+iR2posghHn91fjuq34dTTEzM9+5Kf/EtcZSpIMM45H54hA0t
55gmGsZ5LQ5l/Sv+wsOkDQCdeb4kUIwvrwiK5wArEO4tfKj80kavWRJWHUV5X//u
qawQ22A9S6rhwnewB5kq/DinJyPGIU4rJ7P9f7voB69wx/Yot6T+ZBH33DCzgo0R
8WOpIupRjypYWKG90QtJSr8PhAwzhF4aJT00XUxjIzToGTb0rOO3ujUukAxNWud/
M6binUMp+JtWLh8nIGNVlZzuLAFrJMsYtPoHeaCSGYnxQ7YCx6apqWsnRj+2bt1z
gsNtkzn/+uWK3qiHy+vH7DadE/8BQyStEzd42z3Js5Y/XVXoN8lX+zWVeNNoRm4+
g7UFTtmmRK33f0PNl+zdHfo9bEI+3CfopjxUMG+s9+uTlunExKDAr1DDBF2AKcDx
wfvJJTYdx1V4GhjfALfno7jqq3nKXP0AaCrO9QQBSKSaM5qiDzwfcCL8Z6L+efGv
57T43LrSdGT98MIby44GRZfp8e6ZPo4AuSAj2+dPQ/Q3TyCQm8Dd0ilZRWSNAe6J
R3r7p3bufTBO8h4X96wQXjmMkfg7PkAjkIvfLkg5dVGBM5XOADICDq5VyAxiUA7O
JCkgN9toUe30YQ7FHpLQH6zfyvGvtyGTkDZUO8Y3pQtMPVBHVhfjw2Fu1G+Is8B1
Aza1u03Aok63OWpWZMrhgJy8z1Wb7bIN6/FP410kY8cWrI9ccutFABxTD7gRv226
HLzPM4AHlk2YH1ahJbxmyZEVanEZBv5PCY8/Ec2pZWy4Y1wetuzC4S0faFySLiYN
BDTxdEJhBdaFVs0F8Bhod9NO5HDMHSvNb8B7VQyc6JHp31imxpt4oR3ntzAVJ5SR
f4CNKeJzF92YdkvawWIP1hK/nkQuBDWqv+5vvQFLC+KzcKdY5YZZSmTeDCHU+bPT
BPl1Z6lmyAGTRGsUWvq+R+J/egv+J2PfmuJO78m0p/2gjZtYZiKpusrm/h0rJbrr
aArA2KaIQMHGCwoieODN6v98SuuVRoh3ao7yPgl2mSedVtADBqYKXWLqmTnCuDe1
mfw9AnX8k9YMSdAPzBWo2BoLLkfgCU/QhSh5R4WBrMSIiRxrr/1voRablP2vGZFc
ayVs8iRX+BLHcPo+gSwSf3RL7DXbZZexss8afUmUlXoeKufQLkD7owfrF6nFDQdT
ZzdmjlIV6nHVuVwU7MT0fStwaaDD9ko/9hBnT2k6J8dObl5dEAlBBvNqtCkhJSAB
EOjeLcF0jO7nSXrAV7l/EpKq3jrtaalbh8RbuKCdkYqFWxWwAmEw99hx5fcQEJSA
PxG7UsDuVTP0v5tfOpNtubq9pT6ZXU5ACYYc/FhIghyf7phba9dKxyO5q1/n/iCh
V/TtX/0muKxe2q0RsEkGtqofiawZqCMLJNc5kkmSWbnWVF57nwhL+akPmT40EZ8S
R1+KS05CS+x4jCbxNSAG17nKCfd2Du2iOIG0rEZmbhBECb/zykmjYb32F/1FEFbz
8DF2Cek2cykZ8RCAweIFZVfpiBMFfDDW4WIocZNiQthASSKVVJp8rU6gl1XMWbnJ
jQdTmh1hEJLGW9MIfXvlMm0iEmdOQH+pAno7Gjo8UEKX4tSp0re6obZab91UGVVV
SFLkCaILgt3kUfdUv5ap0eGvJNpt1UoslQQuJvm48Y52+CosSJ6b4FK50moWhlLB
5Ij5Q8FaN52DPFDzktFRoNxq2h8lWnlwAUhByL6lJNKfSihijFeJ8bKuQH1LhnOY
sWdi6r+OUKIkZXMgTi3vEQZ+IWR3271iAnN7+slXM4oIeEBkz2GbMaTjpzVvuojh
prkbUdf0UUe+0iZE0bpTtkE31AKLy2p9XaQeMxQ0dQbSJ2Qfh3Umek4qlmOC6ITk
NyAud4qmmc/0pd/3IrOGdWfWanuEQrGUskcmZO0a1lR55SL/1qSu0uQdgdwvFCfr
4K2wSkujPzSSuC0ooWyarVH09AZzZSNs+DVQ4VdF68uKcp9Keq2GqAPkxzNJPHfv
DNyHXqNlQdZw7PuoxsLOCT/h/yfFmyv3xFR01Ujhi8dnotmXS2xVz+oIsLMUBLlr
UjdwA8+xkxSUtcMBqBOnvAiiFrqF4xDHPROk2BjWwNOmILBhU/JOcUmAiNJV0ONl
YqIewksIj1YOBLiKtKwpQYUAbqahEhiZHCIxwt0Pj+qhNq9m5pWFFyUuiOK86q0t
JkiHbEChBUAKFyvXCKj1nA==
`protect END_PROTECTED
