`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8fHH8g6fxURmkjnSZIQhx7TagMokJ9XUULfU+mQwdTahqbOcc0CKngtUTEDCfeAe
4oKt2SeXCFR9T9CNoq4AQO5oWrhKLYcDep5ffbIe9CvO+l41eY5u9HuTgekgpJeJ
snKAdXSI3GC3U7J2pUe/Tv4zmHCSXMGVxAdczJmdON2D0V3JG1FrLMwWjSpBR4C4
wLuheI3RhKyz6BvaMqJz2v7uJxW0Jc6eURZfK1s7a5k3/tBXBWzaey5NbcY61IhV
mpDQS89qQ1+cUsGEb9EJN7dw9S8AFHq9Dzm+k1OahdSkW0PXRMlgdC+08hekK3Ti
an4gCT9PILrKHxmQqhhvmeb6dRgIeAG2ZFqupRG8n847QIWAD0GOgf2kOlKLsNu0
odaoOwANUxyql4r8ymORogq9E7lnHgN736+TpscRjwoXNAQChJjGLDD8TeZpiRdQ
vQRgxag/irXgusontKQIfc/KD+ztBylilDBXv90b75uxMZfnxaNZlelbSgwIqS5e
i2sxzOkOTqsbcb0jZEdpUxKzvzKIHnnSn4gVQNiXLLo4FyUks723boAsE3pyhl5l
Un6jF3UjChmr4S5tn3sI3C9n2YIFCTK4Bm/xxYv3L+Frcy0SbI9r1yH0BR4R3rkX
xFjbGdx0hGRQqkjFtRGiLvTvA+q2oMpqCgr3aBcrg3CGQLD0owuakuF3txNwVdG5
VF/dosnIbis479SbArTllZZDSdu3a8Aq2JsdHuPyiwPEKfq1vV/eT+2v+9w3xA9Z
aKBCUnOYzZpBxS66WEWDG1nkBv7F4BoMhYdtZCw/YcGCLNjk3iQqAGvxUFqGwbRc
pP0YN/qL8mJ/BIeLMsOAy7128INZUpA9xHEYztHBi1YwTQExz2lXSkVQ9jH8kyFC
WKqkNLddvCwWmw/zux4mzLuBoE3/hQO/qDCcLy03YkgMEqOv/UvEGYjY3Om6e+HN
ucFoDJWr5pDmvQ+q1DbQGu4xxRcJiTAkZxiayxXvvYj51tEEWijiGA5XmeNk1+It
zBVv0VQPtcGN/f8HXKswGNZJ6U7Hdi7uDcj5OY53TZ98NAqfz1GtpZH0mdVYjH3A
nrbz3lvwRbWlZDsjG8RQFCdKF48awrCQzKoO3jR/leENdYula3DNm5Q72J1xCzrw
R30qfbapptQmE6K9MHK9OLu1DoB5tJVaIqAGeYJeO//Tsr6qX9TJ0YRMTZVDN2vF
Uh+heUAheFcax/wxJ1wuKhZN+YnkE+55kVT5LLuYFP6z31Ij/Jj0ueWda1/yNGYw
WP+2rnQjPXpRopvlpPwEB4ss2nRI92yB9dVZVkdTuh6QCMgJg80GajAAKXSDiTih
rvAvjko/yLHoeHjlrztZcxzqyJUc+dvP0WbKohqIO9MdnYi5j30H7G5BPX4+HYVm
PgpxJMXi+vux5YdWATnpvDtzKFp3eagY/nB46jCVyoDTc7oTO29fuY2BHjc7t4fG
X5VqcqNad4Apg3um2GPFHVUQxAnAOfmvG5KYi5YMYW51lsNIZTQjlmGSYy7M7ehH
8OJN+wx/23wjT0x1W7SXCQWqhKpbIK4bX5Og6vIxxRrOvhJTe7NhON7y0ebPkep2
RJKWCuX37eKFAQhSrrnEjpotM/RyltMHQJ9f8dK1q2bTvZkUHYwiZJAvG/ztd2yN
Ut2xQPj293/fY2m/MxFqMVh2M6Ji50Bn3SrtbMQRlHofZgfOT5GTPeb+xtN2I9js
/bcl0vBiy8eazP1KGO5ZL//VofzvaPSb/B836TLti0YZiFhNGH2apWekzkhYSzRc
SL/t/gKmSCaINIEOh5HFutuapnFf97aO2X2JNlYhivIaou8wln4UTfBENfeuNTSB
oxdxPnp091FA0ZD/Bef6kvNab/wNi8aCiqceiAg983npocOY4IZ8y0bgH6g9R2tL
VvoW8Q89lBS5k0imAIBWGm3fdQPTcltxLtwz++B3qYL3eE7F+UeX0Umpg/30Lz6t
PJUL3zXzsGWCCqttOg2n+lY0yFrEABazb78pSbYKrzXtLTYCTRNIi41+VaS15UEK
6u/UIjDm9mrEbqiBFGyqmnUzihfBIGF4si9HTo40gMDqDO2rEqed/B6orfq/TUrJ
a+NB+7CIVRfouU+pRLRhrZ6TrSRNGPtwSGMJYegqPhTHMGS6ywttjq4moggFk6ML
Ija4KmJlwIZcul16ChwzNyxQ+9mqaXtSqi4jvbkLcTJ2gpbhdFQROozJakcBFVS3
I9MX5i3yAmNp9ZwARtI9lO+Glxl1yrvK4yFCZi2Wnn8NtvSebV3S7ILogIoBkEVo
2iCidrdc0+33rk1qM/Mh5/3Q4LPBUes4cP+ZBW8LjZawnuze55OhUzK92BFAnAf9
FzhKUOUuU/NCdQxURAc694iPT1F+MHmJ6TD2279MoQA5woSzs+u9fvA6DLm/TSFv
K3Y/72u/mRnocgZtZKNcYwimUTegWnS+zfgENFvFzYiO0n2azGUnS89eXlEeRE+K
bL1obvwXRRBd2ZAbQFctIgIxj8LfzlLk6YQRfNN17ZmmH+dBLPR+iM+PejbUAJdl
aWs3U1pHaBIoAyY5weGYXCX1iNVUmXmrITNV5tUgXww=
`protect END_PROTECTED
