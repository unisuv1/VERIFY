`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
f09dOxSpnPUnDKCGCUnYnfTJc0UI2ROQ1gzBP8M0epsbyYrg/OtM3UODUX0INooe
CGkLoZj6iQZ48GDgLF1RynowupyfqZzwBGYTv+wnooLp6AgX4K8F/NKC4xm1tisY
Oz2XSnstg3OhS0v/TMRSrUvXC7xCXMZEThGSVZSPgbtn+Sdjg+nJctR0ugxy9UiZ
3xWPUQrXtX3PYaUdKkjgV25W9zhKA01GCCKK5mAaVL/QnmWMMbj/9iLBSOf2jnfm
j3qVnZH6Yo94BN/rO1GqCk1mf0uvfQxewQlLfd0GE+HYrSDqrWj+5KSt7Zh+iipN
McqU2oE60T4ixyjFhQSjmIPx0SRkXagvc6cY1TUYBK1OQYgd9OX+LpPCMzwQ/bLz
eRKdn7Smg37gIlkAdN8369eOSMJLXMq5GJoiVjavpItLGREUk+DLFQccWhP9yw5P
swez9M5RxA9NwD7HGFsFmYN4H8QvJrAr2++iLhP4/Ld8z9vDs/mgP3AvShqtLzZZ
2OJvR3CpPQstEVNhR8GwoKp4TOVO5VsTWWcWgGVuy7TOPpwia+qTUPeVmU11w919
JWRpkxRkp1ovDmbIdqEw8ZpdSa4lWJHVp8nVK2SrccZfKCy7hZrKCUsu15qw0Jo5
j0l23uUDZjBypLMB2c+MiyS2O0eN3FDWJLFwYEqT1FFmfbh4t90VO6XQrqvR2scL
aDq42IJoqcthyTLoAw2F8J3jG5SutsUv1+wT39l1nybZtxMRHkof6DxPMzq43GQm
w769vllQ4CkLc0w/W9qkPxfC0lsQwJIAhMSiDct1N7SS2MBVh/Bev3WIYxvRaQBR
fdPVebjwgsi/BgsSLD6svP90vGMoRoacfCWTbU5NxsfHfk7Nd0+sDjLZC5XUUY02
iMNj+q1FRlloZnO8o2UO+Xvgpnmk8FRJ4XIJeNpAxbVlmg6Sz6XbQjZGrbiW4d8P
bGWZIBTIwgQuxtWSsH0LbvczTFRcf17E0Z78q9N9GgBwPR2u5dojE1J3SCAPKK2H
DNc+XZde/41nTKZL2k7viX55RGP2Qf+AVOTZMr9fJxZNfLmrrEqS94zaJfsNMLN9
cFML0HS9yAvRv0gGTxMVdqxFJnymIwIQ9/FLeTLrbTdDwRHMNkEgce3Xw0DqKsma
5XTavdMGm4o+rj3pUFBi7egfdVFX3qX+HlqvSoZsXlPlVFXeusJFgr3ymvCBOOXv
oBqhAzS5FYUXgwX8ibMwleeT+NoyHemOn+SSFZVrKx72D1+QsVic2AQgNFVPEx3L
z2L20D0M5Qk5nozke5QvGx+8+m26W7tCq9Uq+iSzdUopaU0BuUEaQJC5ahJpBogM
Aqz/licojAuc5+X8OBAcPyU1Y0UHEvZCljpZYsnSh1F8oi0fLt9p4GkTFsJy6wKs
OWzHQ3Nx3CIWYEMx/yKMTLJFqMWsmZP9gxgdmdzMdD0W4TWx8pqqC3DhRcUKk+Lf
CCo4u0fsNZEE1syQSx4BQd/zRsjAThO2+hECsH8u8UIaAkjAfiHrMdVEDsybb2ST
Z3aU8OP+/6bcLgaDWRH2fYrHiHWm+RzAtlT3KTptPIOMP0bFZl6YTM2/p1rm0OuJ
6X7LsNwV86A5tsCObqSCasYaitZYwUbt2uzPUGzBOt2w6W1V9Rb+T5oDMwmmsWI/
UYcRWpA6EZwdB3HpBuK+P0OIlgC9K4fhJiFbOM49DB7p/WSGsx98cW5NQo7fHnx3
zsek2q9VCPzLviBnLSK3OvQZr26FyBL5c4KzlcumFsKkZ+YaPONISoaqBmy4emuo
05NV+o83w469X3GhnyrmqGshwh0IoDTUcxJ0uwx9nN0A78M66SCHIUz9CHvwO6/b
hGN9m2XlhfIp8pAezLyQeTAyUS49X+WuRhjtNlisL2AEzxcspvXN3TrUEZK4jWCJ
cyv3/Cs3JCTv/l4sQ/2afVfpxC2r0Doer5CmiPAIGhZsLspy7uQBthujA9lPmOPZ
BcvXOQPGwGYdBOww9XJZi0YkmSsX0i5gOFtqMvY8pFzABIFKCozw9kTQUWT90QEQ
p9GHDLsLbSMYgnW1BVRhk8/S0nZFjDBYoQbSaI8qw3Hb6NsjNeJgSMuBWRVw72Ae
XOhQdXiQQhOY557QUcqF4+2eUbg65zKwozOfUT5payIB/Fxqjaj5uswjULYPGf29
wo18VU6o+12/v2d0Zu0N5Kgtr8XoLjjtwwCNAhQhr9A=
`protect END_PROTECTED
