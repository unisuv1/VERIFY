`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Kuwd3bNxkcdjCSgZwpDrKcFCV/duIrklR2b6dgwYZ/Kuf/rfLsJd4jIlSz5m5j7P
y25e7vql/QSECa32e6//FOtDgLVb2RZC6XWKNJOkFpL1hTTXhQY2OSe/6m97jY3c
QCKc/IjZaoGYQ1i/80YBqhKob4tnLAUacp0gmBWLJa1tfBhAf+FSqj01aAKj2xEC
lo0PXNT1TzocQaBW4pBIxNVPOZpQPRQ1cTtuQKmMjZlh62xTxeNhVXE1slej08HU
muCVlI41aaaDRRH7FWd6M9/m12a5JdBfm+gqBctJ6r9gtuLGAl0HDHbSesVWewus
QjNXPP/aGFk0ioUK6A5QsM2Nrb2DGA5aI50u+m9G1D++rldKes2LIj+yhvAS17k7
dqsqnV2pYtqFA2OKPyBYlCn9CL1W5XPs7N+CfToxICYo+Q8buAhtSE6AYEZkJeJ3
U1n0Iz2uP+HlRtZVoEVlwBJsWy855P/UqUuAWGlIb8B/nQfmcjQH3ZgX+XICGHoG
Qq16bnSz7bidLf8S4BGRqf4Hv/1rXNJNM0uAmrKCmVJgkkmT8zJIuP3uS14s8YBZ
AbLNFqNO+BdAtfPZ3uecv73CoSUtlSJ8oDhbVc7uDrIFlBPmt+0sRk1LyTs8tDVW
TAxiM4sc38nm0HrvGgzU3I/+alfaXnY7ZoU95/kBedVOJZ5lBRS5gMQdqvE9ZYMX
HGZrOWHOaob5MeAvY2LT/6Is4zOFtmw+IxPc7vlZ+QrPF39jsvmeisk11HdyYseJ
GsO0JyJUaKYyygDc0r0T7dbvvxI3ft/5aknWFh5eNGbrNvlCcbYhPr7ZiQP91FRK
5bD0BzeaMXoQLCq7+6m8R00V9J6sy2D0aswMlbuEIcYnv5qV/2LyK0aeZEZ9Cw5i
DIkVS6/m5XFO0+DndNIsU2TJ+wMgrNz1iLQNnpVu97oJpxkh726yA8vOS4L1HTFP
C897UKH7vYA19MmPAn80KObUg2+UDJPp/8AXHUHXC/XU7Ly+jd0YACAe0VXVxXqK
IG647eikFL+LJrplLWeGRWTp0tiW7sharThgrY6jFYdy+y5xXi4+slZez315msA1
faNkQRXsE5Tu7Czu9NiziUx5XywU7c2cUqwk5VbvxMrPV/wCIPHGmgLk7UnvhjkP
lucaWMtDETCAb3lWRHxU+2EY36pPgsL/LooBaOtqFkJk0na0uUJw0COVZS/j6IC+
VUvOrlPQKsK1JKihmUFIXH3b3Z+c8YZMkS6jSfkhZzpb14JoWr7v8TK0TxgyPIgE
BeGJJuHPaPaJu38eeqzLwEbycwIzZZaIAAOTIGI0qyajEesscQDsEQiZKbnBXGCz
M2n6bCSae9d8VEAk25u/sy/lrLINtz77sPC8SL7GLoquFZWVzI3ZARQAAKW4vXom
XdlJ5C/PcqL60luDF4hAWgfOo625TdqZgiF75DhBnyCS0fZe4TzYAmfyvSWFRpw3
hPJ83fIidoHcJuzJu4UKAU6LEwyrJc23qTTjAeAr7uE=
`protect END_PROTECTED
