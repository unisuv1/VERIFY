`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7k8ZO+OD3QTIu+J3x2jhqo/0V7O/meudOYVlRQFkX8mAMmlpA+SdG4ya78BKDt/W
szHsbnWJVAKkKc5TptvF3NR3zjLR7IitR7TR5tgLyY1MNlzTiHo5Xp00ruanf9RK
zgkuTOEmKAEZjTZQr0kwr4wysVt5jYPV1f1hK2F7rTdam3ECEH+b1lumMXRiWVUn
zqlX3TPk7DiY6pJaHy7f7ZqB4pPztQVCq6/XMzq3xljMKY/2CRrxkZ6KjVu1Erf7
/qT+eFaKlvPdmiFkymyrkcfjnXltAd5RcTAnPNWisrztfWJ3+jLh/n6amSBed116
QBFd6d+8SUBxm2ujE4iC3AbNHsOe3LfTu8iiluBANCVjRxNkr8Mon7JboXJe22c9
w2sheuK1AeRpbi0fxmCcAbb/B08/wvWVgRXcwOQW+01ZzC4dYMxIv7/if/qI6T67
WTryN8QDBknBqftfZNBKxYQkpR6o5gRXA2IiuUrYyHpvkPGF9AmqjX3m5EMIYvTV
dE1UY4tDd5K+RdZEIM3yc1OXiVGHjIkHUY0p2VkQDdWg1WYG7AGvBombZC8xjWRM
VrazOh+R+CGs7/iQzj1ao+YaYuE9EU1r8bnXkhTrNsShqbLca2QWpFRYF23gCd2Z
MCRClpl6YbvsoSROBVeCGjKQNB9JlPbMLiV+dU5Uvh/WN9MzQ35AnsaErA7g0OB2
qJS2pNOfiHONH3hdZrNoCMIC0U9s6FrADPZrI8ZZUDbBdELsO43ArzVV3QMHBbqn
EQOAYlvfp8yB9Vwqb7tAJTkQ1X4sdHhwIHQkz9aOMjUiQTArQlzSby1ULo3vIWx3
MhSwMaGOSusra8aJJ5CavtPdUzRWoYmn5kjzGVYM6TTTo6yG6Pwdld4QUHpb6tcw
OiyW4HKt3iEqS32S9aEhATCkyC+gkqVxCRYzGR0+96Crc++sIwoZarrz+C1xYNFH
FMIFUpuaEHjlEHUmH5bIyG2U9ZfcpIaQu0Pt9WMxfJr8m80c9o3n0b5+6fU+0hC6
gjeJT7oalCC7rD4HDX4ltx9tjpFCxMG8hiaEGlHzzVeQa8fR/15MGDeTPcclJA5e
3vNHev8wtH6pS2g248LgtJVIIQy/EzFv7BiQiIrCF1ZShG8haV7mh/OWAXsRT9Ac
msiM0yvT6+idAJwS/LVsP4u+aS3G76BKRzJUa/CuxkCtvVG7z0Ike6G0WexTxbny
xiXPY5TIoKDNo6SkaQTMoF0h+Ofvark1TYZQ5/g2FidvnRQrLzAOPTRN5ENo+mf/
elcRPwIpMpyDQqo8hVFusxBjNR6SEty54q93IUMj2sNclabnnKXz4H4g00JJ0jEq
znu7MguVGFB/q2/nkCdb+P9sWnhe530Mo/XK9RAk0LHrvrrId+SIMf2jO6wXdhCE
2nmozTfxIj5DA77xRwsfsMYTqvszON7sfTaiQh+Q2t8tWNa/32d6K6S3XQT6JErr
Vy4ZwXw7tBDwQS0baXZwdw/SC/NlxRuhvHqo6TBkB0fdnJDsV5pbdEfxWxwxbYOK
YXjdrkv59t2rtbTgmyVwNsHuVkmhJPooIO4Ia3FdZw+1cIFI2zQCKeziNfsaeccw
hUZ5ykWATC7MClTlrDydzf+IKMwSdhPGxM7/FNZjp0zax+fQ8PvzcA6Z3yTbnfXv
ijSnLFmaKpox4rsJGsOJkAMTAzMK7HrwYWLB7S75SQIiPhOp56MDCdfQHz0LIaN1
xUPJMM7WHpet4bglIl/+3qnj2rIx4a5sjK+zhrrpEjcnONwD8mKX4E86W9TZ+RiP
8JN/ADo2w/CEzcFt3xGLwtZPGAuKoZDVyWRzQ4TNDYmJACTrs3OgdxfGMKMblHOb
0Zw9e7MlFqoAnQytB0cX037Bgvvi5svo7yL1ikOpMbmRBWWUnyU6vsvhJ7HAyWVy
nXfFoz4zsxZddnGMorOGKxSY6WZp/cE5VJv7yHsngb9FnfvZxJMFomjkK0XefUND
AVvBt3dauE9avxzpQvdFpPMCeqUOlRQOaCpOSqPS0EzrNKQ3nL38R3qryUstSE79
pHKu6B82QPS1q56EmrZUeCBKaDHi2tYPzxK/rJVfWPXi0PPVdoRYtFcWtMhF2yE0
2n63vVR4HXsPJ0hQdgbHKXJpfuqR66PQ80Ozfvi/vThe2pzL3bLMgyJNUpzbeQu3
szOkSdpYuKDaPE/UBE87Pn6v1j24AxCd7vb+iQkIeZkMbGg/VsT9vJELP8HXR1Mb
RFoy0beCZfVou3QIXEsAl9+1PCce5D2VTo5Lu2wSIuAPablX3ZSzTofYU8LT9llJ
CI6Um059QVRpZd6wZEck8AIR7TJD4krh/ofmFWko3Z8qG4cRjpKnUQhkESL994qj
urvRaldmRlTAtWyGsjC8I04065jbo8H/vZMyQD9UXjACdR114tsoZcKNixBbziC3
vHEm3WIMmWXHvDe019U1kt1/hsFDmTMva0J6TRhARS0aBqlF+uQ7IF1RuRXCcPto
yGLCRKJTN/PCiCDpIGkrYnEp79GT/vjWNIAncIL3dZpxsNIqmwzEjfbUKZJsyO1X
XfP7NH4POlfK2IW2JtFhLVdyP6kvkKOrat3VsSdDeoUaTmvyXxH0vYhHb3Cr7FaG
AYHdCgi4xUq4NMISzs3QCnU3Ah9u7JLfhFbbQ6ZfDumg8DRgMkE2dxQxWg8QWxyM
6mVgeRFN1zGVTPW7cqRsA3yswL2O/ENsIzUXDSRoctCSe6olJPdB5lSXBIjeCn2F
G7Lbbx2o/QioioKMaABemPQJ+uk4WM/WppuBQ8nul8uJU6pXYLbg1geIVAIKWXC6
YRYM9G1yJ+7VL+8MXjmFgkl6AUGJq56Z7x9DWM8LoJSBy/TBYP1nErJvCC9NJYXX
7rPbbXYo7oKN0y+WKRxKSuZET0spCoCRbQdepcgK7lYwmv6Ig145Epaq2lejWX9W
qpaHaZtNShwm2ILDoqDZXjP4LjpxFXIc6JWDty0Z3IFtGlgXQWi46A/vRx/lX0om
N++a468AHMHszYkdbsRMKwhAKtMpLBiQAs4eC10X8G3h0yv5qy9P1bkFZ//wRYeR
3fJeUcUd8zeMLSFCoGfoaWCPQbAhzfKrppE1/6KLyNwHwpjVYhx8K/cbFz/FuXWW
GepnFs0CeIv0TlpFbRDKBn6+DX7Rh6+dJXyTon+16L5luc8RZpovW2qD390R7l0Q
ER757HZzwUBJkfbUs14ji0InUODjRGjWNNacTaq3nma0rhcICtJOvEY1YbwnYFKA
gn6ogzvAdd7VQOXSLaYO2BofGNIlqhJ1cdYEW+51MIYLpcVT+6vFkLk5c1/6JNcs
+2xyOfFEKyD6atLyg1lbqUB3APWeJj/hKilkKr0wjsPaE43EEiJ1E6gw/LUh3QAP
uwT9tMmPnJsy6jjOf+91AUtWLW47uvXaxRiLD7SDiP2+eEQM5/RhrRHCrJ0oklGK
+HKZ4gVzRSEwntlguJauSQZ5y1UAi+c8t6jid0TXv49AwCG+C4zq+5YgpJ5U6lfb
sPjxmdoPE3+uYLzJZpJ5iMXn4vRtB3tFtmtnUd1YhiIdfrmJQF6Z9h4OioJB81lZ
ZMHNBNegYsL6dddXztxI97+0L6zOyTneLB8lx64HjLbbeirAiY6lQwZrCPDZAakZ
K+4FIDiBd89JYuRc9qPRxEBAND/SlSbuY01GHjKXIok5ICqUfO8KFh8L3glUTI+D
eAvECf7pyLl91wV1NxihsD/JwP7aoFUM/e/3u8rVOeI5PTt1nUYQEHpTCMJ0oc4z
zBo0SDJlKkQE75qzyzi6qIUwNcV0+3QYUVLDGGUH2yD33fliSyLAJ/0Ejhl7Zpsw
a4m4n6IVNK5gpvL26QBeVv+9STT2sAnKZz/6WNXu8NvYMID32VGlACkPAVZ5ee12
lRrPoPIEcz2znceHMFdMh0+4t3QE+IT0sNEzHF0SkOgiQEQ1+clAsg2Eyj6Kp2yD
JUIDSjsqDbeO1aKb1ODrlyTcxM84YzLHbUlBG0jnOUdOACBzTqUx5601uZqch0dm
OANvtK0ypfNMWleYyRd85TY3BrB7oo0ygNtwnWSSmma4//H7syafA21sKkbFfYx3
8PFMC44FnoY+NoKaLfZc41gB3cJxQwht4DppG/Pc6A/YDKyR2/Mjyw5I0nfewGQz
pmeO0alZTApLQWCen13+uyH7B8jvvRoJSHzoaIuSJTymAFIluA4qpOd4vB20BiBG
0MBZj8h2FO+D1Lv0VEarm0LgT4RCNrFriiq5wNh61ec2Ak+o7FlJASzAm1VakZRx
R9x/Hi7e3iz8r+eVIdmWHmOjQLrWC4GgA2sbw9GsdS2o47LCaUG9ss50YGT9/zCE
igwoPcXO7H7+ML2daFRprVZIDA2a2H945BdoGXrNNtAc2i346opPOFKHC6oYbsJY
xkcX2izvGan5KYv2FIs2rPyEWrOr7uJVLaZxUPLLkElPmSZKXDYy0UPu6TxoAUKO
Jf8iV0vdAZ6bDwkHdoh1oxusorLX2WXFDXpva4zgAjRoeYQ5CsU27Sv2W5vWWt3Q
Ku/p9cT/VPnUuF9gUvP5tQr5i95SDQa4WG99ZFdoYRs53ci9wyVZw9CmyOeqsBSe
MfUOaWTZvHhD//HDQB0v44Qx+8iTNw3FAERTy8T3zGlZOuMP6DTwFzM1Vf4CrH58
Clvy6WrKzGDC4Dpfrmme3OfNFp/UdAAlPhCHXFBxiqgPhGOtyGUsut2B4yCwDRe9
e+DMkOvwlFQ0mY5F+/H5yNcsrxVhUPUn6EwMqEl6+EtKjbn9LZGdZz2EEUiFo5JG
oRxPzIWd1usCVKVODL7FGFXwF++/DM5jhr6ZuNXlxo0pmi9l+UFd6zzv8urv6VC0
FugfBQQEF/InjxtwcCmzF67DM4C70yXkSdc0Zz9bQAC6lf9j+gtkwuX8h8R2XfQ2
o2K6bYKuveiCEf9qbPcif0Bfq55hIc7tt1vSupa/7hc8pKRO0PH6T74+dLpMej5b
yuqeSxoDdO7JiPjA2XhqZjePMeGcBHzFQt7OmQEI/+7zqu/wEetzEmtgnssm5hLi
Z7fb2Ws6f4kB5YvR88B4znS7qHtyzYmfHlEbk1awGzDx8fsAL3RbmVVSWz/wd2Pk
p0kFVwPLxh/90kmrZ9nPehDbkBYtklcVWlDuG9/eExTU7ZyYaWIxWQSW6Sy7rQuv
ENHN22YAJreAcxU9Nxj706Hc09Qu9cYqjIAMCfC9pW96el2rdIspM5sK2Ko5pgOQ
5GaGW7dxvjsHHg3pjdlOsPqja32Bx5SqpeFDSxlx4QlAWc6vysF+Im17kCvpnZDb
tqWIoqgaJUlt/HMOhXRtceLRty6Q1jwmzs/vlfr6Qs6UvRECUvzlzD4T5orvCq6a
jlbM/zr5+zhVhjuCf3S40COBk/9XnH0qJUen504h8dcUGRBts/rTN/2kYRZmU97X
NQVuucUCtLwgOjvcd8s9sJhP6nHLms64Gid79LP6frR7s/OUCn5m95PAlL6ESKtD
r3mcpmSvzfq9frLo00PR+P2NzVKyCu3aBHcw4GS1HNo2YBt6z4sCWojx0d7N7AUP
RbxIcrdwfpCso6aAqY50blwXR+1esCli/L6qBZw6I4l1fEBWaP60OtWhJVpYYUGt
9jnyVyxxIMjtPuf4bVFROCChceqxyW2gMET5HVushb5SdE+FZwmxFgBJkDiKpsWE
HHhxloTKcxsd1alxl6rMqbzd5G8GbdvMHCCZ1aAxnOaDzoic4UWm5axoB/5OW9QX
9MqzEnYHzg/mz8g6MD9n51COmrk+/E4+mMMLMZvgh/vpFRacEyDIzbBonosflR7t
27qHUsUGDFWUoOyWKkq9cbEbpbcI0Gt4Bltie/rv7aqrsl/qDp1rwibtTnMgr5qp
P7mucM6IGdxumX8+oIsB3EMG2qU7Yv1M6DDXVZ2WfjANHrXt44yh3M2tKEBf9d1y
VS4Xz54VoKBAPXUa2zI5ix4Gk1DYWPrLx9IGrMcO3uY0XHejNA15FNi39dwF148O
MQ4tkBBArzOPVZCGhA6mOErJjoilkg8/SSRmGcywzOtcyl6zKHH/1p56tC47Zdr5
OvStm2isTZr77f+fNdEeB5Px1P0kBjQrQ0v/F2N0JfCD9PM2HkSS46174P/+cZwJ
XJ0XGOJ/h0M61HLhQCz63saI1ZrXrybPwwkZVCLVpEFP6CPY45zIOtdKtoaEFrcL
4GIZL7Mymo7f3CVnWR0yhcWmMsjTHtiCryx1C4rOGLQ2aRttgJEaVQWB0bxahlJi
r1lueqDTd0jE1uUpITfq/WliEEsNjr6nsoRtkEHjzZ4TGNdNJqYfXhpLlgnD30cj
L1npND4Z+gHNgyP/iCALE4yjPMTmgjcP2fw6jjXy56sPNdwlXedIGYk6VthLDzPN
SmJdi7WlEe1fCCPygWEyE87Ji4oLK95iZ3YQFh6FBlPLMUJda0z8rvg8P3nybZiu
aUXuI61mDdgtrAIfG+bJDrSv+6uX0h8pAvaAMNRZszLluQ8Z+2fnQZWNbmpoODBY
C7venol3zc/VDfVvMqUzRXclIo3811h72cKHLHuE9HbGyO1MsleIBTtXW7MGndWa
VAjtlP3wdbzpCF2oBmmbcWzz3jnW/CdPyqx4M7DFwvUUaMlH8HP52P6BtmgKnnK5
4c5Ug2/C2oA7SOC1HfaE95L6T78ogZkdSGvPShu9Emjf7tsl70xV6O7ZhHHqokQj
bQQvAHfMchtVMZzFtD9elet3SmlDgx5HPeFrX+NRUDLM0+4VYvzeel948++3piBd
a7C/6xfrfMrNj3VOOzF0Eg+ysatiNj9d7iVBwWg59vAUtxdiI4H5pMREf6XWRGdV
hbIvnhyHuJbX7AfFXpiKtMA+mAh2OG6a9T/bMdpjogFFqhO+RjIPPF5ILzPcF4/o
32EHUk8AYYscXeUo9F7JqH46WK/QNkJJ8BtZNvKrpe0HF0Y8cd/ISJTfhFT/TvV4
A8qm2mGisvEiX+HihgI9WsegwjjnuGDgwFnbyOlxKsd9Hqkkn43DBalVq0tqdza/
5CkeTcnW8zMEaWapJ6jXpoxAlX2vhsxZIwi1xzdk7BuEWSzMOhrqfc4e2Xg4Z51G
F7oqB61Y9eZiPvFFsZ7gQjhf9GEweK4gexGP5mdNa0GCbnyCsnKc/TlN2Ah6AYwa
AKthhRXUbsS9Q42/+m85+fR2JOu5fKqGMHFYX5NYgq+Q+aVY8xkLCcPfYyEKB5dg
n+usB41GYDPXd98Xnu2+LpC0RDnb4JgE+PibYudiU573KJYzkl64BHW5hQoebx5q
Vu0HVwyX6xsaBJ3qJfP84fOF3B9BSERBKzjKIQCWLWCbbGTuJACn5MZI9IXQnQWj
9T+WEEUb+K6CpG29ya4QBGUyMLkdSWRCrHnR124uKBWqhv0XA7nH++vx/VWwaiZo
OJ/auWv7dZDqoP4GZvhyPyWqRKZiNdqGFFBMd0ML6KoSW5hbFXIPTbe3OFa3DIME
KDXTJnNIHYS9DzyPTaHYWtcSXCvGkZIE+eu08gEzjoTMrf5mYn/EFzre+Z/32jwS
qygbsjeUibI7OgGZL+2Z9cd1uxnRLDkBF2dKqFLHCnwppWvHSa2IBlOgC2CSZ4CZ
Bu7h5243NiROET8Qn0H0v8YjKaYJEJR+8mfRWpQLUqzn7/2+N8MyMrLAnCnTFd91
3JpkAny0n5+6HAgIklYgn9BxTxMsVxkqGUA+iNQH6Z/On3OEPIsxpPWUaVS7dWJQ
bZZ6GBn2refLAdQNwQw3KfVmbF+0QRHrddyFLz9LjIxqf9Wp/Z8KQjDZ68qeDAvI
QAFvUu55c7u3lLwfr7gWlXMJZ5wA336oCjWvrDDxuNVeoj3VCs/iitbYv9M4lIbi
NajPyf8Dxl/Kcnc3E+yHRmM+rC2lGSMXfrFeQ1Iqef1dMv4gHF67WXUMphcm8QTM
riT3wt5ZAW5M7pmqq6wp4Al29dgG65xCJTv5PgOwRaHMCNXNUM1aVgQ3jYtY4EaC
hfC8a490LIdmtb1rCpZnuYCuKuM1ikoAjFmrsFMyKbUFfA5Ko1OcA+zLEc0wJtVq
QSO2fM699oNs4w9uTT4yEHzdJlpPB4ADyZV528trDP5HOYwFsM8p4JROVHjYv4c9
gRIPkEYjk7D5qTg1OArXUKwRUDITgB2QP7+LlzOo5zQMcHF/n9ux2T7bXKEg9/fw
VGi/YTC7w+AcuGieZ2Zo8AIQDsZtw48R8s8MAvOqcYrp/JYOr4N95vok5KgVjj04
TbVcwtYiZGl8xYigR0jTk+9BS4wJbaOqm9OJ0ImXgVqCuVj9ePm/zkb+dY0JI1Ec
xhFXaGlyRTMEOuMfC5jKVnSjbl3CQdPMLmkvMM7LYiCDzoy0l363pXfWv8o/Ptpg
JTIDjX10CHRWu2F1Gb5Cy4TY6BVTAKJYSIdAnllP0u7wyO9ODAJbdWOPOdOX9hEw
LXemizhhLXzfMC2UCib5BL9+7Lv9ZxhPYXeMSyoGgastlkoz85V39T7OkuwyhEXw
p+kQRUEL94zGDxNo4V2zYp30RKdpEjAb1V5FbFiejEBSqR3XtMgSn5wH4/qx3ecU
TdgSo4rfluBZEXjAFiu/hhxnttEgROdo0taUMtkfjCxRlcx9RMbphtbbZhYg5D09
PFzZh69U9pEnIdWII7WaANTyy+XgwNqfoeYer3E9BXg1xGR3/afGo9rmBlHE71C5
TWJfXhoucdvfC8CaUr2k4pKOsXV773ZXZm4vuiJ+ck/j5FoeXcadML79EUMeb4rQ
cxt2K6JWWA13v3D9rmY5ZTmfKJ1VtetkHxAvKB9KhHQSUHJi+K7StZDqUeLHjtaM
C4b7IUaE6MmCaNUofXIJKxN22rjAMVZOvqrU/CapKzVTcfikY/Kdevwsbe4gyt9g
B4nZvP7FcjANxxxmFw26I/og8ZhbJoYG+Kq6t0WwUdjPS8T3yJXA+toUVwCEx9q6
nX4SHUmOaKt4MVcLhACxJ2Oy936u7RK43zTEgRjmKefGcKDsjDIOSkMLINhrxsKk
5D3TiWrj1NjtAMGfgRpm2yq+HXC/QET1F5MvQtFC+j+ZCxm/CNyzugzi6pQ5K2C2
WhxiLp9kwGLhZ+FfLrWGYLz29kPOhagcPC+QqMOyZmtcz0Ji9X2iGvv061XzXj1T
qtjxB+HjnbEEazWSccmj9sQioOoaeLyATe0tqvuHTkqIfySt5hFoBhtpLAV9kItg
7jtIbia6sLJICIhE4ZJiO7RTAN1bdMfnbpjPEKDk8sZya6VVrQzOFYCkqwwEtkAt
m4iYFM/e0VAZ5ybMm2EnLWs4KiH+Fo9gZBxYtGyjSA0SVCb1wgivFRpMJnbSBbl1
QC+cKlnuDYGklhO4Fv2Fcpy87BJALKehz6n45KdjGcegFEWUUf4iat2xhoRYjgfW
LWqGUWwXeWGF4erJIlyFRka4G6RzqP9FEtW1czRXl02fc24DX40pe+eGaZOKkL9u
10iZnxay0WLxCGBAz75+9vo+X73mc3z5PVU7XK31a65gbFk6ezBfFQbfwUFPij0h
WsIpf//CxZBr5Ung2nxmMmxBf98NQE2rLwqmjqTDqM68PdfFb2Auu0U8O1GxNmUa
sDAi1qsv/cbWlM2+s2DyxqV2uH/iQcV+EHXm8xcrYddZ+BR3UviVz1NPtITQObYO
hYeoQYVqUDpC5V6TVT1f7i5vaf1pm189c0O4r2vz99vq8/xC3rm4KKbQJfE7H2GK
CdffbZOqjzlPH8PO74sMkCK0rCQ+l8l0X4g8q6c+6fCJVaaCJ6vxxCvqRnHZ9VN1
ge5x6VYhzY+cciQjlwXqRsazzFu0tb4NN5Ytz8JrTc8jlIoFU61OHSRewJufSxMU
EMaHVcE0uFBVxulDGd0UvMDQVFkoye0NbY/6JvpHWiMRHka3vGacGle3djeAd7z4
4pSJRxDq2QXFE0blpSWafgG1/is70sH1BertiqpfKkiHjRy1NkTU2s4yRbUASjIG
5jCBTny9uxCQQmpSk8fTSMw4HI3C8uBYCFEu0fgDYdSk/Z1ZO8eeCLHwaT8zVZLc
zYpnQeSkIKkhX17lH0BCwvKbXT1DwztobBwU+npQfq5IAY+VMb1tdc4jKquD+zTj
gaYoneJPulp8eVAwxPuGiMAq7r+vq3pJpL9tTcjecEBX/fPbO5oL4A9zGBogzSo1
bRxAndD8+leIWLi2vSDKSZnZBBBXwW0ZD1SpMvYiMyvtg9Dj6ME9jnraG8xmIeQ0
IrjBFq9mXyWcNA9TG5hALa1siHjdgqCZUoaEkUtsB0SXTO3iH01vF9Wov+wNN1/N
naKeJzXxGaay1VLl2a0UWQrD4i1TzrVxGVRA7ICv4X1c5oBv6bGkIXyFK/zAdL7G
epkJtCi5MpaoTE+0Go8QigjLI748+e1P8C1DXnsgpr18eOd8qnELkwQePnFgSkT6
9XjpjQptRgc3Nic/rraEWrRIdEvB/CKHC6cwgCpCZJ8jdV3Xh5N/dfPPBuOpcvpa
HtqCCbp244ttSXGhVPL13FlaL7NGVjys1XiPc+91IaFQ9WN+7p9wC2LUNj41PpDG
J4VBWVm7PrwN1tmDG8H/9QdpRQgiuX+IjxlOB5w+57BxBKJ0q/9onvH+6OIroXEW
AdbBdl5yQq3jAaT4Wl+N35LyNFTS1okzR0T3MYFEore1m7HKyEfka42EVLLXeNOR
f2OJpD/Wj2rel2nkJfxThpFSDzhAtc7EGuEgKUYZKPT9i26gDn0+8uyNoBLha83z
8zwaCT9Sgw+H5148mK6xmOU1F94OgNijwGdWE0FNDBmuMyjpYWnKi1K9cg+OIhp9
lNgS6RXKdVcilxx2Ezz8z1KsZfSZSvqPwhrth+MUSfGy+p+DJ9AsR/MEAMcy10OM
C+kMQ7XgBa0PMltJnGTQQ526rnl7zhEkhvTt/H0fkIuwMY+5vUQFuqZOuqSb6oYy
KmACxpLE9GMfq7ZoCkWzJDYsF6fUdGdIzmreAqX6jRh0BVm/TmjjTNwP2p4zjsQh
B/CyIExgj5jsbaf6AOdMrW1wHptJeio1Tmgu8s+wbbl1hQFAXXMZql10LlkOc26p
52nud6p7m6xLhWbrdoPT/gc/DPqhtC5Cyd1NJT6pkk3XB9oGacODIKAbQ7IqiUIs
IUrDLa0k0G7lFZ8FfQqeVOpwVhPbT0UrqWBdwD8wN2npCqRD5/b7QkhSlyT7/tLV
itz/tLSNqIxndP8HqRnnYdEHouSzrVWC3BF9BVXrNncfj1MVRspGoLcGmKlQ/AFi
LZjKyLG8yiZa94WmvnUm71JQvOmYPZ5st3bXzuSUhdi0HC3FdnruyWIRro7XhA7K
bx/jHTy96CEAyplP2Az6i8/LwccDCT15NJe4w/A/bhf9b/OAvVXUXEBe2RHm5PMg
ScXYcVLyfIr+vapfvBf+7WbulVynUK1HQADxNtzEVarlqbJgb+oZEI/Sta2U7KwS
vpL1uhkKWHD61u0UIpsQ8CqkShha2JdfkbtzQUAqAfDFZoDbEx9WgBnZxAcBiQ5N
vL1KbHPhXXZ47Jdog2eH4nqOeVPD18t5X4lEQdaEdpQDnG+soiyt0u0Di3AlTQfn
u3f1+fncsQAxMeejtVJLciMggvHaR73v7Y9YNHOuvONUi17Rm2b+dFU8SnLLzLSi
v+zJLwpEkot41vicpX2YxVYYq2rpGKW8bRut5xSon2+66yV6U5EM8Z8YsD2jvy1n
NASS3WFr0s/fOdzFuaHZ/GTFoc496p/36slG/h9CnovacCmuc6mg9QpbAGO6LnoY
NNd8aGln/onLHCB6Qua6IMfMkKP7WqqvAunQIoanxV/Oz6n5c78D2uIBH7yqgJWj
PdDeqsDTsy5hhgc90PE1OW8nrAp00ziGQl/Lo7LkmOl4BrzEzS/wE1y9dRmnYPT7
i2BmrxEmtyV4QADsXffSdK+Z1HWKulMe9OGWOFUcmZ4WzX41PMoT0OplJ27w2qMQ
Y+cSQc0KWAVBiv7MNIF/+r4xaRtO/oYjDjeCHFGZQ1U5gb2BMv9rPwe28zBk9G6P
0u2rbXbCSXc2OJJiX8+R3aQ3qOPid9VWSXrecQOjZUl72UCE9YHetbg2Q/eI73Pe
Rn32pjyaWRv/+wUM+nZMvxsR4c2cuAPLHPoItu4B+AgYKnfP8AVfcABQskK4F7qD
1366+c4g4zE22TyFU9gXJSKEDg9AjUUrPtkd+ChOD0lDAn7a1VI9gOEe8IzP9x6G
ZbSiD4Kkso4+kA8ZGpcpk9+zNSJlX+AqHWsN+25dtGnNoZJMF8x3kfPwQcQJoQzT
sY5Ej1vICqMX+1bLdYnMC1VDaf8vM7jTvPm+eQhyC1Rc/63UJ5WqC3DOkmm9eXMB
4ET9/zezRm+D1zvf9eOl0RDql0fiMeoZXjKdyQPEXTY9nG4B2pYIn97vMgZaFe6R
CSXp4mmSc1P162TSQJAJsFJX7ormdNEGEAxRxB7Dw0qJgVXE0UD88W49Ku86YPml
WMpcEalfcIG9gzD7TIap6GaFvO/om+jKjuS93UAYx5Hq8J6vVNLlmL+aNS+m/Qww
OuJenn/gJNWCJTeG9q9KSiU2dejds+87sAo2b12FLRqmu1DSrvn0op3ujD6+MCEo
e99S9KJw4EmXGlk0eWuEz2AuJE0Lfk8HKbfYQBigsvRguvnmHEkce34o3MuB/KVd
Kag+AP0hGGE/38jMxX69lOrCq6LXeVe8xCQ0XCnvpuH+urScJBc8Ne6h6NRJ2vjd
JMud5J7DwDtVIg3KdPERjQKH3qXm29Bu+FWW3ujHZlqVP2bIcn0/9U0IlNQX9Yli
q+QBNMDfEaL5cCHHWDawc8iSUeQKxI03nJDC0u7DIUG6iUrUwLkFm99KBXN4NzYO
s68xuSJzmjRhRkfesYrRG1vq1TQ8oZmZNnZ336ZfKSay+/cPJIoC25fAI5o5SM/0
HyADqhuCQHUbcmhrfjelty/OgcpVV+x0EBpobK7rfFJZoMc7sJAtyInhZmK+xXJm
ATsOeR81Wy+Ls0zpZGQ0KagFHkZndDNoD5BMw6Wr5Szxhr6aaMbLH65BLPITJZ3I
eueCAqY9mCyW6efycK3Anrmr23XoAK220ymM0Ny2fWb4oIk0n3SXTKpGYssDxthr
BmsBHlJ1f0r3sPbEnb3CMyorFmpWTeFjELf/nBn1Yb/cRVVGalTW8I63o5Kq4N9m
iXgRsr9ytiIT9RKDbcl/jiuE4jhWvgVOKjI+jBUDBnwGctG9RDwCgmX3PSfmhG9R
NaXM6mqskENrbDgXtkMZT/+GhDbOeGFuupGv5WWIekcYW38+q5WUa1kYz8+EDHNi
YZpK7zpBPp6IeIgVS9vELHE3bUIdwP9b2DOMXaCV9k3I8jqy74tnYKCl2fGCT/9a
A9cB0ungWF2JXNmMF+c/r58QK3CXMV7ZT5HeFOuNBVhPDfLt55hV1vWWICsl3szs
mhsA40M3VzdWBVOu4f/t41BRSI4200hvo9oN3eyTyQtIoEnzM67PzAeQx3vSvpR/
PwTgJQrHw1l71L3Wsgi/HnySYoA5WOpZjdy8tN4qjNHZ0TAY02Agc2XBHZzrn9bR
NN4MHb1zDZJcVgQeq5bJqn5b10r0oZ9bp2ZS1405z7JBP9jpLtHth40aPgcSyLUT
iwkGa9jBCrmYLkq0VId5UjL/m30Mh1D4muGut74Ze1zTbNFO9uh2gmxGKkUqysV+
tjtYBLK28DxVLEsZWzGHMuA+PeEIeQzLMhr8PTq2THlxrPVTkmhTVyk05nDlNIxO
2NKq3sFNW6/rAKvv4n+UnjdeEJJV9n/ws2rkQhI6l3ibNjj2F3lIePyV61n8LhPd
D1cetOgHsIsqk6z7t92qlqaJvG6/k0RBibwQi50OiS/K+war4HxnXmAjvSx+bKmE
jdWSwS6znH2dleq4uNsR/4zflVfnm0rEzrggQbN57WDSg6N9xJ2lZit2hEAwiclh
tLxVTq65hxp9XFTSIGtzRuxsaab0gSayTPR8K2bIRjmeEjLduak7cPwoG40luvid
KWo7Q4FPWlQxe05GXHpcVuv3B+LAQcd6+OzXbMu7JKGKg8jshvbycOIXjyNJ0pIp
6ibfs19TX/bhG6Yz0VIV1CbT69hnUrJ7qXGnTk/MlOd+3te0aVghCmveyRtVpred
nyG8CU1z7Dnvs5W9yr3aANau1uRB8QWyNGQCuDlqkJ8s9SbKJPHGgEgTsdV/Uj0r
VDM4gdVnbblRrXBgZPHyXEjU+HmwOnzswKJ2hcIfhyN1DIF3PcFP8LP0tMeZ1FAO
DPNOiur3rukKnCe5/byrso9+cQjEEUuf5qky48mXuSmbgL0V6HhIaHdjy7JGRAYp
jjkQcGglYhGT6KzSN7PXWaCWLa83Po1P2xAtlAGP/PfoxC+KhCEICPyMGz33BE8O
Pf6DosIIeYK8e3vbLqyjvzS7duiYjQ2NaevY2RnWo37ki5vEGoPbnkhmXuCye5uS
jBf/yKHI+NMxwWn5bQ2/qhbMKvbru242Zx8i9vVkvro+KaF02zTwnOaR9Sn3kyf4
tGG/jwNoL0MfmKeEd3/tpb4XDXg4FV5OCMJU3QWIJLg5GrMPMpsKi02jzUO+MaXn
PokNAlt43IqGMgmYOG98fd1PioTJxCaHbwXaLYHNwCRChC+6ES5L59X/FFWw98vN
Ifrjy0CutcUKprTKqpwrhtYjV99abOzf447BXxPNNwHjsfxp7PxX4aAT05Hpt1tE
HcWhXnc82xJX2Al9FloOClpLMnLN0b30D3qdif1+uQCoVdnsm5zABjx+jJe0yuN8
S8C/e0Eo+WrEk/5WSeg5ScBesJ/YPgMXSjcsJV+BLDYLq8rbvcREHjnjhrFg2gOJ
u5FXhpU3xjP72fZ00Q65g1YJixA2AV03w9A5iREcuS6UaX3eJCf7jx61+/qp1fTZ
Wk6E5Mc9+giA65TTZzFHnwNxrPwEXXRFix7NC3gZj/5TrB+XXrMbFRq0ntbqsPkH
nV2WHbLpPZLZo9LBZS65XgExseH5rZU1NdwxwIsSUb8YmH6nXkU1fQSPb8Er+UOW
vSumxaCiqnCskof0IbHkfzcZyjGa4U+TEcadYgE+iGf3wGonxSkLcs9vm99jQybf
zYBMGktpLN78mDA1f+46u2iKP9MjPVHY7wqtfAJnQNlV7GC5Dx8ty0DStuh4PYdB
XQvMIkBdn8eBhOikzu0AuML8Kokc0CUuEVjpCYkhLejIjCXCiwvCIa9cpHl8EabJ
WBpQlddQNOy8qCvZxhZ7IIMiSllpS/g7t/JJSiKHekYKO/tcOqDAYymwgmIFRnIf
cEhSlrOx5q8tJGd2cDd7etO3slw+CjNIcsIqvlUL4B9O+FPeJ9DBxG7quxNN5/EK
YntX6T9uwBt2SHW63us6O4R65X/W1PlTgRYcEiZQ/amciloyKYbt3Ut/2l/bQ24W
xJfCUrHkFXhy/bnd7UXkDaiKag60K3E8/XVVxM/6pQfb5JOmZD0whwW6r6XAm703
3QXmyuMe69e+onteinzMz9iP6/DkdMcWazGNH2iLOD4bwnlqY0/A7AVDSMBraqXs
o5LKx/bFdj5vrolcVqAGRGYqea/wH8xPyMSJjqxU9dRB0DCgTUyN8tqKVj46lX48
Q4XyxtUEb4psp1ZMKb33SoKD4bfxr4K76VjvTpGEaCPl/KhGFCW4P5K7BN89WDBt
GoaMtxZsCoh1JkRtfmK47izGwow7MzY8dVBZVVVLymz14JpwhlL/oxk3j2kBXEMD
9pKPtnt4ncm0SvIToWAIAgTAe2w8ygkG1/sUmBZ4m1dgnXzYl50NxRlgdhtLg8a1
1XjUsd12s7tgam4zhKjqIxrK9OQzPECVJaE1sj4rNPa0Ibb/hAZDtm4k29jDNP4W
6CC0lPHIN7ElQzpdoXerZ7F44hZlYvrOcsSMnOfAMC9CO1raV9WpehM1hwcpm4Jf
5kVBZDpmrJ+Q4umFfyQ1ePjf58nySeW5ukOIE15YU9ZsAZFuY8WmTS+t1DzR6Ohw
UqCEuddg/Q/POq3TGWHJ/BImS0xdcUAaZ4F8soi7V+YfJfoOYUFAsYm9d6URu6fD
tUmo5TZY9vFD06ltADOSsW2183+8J6sZjzz7O3hLSVzZiTGQlB5XMAWkdOpkIhbH
xCRKMSIF/1ysA9wLE5Hey8tWlQnbhJOim6c3dp/moWxmAVHhdoyJoZoKQP9re6GJ
5FSdEj+lbZHZKLwoE3KyfsuqIWUmM0X5bXgTAtnfsNQQi5kTCs6h49m1cRZklAIT
VOcHtKpouR9u8+1Xpuk8LsA1tt/NZpPHvvi9GBwBirLbZeG8Y5c0KZ/XGC5F3QdK
hqYlQwPKnBJVsMWZCXCwmyKTvY8Dtmwv9pzwO50rZtCoeljKjuDBpqShouTgzasq
bY56fJeNrLjP0Zyuf4L1WP04sXhKB2aQe1w0crmG4VF5V0GWJBZYncWiVNrFYjJj
4Lauxbas56iR/7o1u1IcwZ71nS5OVamAfH19gpwgJ/kI8nQ5Sug85PemFApUn+Mf
oEG/6ntdXqbdtcBye2UW68y+oGnEHI7PYbUu7H2o06vDwyFaixZNxae5vj73LuaS
NaYM8/skvIwC5EMoP/4ZG13y2A4Y3bi6xJBVAuKMJZxml4V0ek81cFDEImRyQcRa
4vcDUlApZ6mw5Auj7P+Fx5Bc5cUgni/ElyXnYEKjGJeVJA3LCD4pSe1BdFnFFEGR
7+FLdwSibiRdmAAJFccKFML55Hi84AflHWmSUjO8hnl7eUsmuiKm0SOVL3b2SR1Z
0KqvIW/yhdqencBENf9dh3L8lEvGHm6dKHy5SKN5zShCxohJAy38sikCc4p1zBAC
OcB3veNuEVvSCKrdRacXIjXb5XFEftjQDGJamYRt9qEtH3wjqFHGgseGg9+dQNkI
2qGJ7jahWOBsyAb55jLOfE5OP3G3QbSCnJBe3FWHUgjae5el/BpoCFMuhiiJItDV
HNeeXPIH+8BFqtKoDdWVKQWUDyk5v7eTM9tIInjDJ3ZeWEVHqFi17nGGBS6m6N97
Z5G0XoMfqnOWBU9e9q+A4WytMeTTI7ufLl0P+JHaoK9d4fHguSFaspongIhneHDT
SdmPUQRq2d4ERF8mG5dpMWAsG01GHg2hFrZAnD4/8UbVnTwweA8PwO1ZdJN59moi
DMtHnELZ+GQmSkTjaE/jP5M6mByZWqtA9LshctRCY1Fc85qhC9Y9wRMtkyJlkN5j
OhlES6wB6S8EVXgadKev5D57YkdAuKoAWInOn+Wly1zJGZxkZUafXe40fKYEXAPP
UTxivOUri8R9T4r8Xv1lSdWfcLzN6IIEsCyCCxyNbWVJhMFDq7SCdvxfN8h0RuN7
7VaN8PCaKGhT9kH+WCGJ/qmGV4hRhA8fxdZaqJDKHrSpEo9wTbA6j00J17ZKiXdo
C5C63EurlmJ1quyHB5BLjY7A4atEMxdZxOTTeoW9HLyd3WMPJEXVIkyrlLSjtKyF
P5tXRLUE/Fv+xuf5WbNqYZLHXsfWsjpaaV6/O4Y7e1v4DY1R5jrq6F8rTqAFpQZy
9EG+YSQreAAGhNvgVCh4+9SQKDlMc0Y9SpOtu5SagQnqkDJie1ho+qHakUA29hI2
UEAPYrwkMYN4Ur+VMBhW/d+ucDosUScOmMhlZUyTXgalEBphsG435KJxV11zfN/0
eeiUgfpVLdrmbW9T3F+j4tfIYgGrvU+dTmRpwHW4nuODLN0aNpH6q/XKgTtr3H0Y
etbbEs7/fxzP7S6a5qKO62RerwrbG3rAb9i/BuPWQqmzIsuld5RfdqIKOEE4U0WZ
MdZkor9fCuxzGriPrXEtg7qk7I+7C9HuCZc6wKwLRe3srk1+hwOCxhT756bG5Aik
+SKNMtQyJxkWNr8lVJoNWMFQ5ASJvA2h53gUPJVmXZUJfDcX3MzvFpwM824La4/Q
jkUGwH/98bXfb+lTn+ce003Z3gQrLgFGDRUoIThRS9zUVQ3C6aVGjSm3C0FugD3x
eSLOdyPKS+S8fTJgJdVvsH8TBq04T+ocT23plsU3T2sXFNCR1bZI9aeZEMkjq+jy
wRus++mkZ9yyQgj3j6Peul4xLFQsKEa4E+/6d6/k+miPCFwK9f721l7VSRDFjaXb
55RpWP9swWK6NNyO8D+e0ngeZZEoC2uWuKK1UESl+IpwvrNeU3ty4qP8cDQAu/B0
Q/WZ8G4q67zfUY+5JuPTk4pPcqglNwxOiHbp/C4pBnzJG7Zmkgp5eU66ud8NXTYj
8b9da/Vw5biZ7UEgngAHNe40P9yXig8o9SWlPVO60Bv7EWkv0JbXUkzH/S3Z627v
Uj/UnQuam5ut2KsK747utsx26AmFvEhV3j/c0rLrnwh6xDnfmVCag5+gVAhW4VhQ
cxgYcKf7jPEAxsBElYlvDQDQhaClAOxuZSSYjdTKN7QOhqxPhNA5fAi6yeCWYBg2
OY/MRpeaK80fVgDucD7rJlg4ASIU2RVBamadn94oPuDGOQNbq0UgLdmiwYXBVQvo
d0V8ROYNVSpqR/TgqEVClEPr/lOTrMwhY6l6jfdR7ZN5h8jl6/J2/sZdy6TZr2pG
UTpkRbgaFF2xGCN3HvbbCmMO8gktPnMymbo7XWTK2XH3lkkxrGnw/GYCNI1DptU1
pSvaTvxRjvdz/XXO98w4jiFuPzrtcwPrNAueabMEekcAjTuCLeUnLWVK6d4fDlKE
te1DUJYjuHpwR8+Go6NVtdE3WuoRBqaRj8w+drxZ/TT3Ff3liMECBkUIb96bej0x
A1pt/LMNHf8ZSlZTIOw/E6B8cdXAUAPfUzBm/jLYQYSGVLRSvC2XYrD1DOghZUHs
QyFX8b5iSeiDvxGK/bPD68B2Dfdq+hHUz2GyGyIu2l8+6mQuU1G6b87josEhk3IW
v/RPWru12y3nuW0TU7u4aJIUfec6FqtGneQBNtEfcBsRkeyqDop2jfqYLiJpbhoZ
JEEgtjqM1FrKOJNPLIOK0OfK2DWuHUZjHk2MQvZCk3mkVt8PMuOT8mgeZSQaUD04
9f2eRf8WXs0QBE1iXUwiWiqO+RLnW2pDFfH5WeflmeAsaRNzHiaWuxM3Xj8ChHk9
FiSTfBUezfSAt8zjEBH88OgQfvl26P2s4UrNt2xaDfvQ5gU9PKn8wB3IVF16Fh4R
9VkBP037VcSGrCMKEyjL9NzvkTl5EmcZmH5Oi0rfdc7dFv3CksBDU3ODXTppxTLw
yg7eWx0aFsMyrMV/L0Y/yPMoCzVHAt629y0nP/r8vzfJ4xI0+KY0koigM9oGZre4
MjByo8xMURrGIOk1ciNqulEMImlJGVgo7EVfgPrz+/bqPjFy0/4nCQLvthRpWir2
CrIIzc2GotduLV8N1AzZp7UCn/8XrhDk7M6p2j+LQEsd/tE4/9ea++r0UeSFXvkZ
4IybuF6fFMco++1sKExpZMbNQCi+X9A27HSaRgrAlXz+FnzqpZ3umbrVUFtRSm9Q
S6ZRA1EUkcts4T76h04JBL2DPKFlJ5kxd89NQmjJSsW3wjjg84jWHtGNZJb7JvYo
7twkt8yCoxX9Zvr6v9J1ecaZQMgVZ1hTZHjtT9JL27aFhg6bOSGwdHrkWp8VpuBG
31nujzx/LL5L1RXiVnl5sfQx1J1TbhDr1pzs2X+jGxpGGsoVfGSB3+WMJjw5G+AV
Pg2uEvrocNhj6fyYcmWo/G4zYf1Rc0D6R8pGDi1Ms4EOK6Nz6p8srkSMR+rE7E+a
Y87XKSxla19XNZaeAkK0zhmRZrKe7Fj/smQqiaUfanWgsOo6KBxAM6G7U/7SsqGp
SCh71soFM38lLNcD2Urj15+i/fsHhbAvVJP3am4PGfRFrb3JN2flOALndOOhr0ET
fImfqQQFIk7Jo01TLBpJVQmviRHpuMRAkLsGO9JCV3en2VKJtMjTmiH9xUVicodX
04irwnH5VtKkGFcrAHU9Y5OPGoAh7EaLz4IneKiBfeMG8OX61IU28GB3amyYhg8O
KTwAB6ZmI4lSW9tPYriciEUm/8EnmhnG+ufb+ZKtGDYxCyB1aAbV66RxBjzjoHsw
IMwNaXR3XrmteSMAoKaOOOp0G/dSp077rbHgJyY2MFuSlRleaEuUYeKdsFqi3w3i
mVNRyelEIPqqftReZRKd8K042wthemksglL1Cl8tAncd81/LKn9DQowwXoUQz59o
o3SkZlZsvKj5ahlngJ5uI/M0mxowNWhRprXGLrdxQK/b1RYt+qBzK+57mbp679o1
NL1ZDgSRbx/tFHAl/nxACGFJERN/J0Kqq2tuPfHzMzhuiYHsHbwQSnL4ktCX+jRo
SZc8K+iPH1ORYgZcfr5CWJioNMfqWUz3oFLmg/E8ZOvQODiNudDpDtcJ0dMQCA6X
B0544w8Y2kmDKIdXsg5lGzHmB00Bch6/5POuix22pDA5j44ryqKwrgjAHKYIUdy2
rZ6TU8AKEGt2GVJsjzHjmFGJcShTrtLmamTTvp4UzSNKIzbEZYodFGmaSS0AI4OL
gnnzf6HEC93KfURpTqTIVTzFIM2qiYAHYkRBrLGUaJckfE2+REI29MaKbtFqWY09
mFE75goNANbQ//ad10eRKgtOmUAzirffHi6Shpz6ZK+RFFIinqCIVq9jRnzua9Qv
AfEMiNgEoXGAFrX9/TMNW9Iz/HMZWLRrjkyceu3YBrKLVB6LuPkys523UQWkRBcC
TBFsebf+gIVSvN7Q317rmGRrljoLrvMS8vpbdTmdobcA5M7lbaJc2+Kkd/8skaJv
UO4ypH8Tk6Kct0gMPU25ifjIeFmXY3SYaos2jblVA0ZRM4RVxU2VfiF9mvma3sJd
bZkv7OVj+YxJxm/cZHzKsxGg2b9WFUHRNbXuhGAN1Te05MqO5x4IHRcw3Ds6lpvJ
uh82f9IBVAFEE9d9wsLMb/b1k0Mts+I+PoXOdo9b58u6QKdkRWMkMt42R2Te/GTS
9ki7PYC+Lx2qxtyqGVPcPvAXZVYoa5o7xZe+cFvmEH7vUpacwU/et6D55h6yF2Ih
A89cFsb3EB3yr2NBshSvsBDmR5573hP6lNjdkr8MuObMNH4dOANdDqgSPPR7WKWp
vqx6gWlYbcstayVyvGtQ9AKFYgGSfU/dIayr8bG306RxX6fPaGHh68ZQ0X1BU/2X
vpgNcJNhb6cGvCAnE/0KAG7XVEu3joPuWoPSZs6eIMBhhMmLeCDd3u+sH3XXqtT9
a8rlZc9cBgYFdGuiYG9xRf8WV4uzHaUSxBoGHnyVNfO7T/JVqFAdbIxaeWr0I3QL
JX7F3m9nNzaQEj4bOsj+pSXpJxZogLR0eCT9UdKtZUnEIMsmHRvMOk2HvH4KPJJ2
x8n6uy1dwZfQ9XC5tPAAQSqj6yPDhTSoPXIJtcdXhBgBAEw0SCvdp/U2GF92XnXt
qqYMqsc9FRKCeM8Rc2NyriWi9NmuCpA/tffpIHVI4ynsBvYkzSgyzFKKtRd1Zo5y
ueeeB4IIfC41LQvXdbbxGI9zuHvRBDJTx2XKwsmk9dCJnbMLcnIygVah2OTgTAZw
HjuK0h6ezXy+a06sjlslpFomGwrafN9Bfa4JNNI64iC7VVilWVPJve9fFIbUp78N
ZY8h631/QpxNrB0CzAfALU8XjrxrNT0Mmq5YCL4rvuDh2Jpy7DqC1r7Hd47JUE+D
obY5zTP562KKol6T26+bYPaO1a67YEmZzTi+BkH3kBAqXb6oerHIhKYT2Km/w+dj
aLEg8p3GKkIed2+AeGiL4iSDMd0MIZnlUrb8Bi0XDsY4z3hhJJVgb6k5jCpy0yuR
7hE/gylloBL4Jg/Vm5mU+MDfY/q6wd60LDZkoK4J/SW16KUnf8FQksZM9oUh3Ro7
bN45SmvKVVH/yHKZ1eoaQOlw5YAOOfV3AtHHjKzWVxWlkBShh4n8uHaH3fZXXW9u
2/mTLYfw1fBrQH40rtho7Qv6gzSqIAojZKGibGVUI+kGW7Te/8rqCajl5PhPHrBf
koHnn6QHS748wEX+n7Cvkge9X8hfTyBdJm1dVpejdY3cd2NmFI2IXnIFRQCHLs1V
tZ5zvuMkso0yA1e1ryTm7qFwYWtkvhNf4wuDt9sid7++m6vOu2Y3bdwX639UQRHF
rGc2Gchjrm4RPpRB31JJ8ipuuz4BiaoBXmv/VhT1jq3aazQxxlKpF5bq3dQW78rY
QV0a4RSfDFfST2F1inLuMrFimkB4jEH/czVKClaqRZhRLQauxS3ldHBlzqNqNyXP
y42z6nDUplJ0Rfde4k/XtVEsxGrPThxm9hI8K+mGxMRUDOLfRBth9GygZ4GjtVXN
QK8IHcHZkCSff1E+odk/nzf6iXw959o3QzYfNPGjJuxOsx3cIofwckdx6CvIEWZF
KbUHNZIhMdDGU9QqE6fgQnZvOJlQLNLbjuxht5LfB/0yGWVjTUDdUO+dYX/JnC/H
i0xWKpPga1mw+Q/wnxZCq2uIdpUvGkF0Qj0846SgjVuCss3ZkX25oaEyJtBi8hCk
k/w9GMXvaQUGfEWB8Zppb9c5ZWfTjZGPHl4kWbp29Z4Zb9Zd3Tcj49bmmmR0Kv78
j/eTK7xIv4c9QkB/7SOA0j29GZJ07e+n3wyh0wsD2JH6A4n/RYwPcDdQaKKACFcH
/2Dx8WelTIaRgKPcVTGddDy/Q+jW7nHiaWU5DeNkEMlSSMgPe2rOz0YUq076Tv12
UisJCtcLlaFpdMLt3V6TiXDM4/NvnZ9EdWtPT0xaBHMl+FdDoBtDTsws+NZfeWPy
OAgys5tcyg2Jko5/kXfgJ8qssaEQjzfbB+XGfqDRvK/cdw95DTDY2lOuVHDdLoJx
mjApIlFd17nJHP/pUYkFJTJH/+ixV9QG3LCSzMKl8A7qwhcczaVjZ/slLNER6imt
DbA1Bcyw/vID5+vP0w5pRFH+t4zmhLEuLpjKnN23g4o88zvjD+r0L3rJyisDz3TQ
LH+iZc09iyXOvdRJK3++C8EpM8p/rmjYIW5/9DmORbWO2Clhg0zKjqSrdG1x05Ce
uyxPqAsh3KFn9r5TAvcvqVhronpYm9It1342hANy9E4tKfeQKuO5JMh6CMjZNwQX
iHmk99Hbsd4wFP7fEoW/frZBZ/8EZ/uvmS+g115OMG2h+3bd4PEXxOkHIw+jxWQX
DZMCeM2o149Hc/7iZqVyhdNpQ0TULs5TaOFvHuXBw0DEOPSwHiLi72D1it91s8dC
E88drpwiU7Ev3mqHSRBR/BCwjScUUx0bj7FPdytMZCR4HTkVtSOfdqUkMJwpdJCa
liTphpKpC82HGjCx7iUaCKexGn2uXE2SBOOPqNpUHyf4fKuZmzVTaQyX0Jmdso5o
ggqKQY53WpVlJ7+O8uWPGd+gyIF+ZRfjELjyOo1bsCeuwhrJZ5Gyno3yv/0izSwt
jKK+MVM/+v7fZ78TZbe0HL0/8+lo8maMycAGf7SpQFbHRBUuP1pQS37IU76R2fF3
FcMpe52u3jmuwzEPSWXMqHdX6TIIuIhLFYO3BBEfh3HHpFvF2MIwo4rJOEXeOng6
uzvxPmjNN7BZRHgl8lT8HFngCIlr5UF7B5IEKNKk26vVJ3lClWBuq4wcvkYIoxMM
WBjKEc0TAExs6JLtpx6toiQJ96mj9MANfg3DG05ihp8pRbji0XBtf2XPR1UMRMhR
P0c71wlzW7rmPQTfJarW8jQkdF94KYi5cljaR04eMSzub9EmyYClwSLo5RF++fi6
T3yuFJrMvRsUEBlN+NX6SrZE5HO1TVmKoJtnLj1oYoKuc31Y0uBCMyESB0KenYB6
PfwWRxAcyXmNRvUXhgfpCULcHjxGml6Z6677Cu09jXegvIHJxqT/xjxNK2RGNkHw
y4acoBIQb6Z0bHwxxqBwzagra7NR2PdHNKmteOT3d8bCjeMd23Rv531Sy77Q2O+/
5LrDbYXPMvb5ApWgqjVQk2+rlY6yVULnSIgYkmjGgaRkQZnBILM8xRN6RsBR0oWi
O8hESs/XqifoVQP0S2Y8L1qyOsLPB24W4DCLDIaQ5VlYhzhaPINxpvIoReQJdGD+
ipS9j2ZyLRT2qD+0dB1Y1D7NCoDIQ7tvh4scmCmrIc2Bzv/ybOHHkds+/Hc4PyHY
fqkRec3mLIzFLUQd1V+WJy5GlGQbdSc6hLSwYsnQrbDc//6mTT6B1k5dVfG43Spv
0DHrUfoIVjrWzxgP6WwRycSNU9nGLkfFxOGfjXvB0K4qtmfOS0ikfIFJqs2u/AGv
vXnY7kBWFHtOnHn6gZkXbqjhctgk4RBbuz1dzuaRODiadBf2JFW32saxGjFq7tB6
VSvqGgXBUA8HL+tZywidj7T6C00WHu/awnkXdhASQ8lzchdhZwgZVKFeHY5K1ztS
Tx7IEgve6MGmAjfTUfZOcH+XchLq5sBUtXYRyqchOiX736R3QZRLbiyWdiQFTx+Q
IOU/JD2RgY6dgriFYqyJHNg9J94rEFl1MYG4f5Yvra1zT497jwKwxiflcMaPEQp7
gihANVO+PK9+whBnBpLPZKdwHMBbmF5SVujMWa/gTKfOa/L1yTnA8zAs0P2ZtlC6
HVbDr1h7aZyReHD4+GPbXlG9oip3wAiB00flsmXJqmeMYQf8paKZph4GU/8k31Xp
yESjsU2SFjA3lxYAPlejz1QFPcqgjGlh0Jdf6NcaRbb5xr0Up4OAAue7GdXx0hWW
wAVjTPyVSH2he8pUK5fciAxl7kYMVkN4cIJkzc1F2BB01VcFg/SFvtqrJuUI26dH
CTmtwOHZk08obbvJX+9+qWYagcNLN+6MEGYbe97qwfKrianS2TlF//9F/Xbg51Kl
WXUDoJpts+6FH22C6+zkOBRF6HXEIUqnX4Wezv6Py3en640KBNo/FrODOaWKRVLi
g3DGnLmSX1vmhVFc6XWYaoKx59kUqEsWmk8hrNLC5D4DoPI3VYgkaEIWZxAFlixl
tV6SIXxsowJHZcwlM42evv0weL3KYY2mtiO63cKHNejmEen7sJ8kE6hfHMUJKiPQ
Og/+Vn0HNksVICCso8cPN46+XxoaUx2l9Uc3B46eIOA0bCuDv5Ax1S0uZ4FcUFIj
bbbOzSx8a9Q1Bsx4FVL1CjMsuEHTNWHBH1eWp6kAd+jOehK36yOBAmgdxwOTVo1T
mFMtyxIurgwkxEDejxzwOABcwTTJKxPFyb9maxvL7TOp/jc677+btM2xSa4qGEzr
9f8ENrFVLpLcrKBZvwwOqWBmwXZJiSHjkGXizCzbi/o7g1dWCWqTi/XyhgAvBFuU
ACxEThOGucJ5Ps07Tnx8/LlOJD/Iw0C2VJigNA6f8eK4+L1ak2OaOkMoTbS728JS
ve0A6NmXrg8ixn95yMbBWv456LizQ7rrU3dPH+5jhaz1LhYJnEQkfBdyzWyd0sXI
BiM1wSyAnbXisIhEIz8gRopqh80o1rW/kCqHrKQXt+yNGQ1JDfXBgSQQKiSi5mup
AcodoHLBmmZkS8AxiRb2+zdPuKaVFxYSZYq259klK86CoOeuzPyDFinMVbuGuN0a
6RDV6aNksKScLs+B1KS6q73dxpeqLLsddPRmAb1NH2MCxXentH8TIJArysM2a8Lc
ei8oh16ud2Le1VwemvhASvBmQdskXT2y6ismpr2y67ymI6nKEe+WxNcr/g7gTrlT
8xB4MuS8zTrG9qGnb3KRhZl/Z1WuPcT9V7fs8gvH8e488lpPNfZB3UQiTQxkGBh4
txlgLy1h4B4LioAqR5dV7b3isUf9trSP81XwnLGNEBg6jnSlHATmktMECkk0/rtV
fkcjXYY0jgbKeoA0cM0dzOzh+ge/VKcxfCl2rStPVNkRWh2s/Sgb5FON0juGJiQM
kPPpm2w8u+4wQrnWZt/Fy1SPLOfaaiiBnURk5jxdv6siBt/vMMpw8JAATGffEOLV
kF7I9ePlA5B7JCqo3P+MqSkNnMjnoEXYyJz9VitLkWRn+sYUR4XZ51b07KXN13g8
lkPDZBB+7ljJifq//xy4NhnOLeJ9HK+fw0i694C9bWaDIh34JIOgGno9WSeV4GND
IWJ2IsayPNgY4ap+qkMx8xwWm90Ytyy84JnvLrq3vyudwVwt7ljNvvwzBsWKvdfY
qQkAyRCaHAVPkYacSFFqTClUh+N5VCsh43XogEBFuKaxsx9rLSA6PpQNZ7UnDc/Z
vEh8ulw3gGp45IYnqryUeLI2c4tkjP/2A/zGGlz3Zy7zRpMbCfT5chVaqtTVLzUs
+n/GQKWBMCSDUDV6UBmznYF5DfoHpdTCt2Zr8xbqYt9wSMiLVYQ0c67LyUT8PTfk
tQ86wRwL5sbhdp9VgOaIoXhoz9HWQ3s4Xv+Byb1mM2tVLgaw7+0Kv55RU5jcAn/5
hl3Wey5kwpXcK7vx8BYYVa83arQku3pi9CdH/n3R1iL12FEI6F0wb5/YD4fmcul9
tHCxJIS67NJO2UUlw68YieEUnMRFYEJikq4Fru0l0UsEk6ZvLzw4d3taiEs69a1C
yWaNSSHoAAL5bIQtBx/yCJP4bitP6xZq9jB8u/qS6kf5+VU1Td0WM+HVSxkB2ip8
7ILmwgUDhb58e+p6eYpe5RkTap9nvjRPSrglgrLngFn5LtPfdd1YRCcdC4PtEjzZ
ZwkHXG4cs+siwjvxMEMMJWVLJdpgfG2w6fpwVoP8T6Dlu4cup0lRmI+1YkJzK0sl
L7lW9K267oVSLyBsTIeuHDjuYMeD4gBgtaA3LlhRVd7BluJMzuYMzDaPfvqi3tbD
2uDiaw4IxhFN0zmAB1f5p55NXQSgaWWQa9ZnBnE2KqIV73h1+H8QCjNJwk5e20ef
bDMVd+M432ze27kAJtKLCfsG7gu/hpZX1AYR3hDyFSeIscbj6qu/B1GpuOcDIKXY
dtqkhlUukeK5q/GS2UQreXghc5BdrsZh1vBXqx09JKjMvuRf6K13J8xF2k0FZfgr
cN6zbB0eGUvDgQecWgF+OC8jOpcDvkcMQuHheGl7La7m3AWxl8FoSNafYgVvDOEu
5Vt+EzV1duMlJvZVNJlt9TEllT4MUWAXosnBLB4Vsv4Bbl7kDLBDhBiXCmZM/6vW
v8GqyOxkgFiUDaa22F9eokT46PMTADZT/zC9cDF+kspmkya240xmIrAT0A3lmE1W
fyy43lO5BcQZ0Wdz9LVMdI0ar7lqTuNvboX80Hpu7nb/GbhLUdoCdsz+GdkGPZng
mnHz9EFuPlZxU8T72A59kBUDDgoCGrQObj54dm9+jEXY66iypbGsif+++Kc1vgND
UFQ2Qd4+IN7q1Br+0W97eqlP7qlNVQ7qvYiL5USvWUtgmQo9kwQ78d7wJve6XbVf
06QGgTFm3V2nIfDYURvMcPn9GLUXGa76MfKStUb1vFYrrEWpVeDI4SVbpLaAR+3G
qIjSqL5e6zd5WJAJ8kftqPgv2ulxHbnbE8H4UZDmYztttM83zK3AxE23ODoIxaj0
WNQOP629NIX7yB7hS5YqfV7CCuPFjtPa3EaodwS8TXcKznfMZcoM35AvKzUI0ceX
iX2lMvDzE0ngZB/miPtTrULkte4M7MhRY7Yr6EQ6C4zfKGUU6s8DSAMPHDIWL0TU
lsoL65Qph9Zr3hUDygp+jUXFzMXoEkvhsYm0XHVLNCB3dZeTaAbhUll+cb6u5nLj
ciUR5Oo02hZz1d+FqtHpfZ/Kkg4U1rdb+Wvivos/dRgRp3gQ9cysb8iaQ0oMmK8U
yN4yXJ0EtapHeOlM3r/Um4+UJBSOqe7P2hlftM7NyC9jC1JqOGXNRblzFQxt0iqG
7czruYdCpvv9wM8HfXjT+0dD504fdmGNpZrS9NC16N5ZCfpPwWThEUgULOab0dOV
XxCDsJQYx8FUSZDwnuWjGTmeql4Af5ZEZgyqhWBkhb98oB/pdNzOos25+oQTHkkQ
9dRPq5b8O6pRUKaiyQNW13i8BuGG+8vsv6t8qGkC9E/DjXxQPpsW/hNlONrLBoiZ
+qP6FIlQDUEoRgLL0NFBl95QLjYAXYtlCuR7kPoAtqxWkxIq9/JWhK4YSMYf2tiW
V0aI/u2TA4h7B3ZOtSdxbM5p1K5IsnM8BHlNkcdszUQZFPb2beuKrdlLh419+Nwe
1DsYyB5JnvnjQP5nRjxsUCYmr1ag7OZgRXifh7uyFlcLCwMD+21+kwsIU/ayc5th
Fwvkq+aHIxOr6TFzgD2SGmtg6iyRkpPbuQYc5uIWDjz08crNM6mqQdtHwqv2HtZG
vhitQ2t3A8rd0v/h1gGi3qwWccZDU3SogNNjZDVuDpHAero4JQhO63znt/QCJQdt
NbeAohmaz/HCJUnwEVWkp0YR1YGIM9eCXGvHK3+PJ8yQ3ixaDJ8FsjoUfD0WCxyd
9wMRmYqgJc1s7EBRmj3E14K1GdeloYX+k+FvD+aqtdnSJI4WdGSVE0PGcXvGKT6G
TBvTZ8Ct6FJiDQc9FIn7rV94NyKTK7brnZRgsxWgzfXQ6LsSQ2Ba+nbHul+vHiv7
vJzxdKIdqSXbYDw47y/5Avdn9S7SHLRnrlGuyEvEPliqczWWK2jYx1fXEuj74Mwa
S5T7Rw4BtaRumTjofxs5ZzfB5p+1n3kzRNjOwp/Hf0hSN8Gg0MySKREoHl4XXO2A
ApDThxsJJk+j6LEYSgkk/roH9sM0rDt1kIGslRomU7dPAyPS4ItpJBdfqhHHSJod
cUDKQLFqwoYa34K4k6wp6ApvnPKCQA1T5L1iTCtInMA6ge42HlzX8bI+dPGZ11k2
mYpVLcqNKK3katt6JvwUJ8vqMWiV1WHHKJfEbgxwMRE6qa5xdGtJh0P6jU7b1VUG
QODa4TCfPJnUyiDbLT9PZuvIZiqhFTkE/36SUUpiXnuBqkzh8DeBat9jQVxc3isi
UyOFVesJYlxdE/omz7OoZXS67ThMcdWzJIp8WCb+Nrx48llQfOosqfCHmJABI1RY
4mwhd/qpP0jnzXFSb9fii8D8tRTeO61LefwuHPhU+lPMce9EcPpv5E06mbnH8yEs
jhxQN7oQucoBkHqABFlny9gvSe9HXc1DtX0Udv8QxSTBcVUhNVUeJZ8uJfMhUCMX
FslcMr7jvOTNC1fkm8bQJrMIsGObywZR3NmmychpMHubHMjtP2PV21KLzOQK79W9
la3DjbnWZK75mk4fjfFR81DWvc4s7RbRW6GsdgqecDgagowqifLZtLRdDjcdB+0O
rv8yegyLoFOsVK1YE0q+TYrndJiZgfinItDeqFIj9YTVpV/rYl+l9ZkOpiSRLyaH
wamZf2hmQqoQXY6meymLkyuSKpWIh+giHBMwZlUDWQGjZJiGR64wdvLxUHp/NLHe
wbLfcP9VoLYDDcbruz99IZHNATbS2b+tRxktOBBGSd8lWxQdcwVIFTOn1VcJMnVN
qQNJ4j55Ndu7nlZDvSU0J218WjjXnywK2k9Fd9563/EUK63a6wRTYRFtKDxQpEu0
lfBlrtQW0187G1sFTZIbhe4I4nj46izp7RJD/ou+28H8c0C+QKFZ5yZFUENrifEN
t/7t6zxIodKRGzIurBg2TC+E/jnhzJZ/9Y4PRiKR+l+uje1tUHvjnWe3GSLBMGs0
lBMFO7suMWK4iTaQpL5Vcy/RGfS7UScGbOFBWfPErdO4SdInnTvLdg5E9EP62URr
GSMiGgtobI99ELwwBzdSLRrZhFcZfxDohOqtRWEIxTwu4pc9d7t/CuJAb6gKhjK0
PJyqg3cNp9aYLDWDtmQfZUZtfVmwTADSDrTvJRFDqeADUOYyj4Uq8OR2bMyH4XC0
IRxHGsW1TN4uAmjcZbKKaSotuMoUW4qyuyyYTz+aDsQGWm7eunN2DCiC8MGErAsl
VapcDwEruj1yt1/Td81fsW5wKh4b8MRrnfeGt9/RxTDroiKLBd2GShDoMqnkKWjT
7qdEdvBVs0bxMexx084tP9KlmTWb09daupvE9DFiTIz0T2HN3AgoLe1iEU0lmDRn
uSaaxfsBpFZ0MNt888ISafvzWpJwOAgpVgYuAa1Z+O61AmJ+4z0b43zcnbVqSCuK
PVDwa0O0zJTIhGKpZC/tCgVogN5TfODDvyU4XZ3OF3dG57eFkbP+Y8po1taVc+dU
vM3pDfDZi59GJHB4dl9E53p3YQc7QYNsmt4Fb6qpMmDFMAnpjAzO1JbtP1mnP9Wo
qmeI9XGtsCZE6Lh4M7mg8tCFNkEEGrqIcSvmMfk2uhaTF2Hot+9oW/mK75B+l8mu
sDLdK9WFdoxFi7z1AHAJ+ZAS3CSuxWYpw70OqczKKfAPEyMvQ8xpmgd2L3vrhnyT
9yH1J0RvDUnSCwJIcKLnF+9bw7QX6zFNcJIBezbWaEoxzOCBQo3Tiz72wSqbRSCK
e7TvB5MIc/ryhpS1+MjnngwOafz0v5BiJhbl+akO8eg7Z5fp8eB0Jy0UyxJfvNS2
UiCivWzIvetPSzf3Q8imWtGolHsUf6IgqgCzn22WILr2Jcl24OWCBOozF35cIbFF
Ntqc6IcwkUNzXLXcdXBYDUCztaRFV2pIPTsUvX26uO61cp/RsRsmgCeL05cKwE9S
oAZvZXaUcl5qjwkCnRh8y/LZnnm++000Xdn7kkX5TLhWkgem601VTlOg3p6ibKYP
gTpo3w6LoLSW+NU/9ApI1HhzXfYrBQHgo46oRTO3/A6kz/eiJVGxmudgrVqXTEYh
owb2lrXxg0Ej6QL9HFdFc12TEs7I7H4yvZjb+zI1UrlcuCJhRJJsQR5tqfaGhdW2
6Bouz00i/66ZyZfr31In9IYO1aWcQprE49RzIuXNa7PMeV766PFS7lPswlocDYO2
Nl2+LGr3+sC8SioeJKSnWuKyXm6ADpx+7UVxeOjaJgPi4Bn/AAlPYhcrED6JFEkf
cCP2dTOgqiSk29UVWjr0yKJTEYjkAQsgnoMbnGy1FssJbE2rejgwcXf4RpJFKQGt
f/cvGzfh7S/A8bmKkvGbV50ZhyxnQpDi/+1OdVjm4saoOGlQd/kESU2F333IO0Rw
2BfSD6X2kM797RURWKzopPqwLlhV5Hmimg7WvRa4S1+Luo9+xOBQOY2L3i0uSwo7
buIlQFmfhPJZWSGdmr3uRpePXx0W32NDIUiVl3REQALwTQGfcsoCO/QFEFGxSedE
7H0LkpQOqcb8tbFWCCvqfzGzCMkZBfkMRcFb050QouDCwMpGiZ4aKvDcM7FwKMkf
Id+sSroVcfg0g/7gQHlzgKe6P9LE6EE7/MVB7E3E+XTXwYOnL/iwgSypLhEO2LGl
DRPkZMLe2hrYASNW9hNDX73wTvmu7uWmydiF7T6j/K6NQYeA+S9fbrTVoxk2a4iL
Mf8e9srqxt/s5pCVt06BYm2WFIM5r5rNEBcQYMBLhhBJW3DydgUv18SnFYAnl5Qy
r7aQ5KGAM9v81HkGSZlfn/VfAyoZP2tIuSRd82IkAyOQVR9fVvi9zO7lIYRL1rg6
nAkU4G92wZMuswMkomuGo4uyrz7kg+va+i607PSc8qVFbcTzoKpVrcIVAVS8Oe5z
/knXARWbC03RS73rNuZD4haPFek+8DEjjiWBXdOVMDnQAiFOEQA8pT58YUW3wpyr
A/bOOLLa0IizXBQf8980ecqNzQs1YNYbIPOvjvfIwXLMOg2bGSR+FoYO/LqN5vK7
C20Mb2CKEZ+4fJ6uux3WaKVYL0onl2d2vFTzccpBrIUUh+4O7v3uCITOC03OdHpk
xKjJ3DJ7QAjTHPtq8jIHCw/4dAXmiwY4LlL7RxbkPdo7dhKSvDT+hARDwvN9zqy+
cqV93K5vLb5SjbxgIeRNOFN/yBGlQ/g6Jmu4mpUY6N/WqZjTQ46f4oNJYWJUfigK
QAd+E4k5udP6kEm/BvZajVoMN4m8cqIXBsbeVpEkih8OD2ZaqwMnItDzEG2yVT29
y/Dk0GSyFNZPHudfblRP101TmqE+JXPURxZ/Rt9CmMmsj7Yke3sFShqFsHDcvYTA
vaAHC0qv0DMJz3XmXMd/FAo/htsHgWvLIt7rSA4cYrkXa1T88C6IxawxpGldJe9K
sTBbjYIgb41oKkV9SKZuFu+xhgVjkJeQ+yAuYl5voR5hXuKvOHiGX9wUPKl5m//k
mcMlVyRD1F6PAhWYMh0RdAYpZOzSLFnCxWFWSwdSfNtNtaL5zkzcm2kUBpW06SRs
wKhQnBwXkw6wCc0Ovj5YMqpguWW+ROyQ2BSPT5jeubiqhax6rDvaPECo5JU0oYBO
FbypgY90C5xcoBPmSqyf+yoRUo8rFnyI5DJ6WWVmWgzB8dqSKYhnyol1N8cJr1CH
cuMeAVczo6Vqyanhnx+Y4fqtKtJE0rbZht/eHDGdAnoJi+oox70YpY8erxy+cx5Q
bc8cXP+JTZIvLuioyfREZuwnier364++V/VwcfqCJgGS3GABgekO+ycYO8NjPZuf
a1+ISQ0Ql9HV5gYWF1CxTsk/8O/mpg9PWG++TR9CBqWZ3GL9n4w9Y474v7/7FuIA
qNoOZGWsiZx9EfaFQofBS0Io9xOhkTgmnqkxYgFqPq8oQyINUQvUL7H3ufnf1heM
cDPzI1zMJiHfJMKowDnrpZsmwS/zDMHTgs/BLXLYX9VWqKarFCBS5ZKPgGsewrq6
FsqdpsDhDrXWXxVHMam7L5zn+LbNnYB2+gmOAEP3So2WGnR8DuC4Yt3lwI4KhpGP
RaeZEny/RaHeFckpMsdtZyzknEOIuS8CjK5SNOiw9esdlTd6+1pihae/Sb10kooM
1aGu4LAu8r0nYxXD4zhb8V8f7j0a37tgEzaCb9s8tu+x+Y/ssX3vEyzwsRwJkgGO
1POO8m4SguEii72uxuVCPvrrqcmk15A9X6Kbt1MimDfOKoWDhoo3QDtkLPKBmX7A
6D8CZ/6E031Go0gkFNcdjWiyTYUxwwH2uZD7DYYmq5+AxiiPzjL6sO1/gBDqE4ep
TKR0yQ6axToFMPxEN4dnKXjh2xfuOUitF2JMkrHWkzGkk5naDUhdGoUWOJOdPowB
iF5RsBFSoUBjmdPG/lLigApuAiwqezAEX4/Vv7WcEd/YBoPDO9gQ7+HMQvIuQyWP
+Ax+CZYJYrDtWnI+4xOYXTLMTX15f4JkJEjW/p2oFKhJUR2ULUPVKFqncVaX2MJB
Z8dbLNzM6J2o2ogKOIY2o2iwpWmE5AdEw+B1brlz+oyVI9jkFTQbpbt8k39wDYs+
S4in81PSBZX+sz4gB45OX/CJ0a2/tYHS19qLjjMRgXYrPP/LEAr4copxx9ouMb5a
gm0Gi25MiyONU0mKmLjlBHGKuPLZFlZLTXtp1u6ziGV849rbdVeYVm0PWg2wZFif
/uccH0gL7f1NX80GRANIUlmivE/KV/2tJ/z2Xfbr8R+B0pv4q7eztHW1V6LFiMnV
FDeBI/cmQjDaHIZZt99rdFaF4XYSvmnKAsOBzRxpHGrpEw5J71/ssgg1AxTNa5rl
I6Jz3/fBDXCXeTWCLClIuX9LgWTW9qYZ5UxWZGRJbPv9cNXvg2520reJFBcwahB9
S5faT4I1dvf6jl1sOtaOv4Q19k07QKxspcCJMqqRHmp6FoUaTgY9KDh8asPd3glc
Km4C+j5VvrruC0mawHf5JNPq2DT93t7smj4l+vfBHWQ9BxqhEkuY9MOSWBLCg5kZ
SW895Zu2XwEPAWOxT0qED9dsPWxVbJcQd1FHs3jmlBsaj7P7TxTK4QCdlet9k2pi
oBaJQiB7xsotGDiytIMb0bTdBRq5nAEiST2oirCu4/nR+pS6a2payPntXsc5qmRl
WGAfj0cny0p+8gy9Ta8J4aXs8VQ/8U2SV4tv0MqUDP36gLrWlk2HX8OY9Cns8oB2
JAKcrUZZkXGdYWj3oLB0ijW4tUIFH6PkZTb4pp3DC1/hT80Q58vJ941S/VMWzbjz
axn62ytFKbIWPD3QB7Dd+GZwoHNvMO9saO8pUf6Leqb1ATXusSkRmU8XAWGYttYE
jZhyh5wzsRBh2FGOTW6Yx/LRmWuQv18rbN6g+3W3W8QORjlLDz8n+5KCEI7LXjJY
Y2UW/5EIag8Z6QoHiuR6sTrKihqb4ZfR9zq78yTMIT1gLV76IAqyv7fZhHhMrZyy
HYdXyvH+qCddyyBnXfy7qYKoasddw5WSpc3ufzB5QG85EO96H94KC6BsFTDyXLIe
GGc8nDC8zAFpbRY6Sfn3iWU8VGvN/S6BX905aBVXyB3gf0LRT+F1NOvkQdc6qv9P
cUL5MuO68pTtJ+JocmsbTY4w8qeQu2EJbU/t18U8uF6ieYXfjf/3NPclbCLRudNW
OWxZfYM0C/vZ7p62o8FPoWWR3nQyJnthm43ee5BPjoHG8TU2cxc0ilO0pAgBkLG6
VjJJ81HDCTt1M++L2W+aqwktImMTeIiKkuMP5qdfdI2s2z+CUKxUsHQ8n9JrncYB
hE4P0oqt9/Jh0PtTnZTt6tVBQeY9JHp/F+E8UAN0SZfY+k0N9lTI2Iw84NFBQaoa
F9BRYXIhSMGg9adjxdo8QLiXatSFNCDsvfdXp32rspFrItQUXoOOHV3w26m1LzmI
is7caDWrf/RHMbLx/6HVGpI02QgGQYjGHVjMjpO3tfTX1qi06HRMChREC6ZAqFJm
FCuB8DSkMXpDIe2QIPWMXMpAqkAooYzESd4XcR77RR6tUzQq1v4EY/fmMKSoYxAu
baGhzcBhxcvUtky6yn3O9zTMPdI4TQYdpAEZKlGiC6SvwhIrPsongYs2DnSG2ppG
cPyFFwys1DVGivZeUzYEgpnXK1IgXWOylRA5AxXJ8gltH2fK772aFZJ605Z9LV9l
I1bGnkyfIw7EM2kqmxzTaF/J4IoOCbroWrsSZVaKu1nam7xcKg25a6Yd5bdth07d
oCBrYdIrbmgd9EGfKadaBiSBtJaI5SBcUqW44+7sQs2DicjxCciD/dwZ2J8g/hlR
vtdxjSl8tMsgw+6GkCHdZDacl8O+n2+3ZaE2k6iYUeH+hWMwtfAx5cCeL+tcgJ4T
hVoCVNSr6yyd5azm3yIAMtckmC8hE+UMF8hiEWiPLD1d8uARVK9MOZcu1BBxTXbB
ypDtgW8Iyk0yeoczVsWhqgfUP8qDS2YIMUb8ZbgMDHMaqbxIKIe3hXfSLYWsOzya
UqjWmQ3KU06F4ol51V/tKxPooCA5zv9qfCGRjJi/PHi7MexR1P0qzn+3JgmHfaA7
ziQU9FIbbaf8BGb1YiH4G0YvEEq0iMO/0zzP8H78ttd7yVN2ifPsZbJxIyXOO/QR
/P/Sy1JJF8mAnl/X2MPiRFlKnj4TC9ehADhjSBrNurKuJ08p2WA2OWzpNifK9stD
7OzNoKkDchah9qaOhUNGSzhc7+lNRfKlZ3hPAv5hsDN4TmcgScURJxFoMOW28TEi
Ig9yAEddfkROitXfHinob6ZpnD6bO7BOQUe8U8wVhBSQ/83DoyPcc5fdpJVhTQB9
9rs7CvsuBnzsj33P90o0+QMRE3GJoxK42LZUMik9Hz7udfQQCrEOL3sCwD/eaLs5
BQXLnUsQFfFXKO1CkustSMFC3mm9POiODAMaN6ja+JAB9bJlO2Tqpq679r/eMXNS
Iyp79GguBLSaAahHLU4e3iMDwkEkDxEP4OVpowqTBld+cJ3kZ8nkgpUNPrqwoU45
M6VIDj+o3fXXQvFIbI2wlyn4KG23kZkWG7iOSKvO2N1l1l1vNFmTNirtZVXg/prv
kEKmUqKSkX5nlYC8VcbyPnVyEiaeH9B/8aYfCJT+olTw8dmOcHNh9exrklc+11T/
UnJpHHrnimWYtAQdDRzcjf7DD691rpUJKM0NRbKbr50lfsqc8iEx1vZ4nMt4FRUP
tZRj/4Pr8EQxunmsV5d6bv9vU4WuGG+p92WqoyHr7NKbtUwbJZlxr7FxNPvQ+leq
m1/bF5MA8oAeW8rq4aSC9nnf3LZG6slumg0dXfqhw34hFo2OW5+puyHx2ZKTQ1mj
x9rPEaxADMdOu2ydUNXPlDmUwWmbCXXcYXbnle3RSYSaxvpTF9wW0EYA0rz3SFd9
Iydk/xDjEoBoDSsXYY4poHsoE3yzENgp4qCm9VNJ6zKvMBqyf8uWaHPTQQ0CJ7yv
7JDv1mt/O3rLNNNQmagv7PdEyzwx1EK0/vhU2wiHeZepW6SHl/LBNdW20Um0MoJH
zahL/6U2H5z9o1JC0ore6K9zAwtLKVhfOhbz830Xs9iivHS0zPcZdXof00KLoc8y
r9nEj0/XN+oJJnARASZBZdZEHPTr/nk2mW9tb/qDh3Lp5nFlgmzACcHMdGzy7C8E
SgpJdGInSs9wb9EQ93GR+f0sV7aP3pgvpMzJnrNnxVa0y6c7r7Cu6zsQEtaW1GtV
D9eGB9pnOMeCXuA6XnxizC5TnPd59oVyGVHI1gUttzAPKGNr3yTquoofVaNW+STv
NpJ+6m/FDLOxQECKqDwPt159igIymiykrNdClD4fnWAH41yYE+AZuA0UK887C2o8
ms8VORYVaLZPVmocrc2lQfEYP7zDzGM+utms8shmN05G0dV52OI5nGH5ISgCg1T3
44jTcc/k6jl8sSV6qAsf3CEbJyj0LCr4dBFEIyvs2kePnpWjCM6Vdee9+eFMK0tU
OX+McX1Wc17JIogg+JFwxQPrQipzT+elGSKPOKzTzPeRZ0HWrRYMTszSJUZsrChP
KMHb1GUpjRSlMDUo7n7M+pQCPIrcIosOxvgmYix7CdAXaMfsc4fzEyv6P34tLYdi
Lgkdf+50r9zea0LM2DP0EA0ncfVQNyeFTv9CxKa0YU5DV+GreIIcbdfR0BIbzhh9
a4vzcdw/6iVhxSbALTY0Hf5vKxYH5InDXV2kIXY+3fmT3fAftJGMqeH1khuhpdHu
NMlrSikQ/Juswob0miKGy+MiuMOLZD3LYjVXb4EG0Qs5gCKT6c5iJm3wW7d47cQ+
fmsFHCelB0Yd4Jb6Kh//bCS1VGfDK1wSio6i2WbWT2D2E20bt21y5WAEkM5zg02M
xtGusQbvEMOE3FUjgrb8HNYGDcFI1mUOAbElSl/eF9DzebhpiNbOVc53oEYfr+H/
rnaaw7GXNqejhMcN9V2NKXifcYD0z405SaHXbG5g6tbWHG3zOMknK5Ivk3q2hQY+
RKCe8RADmXDqzGSyWkwqNO+ZKHIs4IKwnwS9iRY4PStn9bn8MiPQaSVQ+vZP5eVc
hn5UPK3ytC15iFasu3PtMe8eUGb95TB5ruKe9d4nc0DzMqvLQ0ata/Bozpg9yxLv
7UlgsKaBvLlXqjHjMaEhmo04ZSMEe02zxUKVy9MDqnP4Us7LcTYjKg0qu+6kUMfX
PDp1HBFe/N/UHGKGGflWnp7Dre23kAPVy/aDZrfYw8lDXxo+6ZTjs0jizYEOlC3T
yGumHZIC/tcVdmUaa81poTqqopACHuBftCbTn5g3qkqtluKddwL3ocYP8Cjwmgdb
60Dnn4cT2DSH0Lun3NNgD4wT8tkGHotv9mC8GZI9FM2DFFf7xrSyVRtNzQbzXJua
Jfd5/BlQbFaeJACAWwhmHydjcjPliQ1YCrZRx3K7tgjW/prnmH+eHx3QKbYtEb+r
+fPXi2n1w3lb0XztJocM5AHnc5ZxD5uBZd0SBRZyJVe1sX7JuAZcum2Kpp7/YAr/
E3ANMg40rzYQ3T2L7DD6y9xsX5CLf1Jsz44+Xfshx2nG7v/F5B5kpbJHjM0h8bLP
6I+voGBxBqk0VPWiiKUufPFNw35YYCty7uKnWzSnoV1es7R4ZD+5eia7rqtT3+TD
iqd53WHbm5yR45Y3swvOYIje06qbGy+nzDt48H9jgUQNVrBL3URDTirbZq0hgM5I
XE36xl/RsJZhan2Ehvz3ipYnLcD7Hwj7AVEa1Snb4hzpywRRzYbn2d4kemGtB+/O
E/2jBJrBaEhJdXn6ic/tc/sFNWfWUH3Ed1ASqS1xRA1LU8xk8qA2LJpU9fFkBfkG
AC1KaGzKnQXQc9V6KEeBh2J/stzj/E1lx9fgc5q+4Bisv08I07TPeDjtl3UoCm4/
iFgkZa/OhaAM0SFAPVRzK0t7mvOWFWGSj3nY7izI+TPpvKpabWvrkF9QYTSnGb+Z
RQPmenBWG/ONDuf0wZga8h+Yzu1aSq79FjRkJwQ2qVwbGHdy7/3ekHBd4w8kizIm
jkN0J3/tH6OHWTCPejkWaUtDPrAdCfROno+KQBOL6MABeOG8kwMy+MUabbVtCCDP
ej8PHL8fnDHbD5A3UJDQupXY7V9L6ySIdy7j/V2omuCSdsSY0iMBZoVPIQyhd4DP
Iqwli6j+dfeUECff/PyGBaFbBiyMpMvOM8+F1+7Q0/MyVsYiNxrq8T6DdqADYe9d
c1rJOjR4tbUcGCmERFSJ5vxFD2ZNRCPb2u9EWHA4zVhrnA5NQzziUL2f9XelfhNx
F/r6ELFu/NJyBqgoOxSgo1tCqe38sXMY2X6IdfEJNCkxPTpTMDCPcegw8V4g2yeb
QNkUullFbkdJVmk6drdbm78pBzRjcuc0KFfcsUcisuoTHrrTl5bpMraYA05548hU
YotOe2lViFn/dstqogj0x9OzvH0BeLQQ+cdie19k39xKGL4MawF/si7Et5oeqJ6j
jbdi9AUb0N2RUaixAhe/8V0LxxX89SVEQ6b9b37vTptRyEc1oBAxoLon2g6nF95f
MOoEpLNJ3ZJ6h9XKhtPRvEN6KxypCfuF3qfSLbo15I3FgJG+dNDKn72Cb9hRv4mU
/QUzyGRDfm51o7dAY4LI4AHh+E+hkhn92vajf135qtN/ZnugCtjUly1w3JRwhKqM
34DQclrexUbZeSrgdRom7FgP3LdIkcvuNN8RMDiq/q19HdFi39e+Ec61X8VGWSmG
YTFGuNhxrTlkvBF6z4S8fSD3LTWoWXaiFPrKnc2j+/FY/aggqYVh0VkSRTGXrKLs
nbog85r33j/oPvH8RNOeqSsrg+KIWgJ2RNIPPH3TpJpB98W3Av3IK/dtnklp5bnP
Xyn1QvE3jdBJ8QF/Xq3vq2Ak06TTekvHn5PqVsiB4BMhebVN+B1YneH01JG2q5D9
tIeds0KWQSwQN0nS7w8h9n7KyfU1WlOcXOuYcQfAXYmPzYfORfXlouRRbDCg8kQI
+B1RVtJus5XtHizm2N+iMbtkqM6Nvy2LGNyqeJ81Z/kdED0lh7ZzD9w2vGk9LV7N
ayjs670mwaBULndT/3Uz0JV0i7+/oQika4geVEW/5MDkHKJAfEcJa/TNMxePH5tG
j+pHNgWNfjSg064v9E1pSiACrieBg2/ikvuHMGS3vlY3MH+EzWwgx3tKBMyo8LW3
IgGDM3ENt4sEUlhVXfBgRUlurQIA85Kx+/uAIMYYfzgs4UMEVaDooEwWScN3YAwP
2YqaqGS5+wR4stkklPbV//2NbRO+v2yX6Zx2paGwZcnKQDrCRCrObGgVLHIqPScX
vXc76iF5/jTUcplWJleKDQ8Cr6SnjyJ0UXKzvGtZRxE=
`protect END_PROTECTED
