`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eviZVdwJGxArmmFI3/9OWWvw9zm12t7GhnR1WQMeZR7LApcbar3lR94HpQjLyFgB
dJDpWph+4WirGP0QutMVQJV3t+l8I9z7+h47A61v/8tfSKofOoCpr5Sa4wSrMeDt
yQUakd7KDPg09XGz5Os8Jav78L+jirNjruAL25XkST87bhltI7Vno4gtDWZuvDTb
+5v3anh5v6NVISyhwY/b0cds+30ChrCilqjILd+Mn1/inD+qCl6zMSEXGY4p+v1L
1DxnhsSsCTKKt3feNgf1Q+JwOa3azozKj2GhkDdzcbXWV+ZZE/1A3SyQGWR4xKM4
F+f4d5ozG+nyS5DYVFzoSQmVunT2JcSNTFPN8WVLMCAzp5yb6a9PowEQs+Rpu2LC
7tXu35aZLYzxtcRTP9ciqAt7pf02kcMzIER3Z+Fexh4sogNUnNBKR+l8atr7Avuo
OrtOn/VNGdd+K+PS+28TcUsn4zKdJH9UE+88uPq6NaAQ1mC5UFx3X537CW7QAGpq
QiiZhcYlDgCQBccm+DBS0oP5JYJr9UoY0RvNwLTtydwagNL6npbRB1lqWgAfM2oc
mz1SBST+DUEU36gKaLYNJmbEjd76Nfj7joYfP5QJUNhlAumUr8Vzohq6jHhswUMY
6A2FUk8j0SBZeUiPSePOXvBd6blhgxhbJ8o5iXBzfkfgEvO965r6YgxLLatut4jk
vIzzMQ+SxxZ0mMCTta45++A/EuN4LRkc8/C2PWMDohjcG060iogUdEp3hgvL6nkC
rXaaOCdLlI0RXzUAGWCGEPg1guAUdaW8QvlcxLY98amVA4DNzG52GBqWzoyIsQap
WoEo5LbUaQ19lcvHDfBFDprHiJ/jEifuCiUEcjueYAn9fBXqYqIhp89RL7AMEzMv
yr2hPZftE+WvC+Gg0iYBh2ZpnN6BMaH4iOY0RAKuv8qfmFGnCGJDcGeeMIJdyxO6
9drPpOSuXWJ02RL99JW8Iip4D519FEUhxf2b69vHqffrCQAFc+kwMDvKF5uKY0LB
jBYLcYnoF85cqqA3mCtZ7ef0kzVsiask9wGaQRpzRo8yR43tOWhOgvskp63Z5ixG
IybAKwZviGEEy3gHXqhoTlAoI5S4d8QixxLLssoC32zfGKtFjwCw0jXJ+zdBI0DC
lnE43Sx98l5OspXH0tKwf5qs2wGmkQD886l/jMrNz/RCSpqI+7xr6mtUf5XQFNg/
wV+XAgrsaqrUGCVhUzxZorHEhD8Zx5yKhCpJJoiBRiolfh0V5sfXOQKm0a+iWlhn
DSoF0co7DfrUfQTjsUczrm+KKdLG48moek8FNjpV+DdKHyBruJEZqHdqrL0D0+j5
rMcw+tDuOlQrxAYJic1CaDumZGfY7117owK/oEQN2OzODcpceH7a6u5u3gW3u50t
Cal55xHJVCIDt0QYPhAVSiUln74iHTUCduWNJ345t+dRS4JfaqiNefdrT/NNAjw5
TYtfwsnkahfWBjLZSn+UN/T/W0SjY7BlVH6gVzX8ZyNJ426/kdUxnDTixWXE6gIZ
eWWbC5ygzR+KIZZg7mFttd3Mxr1HzEIoQIm355TdW2W0SyRnXM8kgldfzWI5xLfc
rOGpogt13WB7gAGnovHBUX60yrYesL9xxgBknXDb15zL01nq2O/t0CLKf1bJH+9v
u6I3qwA2AIxMjnuIOA4HnH/2BlDDur+clYs05zzIEipV6QE9rrWL6GJLrvHb90RU
IwGdXYEdHdpacINCk0+3EPpYLLBlUEqOE8nhk8fWveEYtWkUNQb5QqV+exNeqIWr
248EdOmM75//XbUounctf4q9uX/rfZpeWUR43dFC/q7NHXFoBCuUbnMOrntjNGxj
LlZuOZhzt8QtNtUlTrKYP2wAlZnqKpeET0fMBMPZq+Wsj1jUW26XlvPiGgCnhDwQ
oGAhCxiBq3KSwQ/aL4siGigKMEHzcz+1/LVVgh/+5Y4VJcLNJQ2vuxfchvFBWDrG
AnxBwu8eGZOcKSvWgUPPmojtoH4pThTomoaArLjbSyVGmGKBe+pRgyVmp5mp5MO9
hVr/DJ5pUaYcwWfHTPL8YBwO5ZcMbQc6pLHYn0s+E+jjgbybGOoxgPLf4D/sKO3n
IjaFZQQCVZOR1qi2VinlbdmioiwS1cyPY6qD+rxUjCCsGmgQ73JyhC6I2kDYcZ9p
GYCy8dQTNcYl5JAEBARhVj/985RF/CT9Mn94lgYNfDDGRZR/fnIJkNLxsZKGnA4d
jq1xr/Mos+JfmJcgLfqi6nuIYFjUZSyytX1NMjax1Q7G3P1POTigY3Qcu+u49oDx
9WwvkGHyS4L5rc+gTYURsgj/A3DAJqOCdwEsUPoLt8uw1gsNJ8JmqPLSwtu11hJ5
fsrWwOdx+OhCsuLCj3rVVOPyC80pXgjis3LA20kKz2iPz6ksOIK7vISEgQ/hlsuy
hwRRN20E691gf3QPEaFCrPKlAY24ubfLW3/63k6c6aSwVkaGlcl2R1pSxk7nEgms
wZZtRMnPzgXZmvfmTMsBsaymGK4lEwfehhdL7YEVWRT/bAasKrK3S72p7pm6Af7m
7ekCn6FYetG+PlrdNa9YRPLHwAJSqv9LZLgwr3qZFF7npx8El7ve/XT/xJPBwszX
k2DDFmhbLYvvsjsKZr/M19WFGknZCdi1xbOfChh+GLiAJuh+rSiQI10+93dFddIY
4rC3uiAhCb7ZIFI4nFA2GbGkdxNh7QN7XFJLzpIM+zcyTm0AeLmcpBEW3T7swgWB
XdA2FFqmI1kSO9+b0D5UVHTQ++uPWuDJk5wna4XdyNjRUmvsNSoR0iI879Z+BnnY
4NKGgEVR70gKRshbBDmEtvXd67/2lpiTyX7G06+wDoMenK7JzogpUxTE7uCdCB7+
ncJmMO2KUgLTM2TAdIkrqc8bUfiS+gM7upOFacxAEinn8+8jIMdHzDTllk7SLvwE
eO0OMYAGQxQJ7O1fvqlhO8S+n1Ujp5JBp/nz3VmEZBAQ2oFanBasstiKkq84pphA
HEdZL37UYo7qwYxmpk34505vxFlf/wAnjRR/mEWeAQB63SAApSMptadIstIrhIa9
3QXoV5XXsnFidQ0Ft8VIpjP6rsi0KY4232HItmaSrLgNPey8QpHI0NTm0fliVi0M
JgD9tXnBHiqcDvn7YXXvXll71jE692yAHcqroL381LlP9pw3sjvDmp/bVxMXR17c
BRKA/y+3mR+uxWcU7QFNEK7ZrUqfAc69KK+Pm1yk3X415tnnh6smaL4sMTUBBVS3
EMMMKZBjuxvU1uCvWkLnvsYsadhCN7UAyNTfOBNq0WLQau8RtpSm5oKMDDr9hDgQ
kgl2PWzTC3phxb+HLVPnUpXVejxowFympzqBbl0bL2XZMlu5AJzNjLFU0H6390Yw
9a83JvVfgOZ8NU2Bv0AfFPOzXwCrO/x8ZeKLK14MGmr+PH/fJPuaZNu5wfkKZgIj
668KXMyqLHmwaWoPXF1kX+mUi2UA1IpNhX3y24R1rve5x9MXtEP1mYMMhX1Pj9K6
0YZ50SBME1U2SQ0eVTfJNk8tdokdwv9TbS7+ZvORHWQWkJT37UNI6gQUrdVIocq0
Uqsiwgf4MRLNmqVHCIESIIWbpGduc2VxH65Y0jVy6DuBBIirPRHJe8AlCBbK/gbT
BMmADGq2g1VePYyx5CfBW6HXQdgfx7I3YL95l3tMFZd98thB7DORbEDOwhdkboXM
T+Fgm2pEFgPVE2u7pAwqKwIRR8asC3PMban6aDMskAFSlsNwimwf/eGfimMc3MGU
uzaFs0qxV688NvuA9y/p3wATBcs6/B8Y/vrBefqgvQsW1ED7n5eVKwRR9l+2gkub
TLj0vWo6r/Ys02Z1tk8JE0KfFIGtb2d0WtRrQanDhuVhLgvahVhMSjNVLk/yTsNY
WOXGUyiLQtxxi/kfCL90P23zYECvYM9eP8ahaK0Hlu7dSqYcGdHxVWWO4/Mw+ASH
7yp7lGTwmqDABxb6f0/v0z6N4smICocO4C1fIN3NVB7v5eK/SVXdoYWUHZ2sCkUc
vknnRMcDti1u3J0fJfiOyqwMrUM1e1Q+dROp6wF0l5qYUOzjRBVovqgY7Bd52fOP
HhqhollvyafLlamgxU3rMuJq4oUxuIhDhybDTL9o3NR13KwrAgo6g1Gr64wCMkz0
oYf0EE7dIQvXh2BeyiyHMKSOGg6UoadeXFA0946VOUyN/41y6ievR4tQrKARylkE
6vgCICfPDK1QB9TVyRrnqMpv4OGmRvSCRfMTTOQKhwrUlnzmP5BwXaoURChGnRBx
WU6SvQsXVICInV21zvLHQamLC9B6l6HaIKy+Pte0GI0tqJblq45WvWH3vagtfOkq
4ZF3QMU/O/sCZgbSfg8Lh2r/RubFj69itzjenDy7K2f6e5U0j2Iar/C5vlTHMXKE
ewQfmv71dP5W7tA3MFxNG5owvnaf6yaUJEedTXq5C+DnmHXaRNTC0iTKvn7NIbVD
fDdG1etkj36gO4IGEW1vl/YcmOhWmj/rmh2kRTHqiLIwB5timVU0b1aMgQgt+Mtq
BMsyI1jTyPPSveJ2mxZ88Ze89H+bpNX49k4xX4FJfh7ZnvWjk/yNebSDLLtpNOkh
dlcKilTSFD8c6/LN/+6L9fVHZZmMMq0ny5CdZ6NRUNWuI6tLgYDvoTUMXfqiil44
bwJA+FKQhkPQv9S81PPj9B979cA6huJQZCVB+NCQ9FDbl3zYa8WuiXvmev0ZU/kM
v6D1d1+0jaCWz7CHSILFijEw0hLfLH+YAuutQMB15Lw5cbQcQmOVIqtNkXuLM/+V
9XJSE5Kb2ogdNDnaBBBCrwPdxH0FpYTUGwuQiFqmBoAY5XsX8a9Jad5awBIRwdzz
KD13KO+bW7yIeRNQHQEDSi7WzMMbfsCyw9h6RdSedOW7sEUfbuwA1nfl2bsIX+sn
aDXEdi6b+/+D863Je6VrVSflfbLokImy69X+buKlgA+qCMdqsM0O9cu9ACkhehNN
RQ8x75QpvzXaUleM6RAamEizN3Jb+p4d0aZwwzehCiCylpA/WAfDtpO75cRfvpjS
58beDFFmKxgMR4kmOmlkiysjizKoKuqeNkTE113WO1ytS93wR0Ze31mDi7ZB5OKu
a3tye2txmOqGH+1QzyP3cTYFci7mfwmBm8HFB89ifBqG1mCfiz1T6G6wTyN2Ye4S
VYAgLAGB0EsbZdSiemxIMeawNuwe9Gg8lGcOtoIeMmL3+x8PnCsv4B+/Kj5f6efe
Vo/zEQ26uozdzSQQ2biMMzb5CVvKRyak7A0nXY/ar3GSQxTf90SuwwR8INze24qG
g/5CtS7gYmrw7jUUcdN34PBaUoMAsZxx5hwAQDZwhiwedBqzM5/9I5I0FkQPbYjB
apOTnaAuXyHRB6ZkMrqZyYluZOrZ7A8NonqbtE//pbNgYu3eO1vZzyHJg81aLyMJ
lduHD0EabmDLmAb8DhiMagnj8cG02dQ0ZOtFMMYoum6l4133QBx51xrDkkSXGJDS
tyT7yWmNzd13tAzI7MUduW9rctuI75mKPkCovgLpEEVqlD8JNAqlUaidzrPowyCZ
6SFneA21EGDJrz0lg30mRLbeDKW1bsfZdA9IPqRKh9Rd7TVn3kR2NlfN1VGEZ268
LjfyY+4rOpTXrxmedQcKEbrfkVv8KCt3ovC0XqRyRiAOcwvqvfkQOB/f+jxVONvD
X57DElOeRhXFWRg4dyXfpUa2S7Nck/iNC2eq8fHl1SYpb1Esw+0t1KogibD2MJla
CUfc7/QiQf2E2iHpFsraCL3RYWyyexkwNaXQUjYKa3duWOKDa9sPE785R/addo66
La/4TUee1Dn9hjANQFw+op1U9xZbgQ/ekAr6h8n3vk6ILoee12AyyPEijyO/rhlc
TWqkjqLFku31ChwdW5osQ0+T1C677gLraXBgJoy4invNb/azerUYD3t8yibfvhPG
ZbUVC6BFTDtWPHcJun5GPSv3guVW8TFoCJEbhRjhVyJKRM2vJzzA0mdMa0uOQCM+
T/hGRwrNRyJI6IxWZ+cR/RtsCd3TL9D+6W0a814pZtxFTaBF8miuLR9bl51PADlj
w/eV8CpMF12XJJKrECHr9zguY1A/KZ0O8pxWRjMuwCQ45mu9lxtyvP9oof4qqadz
OpX/EMnT5+u7zec6RjiEQyxrS9xcQvy49Zk8Fx5Ykt6AkXtba72fCumaqX5TlNYd
IThqKfOZbbUK4qxzuYrMnLDhRsFE8aJiL7GVCQa1CPDzI4uH3beHbv88t7BR2VQP
72OWjE4XTj1frVoBZW2RymbLkLNKOLiHRrbVApuktyWuHFGyi23YpHa/SESKz0vK
Apul5wgCZ+Th70d4LjLM1wtKyMbkICFK+QS1kx/VkRph2lfiEnPDB66eLlMVIptV
DX+Cu5fen/wYmiw5XROeLvsSHF8if7J/bedAi4ljDxLVhgM5oIyX+CAGkpSD0MlA
ChJltTmHtPaRQPKjd/KSRGg/m2jgoHJZ53PRaYtn8mE71pHB9nUZls1gE2ROwzh2
TUooJLt1a5J5P34Imnip38Qbm3vw7PnmKpifsGj5v4DP8PLl9l08P0TKYGAEpT8b
O8/c5VP69d/lChYopRR00tNetxs/LF985LVRqe5Ao3T6WvuW3bwd4Ml3m6OBwEXQ
/zXigHAJY/McfdJn+k+dYmUKCZuaCo57emlxjVF6cyJpdV0JrutgSFEEaxmh/z7K
y3m1bEoLFG9Au0x30zfaB7jGlJoBpvdBcgKWEwxHw35a4OLHK5l09cDvI+n2T5MK
S4cNxMMOUx9jOpJax7Hqgj6WtdvMaqUyv5+y280tSUoJXtQSq/fDBCsaUr+1CUMp
gXq0ErfP9BAFZKb3PCCTjFXJjwG9BBjX9ru5aMoyUwf7oTImLkoxoQOmZiyFNgwN
VYSdFnvJJi7L1wkqE82jo3q9FNqAnNyHGHsrVbAJk42b7cVq+2PL402qyzrvr8mj
NPEiTLJt7XummvwoIJXnvxOTYluySUj8VYjZfBCPMF8ID/PqnqSFKm0/UXYzYMMc
MacSVmuABqZOUZ45bwKIPDFCJY+ErJjYboiPRp/t+w6JQZDlzvnlAEMHl2lN2GSn
uNALnUB7FleKMewldb2Qp6Tqnxr2dg41snZU1cSg46j5eFY6W+LFO6alupdt6dkk
bzkcCY6qMijBn5M/9h9b2qBTReG2+jVp9qmtddGC4frXWdwGnWCippDdeGAruDBC
pyzk8thInak3hirb9g2P74YH6+WYYAH04YRpYKEhVXyQQLQBW5nhc8NEZCnYOLeG
T7fv1L8f3IMWbsNn2C7f5j8doAQHMrvDiTI6ETQYxEc0hF8uIr5AiQmKAwjb4sNG
ji1nHNUVFIHYRac0qmFQ+2ZjRssciQgHINK2pyw1VmpCcY8GBST131k+aiI9rW4b
VxPajbsK86IQGBD9UKt26jeL6kubPKAVRiwZ86brnVK+YJWPP76YdysV9JAUH83/
wotBCKGWEEwroMThbiTCpJkI8ycxwyMcS8m4aRfpeP/74Tghdu8u7eKKO+MhE0Gf
k7LRalE7XBqChOhqrGMfG214H4JHHi5z3ZQfDyB09xcaGZDekPjX6fHlwKoYOw7I
Xq2oQt5gqaz3GDIaAi4dKKqzZdTQIeCEF3mAScdP65igmNPKUuRTa59VI62vC0sV
N8tVwFDtTuHJ8I085i5LCXszIVVA5K4fWTMfO/WJaVuOB/8K4IebTxqvokDjfrSE
irGsK9Qb+d041zl1MjArkzDFk1cxgOpZlstwwMzy6TMPBquIoNjVsi/kwF9VVzrO
IW/IqTHos971UFa0fd79nBYCGA515zs1tnlVQZlV3cFTWlTnU4ozbd9AUqlVBEqV
AUtcmtVJsje7juC1WPcgEHyY8wQpWOXc7QZ0Vj8kEMEroewyu4LuP3cahOx28dLu
lSv7k+gfp8hV+NI7G+Q6izXKP3xfioHuL4tbQbj87vj3/vAhwtb9eEu7g6hcHFL7
7HlaRuACqM6f4cYhOj8ECY9rH0T16WLHdfGjh/BcqOswTL82zC9uF3cIFposlEcq
C3EusMTgpf9iNaLCnS02xS9KKIFm/b/7EgeU6iGHD78RcybXOTOyetN2NBdaIoDd
mIIfvBNtVi51829uXeIceWJjy7eZWGQsa/RaTcTzyvP3x19qrmGBbXa8/WIkb0l7
LrbNUAvSjTMOabwxhqw8JD1CG/g4MTQTZ5+E6GXFzyn0ZiGISqKCc0DspA7XB62L
dqq7NMS4yReFdQOd/7tnluKM+EiV3gc1SDNLOx+L47oXi/I/DeYvg04DbH7NiHyT
jtL+MVEyMAxoB4sL5YEco2bZq6wQ9/n3Wo4xdBcwXWbNGqMX1iC/s34LzrDMdjXP
L/LQptgT9TjD5++VQehxOHZpDPUtTiYTpHjoBDfNzCLrP1nn1eTe6cX2XECuo0bS
t6qtqiaKL9PVXUk6s4wTLHL4Up9PGROOTMfxXBFjYehK93KJIzIZI4jwEgzgfrfa
cmxFapSeZMQnIop9tJqpbmjfBEtKxB5xCGDEosQgNHunA6dA2/k+KmoDHsg6qJm2
TDcxIfBuqskNXiXIWwrEfuYHNDNCZonS/iudU5jKl06FP5jq64kaANhJDFXVAILu
gRCRTBT2ceeHfAI92dl/XQCPUZaqJSXxxIcjnopoYIxkaVJVsDVCNZ7meB8ZyK5r
trk5XkCmAcuiy735R7oc+MbOK3NBK0Ia649UjW4fER21P93d0M97QcpweH9ziWGa
ifAIDL4TYMqYBQ4qStybPIHoiOXFoxy/gqtYj7h4X9+EW3QBR8lWDy3eb6AKEfei
L4ludNrA8pthzJ427H6EDorYnVZLrmBIFsSMb+w5xIiqLdC/3KhsNIVr6Yboqk7c
RBHqTw/RRShyNCSiL5+Aa3BH81EVapXfRI03Z/bdRPZSvdd/oQPkmIt8v0WKl43I
Iez3GxPk4K3CW4meJmVB6DVn5aDXisLibl0AIZfd0apbEKtWmRlf/aqf99we7Ka7
F+l9zTkJ3uOwqFMODYha52UZCuax/YODevvgWL7FyxE4ZAotRlQmABTe7lpqoTgG
714ybaff46iOykY6FS+JzNhmuWlaZRAhOZ8LBO1R3+zW7LhF4qiyHIm7z/5u8oBF
Ku+8qDRS4xToY99EYt3EQEMktmV5kq2J1EiEszqyZoLTcJZo7/1r+IlEpT2Dd2D7
EWH+XvxTuIBiEHFI6X+Sr6SIFq2qzJc8dRmBY6wQ8borc8Udio1rag1JZERD9p0x
nEWO/FmWIVGtV5h/yBHgwlGP0x3jDTOLJVI35mS00J1NLI8mxLNggD6ZzlDzfv9b
GVq4AEfzov6d6XNsa+JxybqkpgWSQGv5TdP0GEVJZoacrirDDNkPPzu/GJwwJOkH
10WwuM6kyU/twhsFS/9Asiwgu4UMW3y77th4MGKqmpNv/pBQDYfySf+T2bjesJXh
4nccBKgU4WEUFE6NHhS+rya57G9SmgfktddCS7CiOsRubYdRb6mX/ZjI5snOARsJ
sNqir9XlKK3YLXsx3GN83PiuhDaqLiCd6G/Z7U/fS1r8LhBc5gGZGuzwJcHqC423
UyK1ielIYKIKFdUfUIs3ilIJwMv3+6TMM8+m2CH4dvz/BoGaN33UiOWRo48WuCul
ddcnZsMz4YxlYTOTj4OWQlBj4v26Zlb1tcP9BigjeA267l8u6A2mKalxsUmwBeL5
rhKPVeS4Ne8BWzm4txQ+Cy6y43QZOF0ms1kMrW8uCzNfhB/CJNIC6r/zBCVtyZZI
4PZWxphajlVrWDNyxNPOAgekSNV2WHwLkmhyBbTT5Pi5MvvGJ1GBJUeBkkWEz3nr
qOIoGIRuumki6N+p2cAS52Z+tSaZSElGeyKI0boBJh0KEWyNcR8imV76FttBjIMH
u8JDXNSI/EdBUv89c899DWnhpJHJepCd/irR10JIWey3KKkJkIwydgw755C3lH1A
1TT+fgALd2GdiDyu0g3c2FjvxvZjTnkgWC1yGQtWgds70MUi4dK5+Zr42N7ZnYiD
RkFXJm9PNLL4T3SOiNHt0xqVuUqlDqB+VqNHmusiLtHYRIkG75FwgQLpDJisatlD
oBSUARcS5GwxWfpBp4AiFw3gDayrGBBSaI11w/t0gczFrIUvVaXGBwHXToz2Y3iI
arU8kh9xWII2Tjw1Ia7QOrJSDfWyLNBmBJ7UqOWTzQ9ayTyekIS5FyO7BzHn2jWK
hZMhKDpXDb21tLHAiPpywq4iIzP3nlsRiMyaTyxrFPs8YAyZfFBFcBYknJn8WSQD
A7mtgnDW+UdJXtSHY36OU9ZqXPIFVWU91ETKrne2lN8HroxUhnm5kyhatX8wj+Lq
8sqPW7Vl8HQyopaUKi2Riu9160+ZSLVjgFUHAogQYNfRp4RiEm+9Bm46PwMck0/r
4ss7ApKL1JWZ40kq8rtupqyXpvjUVAmGPTyivIeT6iOFlv3UgDTPsJC7tdPaOqZh
/8BhvI7x07eqwsoBVBNuhYacm83zgvqgAsNOS9O53WYmUrEONmTUUDkSc3zjxFAU
N3+qE7hCv/9q6EavfdIC5fV0vuDAEHTiXPCDk30Hh2fAelmiaKGiL/QLyR2ro7v0
M58js5i7/+crIRG1QZzsVyjxostmw0qbeekr3vFqPECTTVQC8TrrzMLQyeC7v1iE
wknqHWjTxaVdvOPifNkA7E0r7hnX9BzGlqeA2fTIeICV9EWLTb112yIfMPBk5+7n
+wVvptp1D/09cizpI5zI3XgE6OfopJR68W2Tmn3j6fSNlwpORMRqoOkfXfJ2i9+N
S1TTvaYKbnLwpj9RnuQy0dkR1nK6LTZ0+lbzkQ83GUn0IMDAmoRG395KgyFG8XED
vjzQ2PHNb4e81mLjaQWHMVMAS5UZQ5sUGwYVdpBgPnAqfiy/p5yExRdvt9ra34rX
ozcgRMHfsI4K7kG615h3t5dtuUWmlyR5+rzvFG1GJAhQJeRiTpNr0xHGLuGgxAWI
i9LlSCeZZoEZEMx9oQHHstmGVIKEsP/F5Q6angEYR3t1kIF/yEf3rIpnny+jW3i+
asWtuXo/LYhmCppRojuhWYeDJrFG0E6TJ/S0mIrXax9YS3SBuLdz63eqUH2B5BIh
`protect END_PROTECTED
