`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KGTljZfnFv6INHiF24b/d5pSb9pwhvwe5sMvt8pFjG5slUjVAlmFBMLSr72FSRkb
/Ni9sfdh3Btmj3hlgH3lfKUicK0C4EfCSgIyC2M04YsH/SZ4qZjss0bmRVCPZGQC
oezTJjMCyEzfsw+sbj2iKJrVxF9CHkech6lGYc8opNINKAU9NjZrVNBE6YsFjOzd
Z5aVfROijNDefidK+xHVptzzYYOjaIXFywJ8ZQgOi/murK+PNvEgAach+uxRoJcA
o9W+7E0WIHZZHljDln9ICEBlhzgitl5Dpoyo91UcJMk3ZwxCl+b0DzrsNBtGCLXq
dAg0lhxvoZet2yFApwO+mCYu2DIMIMoKFJGylCdLJOwYbzo2zlKdMAxVwyb2nWqP
27C4zFpCF6jW7j9WrYtb8A1gRis7+3eiCBBv8SMIeds8i/ZuqK8trrthtvhelhas
NrF/ZrnyZVWiW6MHWWde8Vdjm1YFWBRXGeOFQKAozdZ3syRazPk5ITPXgpXmwj8o
EBtu8Zn1uTZsNMYMPn4jb/gqcZIAxNhZIRbxBORCdb4DeF0N8QsEBzynq+Tx1SHz
DgzPygfLRlzpDCAPoCHU9spjwQZ/A3f8LGoIwsgbisEIJbS7oTolW/9ZSw31IH75
E0ylOmheEiHtJ4yPkyzxOwqujgL8dZDzVletgcvZAHO2G2e9l/HB4pK8jIYe8GSA
iYcicq5t0x0oJBi8s4pg7l1u+Lv8vENUF22hVGSEbiDsrwBKGZ3F1+soTVDeBd8g
I/YFns1L1RA6jNK6emfx8VZL6FEuoRLEptmsZ2PL55Z57BtT5sLFv798eLy+Mc5Q
x9P0ES4z1I1xoCgNYviT3p4ptlM9k4JkALiTy+uY/nedrHs2gGZa0FnR+v/t2Wi5
vxIsEqIZrv3lmLj+Xh6T0cF80HpQESe9ecS1ANjqqbJOoeegpb2sfe+ooovH8K9y
eSHqzKD0hide5g+5wRzuUyrUqzxX8R1agrWTTP2lYglYABlOtmqYE6W2WRh8NT42
z92uqz8tHV3YVGhvrONnuuaWGIuDP2bwgW9BjT9/X8NrZ+LcCXxqZ6gQ1QP5z/B0
44YzymDHf5mSaUg/J49fpY7yKVwiOtJjL45nD3XHfogO+oyJsqME4v7jRfA/O7AU
5ndHytVYngVcaB3dWmSjFqbOCrVZIYZ+kxCULN+b0w/8p2CmgXKrxLxk9b7FM0su
bfDftQ2fn7CxuAFodIEjlMNU/jBNy6RXi2eGKR7ZtCZos4EngKKb8z2BjW953kT6
vtZeWCFdhHA/7KT1OAFfubZ248eUuCVeOAI7RIV6M9cMaiYrqINXZhBPQhx/Bh5I
0pbabj+3wFw2rLjslZvpbnnoVHCQ18eoG792j5uJLdHPJ3u/NihTSh3q4ToS0qGC
qxqfAPkNRLBkQ0x02ODR46GmwvkaygNYDRZnFluIJBWu4NOHG/BqpaUS8VHwY1om
xxS8BTTsmNU+HHBMRw6oPxtGvcpKun36LgDfF1P1933zKocp7KtTln63r1v3pcPn
F8AFcz4qAR6nnY5EKRqmGkgA1cHMnp527vJO2qh77+zFvi8ygQiMRi8i8febtJeC
e7+l1pUpSp+tqQmUrdUB/Rx+tsUFZSjN8MDvBW9ffp1kaoooda+lYvWcFoAdexTu
sAO+nCjZDe6frTFxFfnxXC2f0wND1VbM4FwT38LHL9or77d9ljKDIpc5jlEtVGVl
SceyRGYh/GsOW1CiuMSluTbaU0QuhYPkYZNbRLcrBpYB324bOti/udWiZLZ2ux9D
qCXnq1G9J1p79o0THG0+rFP+RHX9Fre3zDH4xuzDwJGjb3BE/sJ3xz3OiohI5rey
K45SJTXkvUmKfrLO8MlrV3KQnQVNvirgls4XwdG2RozOz7UTPvWjhv/KwtLL3Upo
igvEKMgG48dHENYoTe7/f1fDU7aPE4ZZJKIvMFnRyQzdl82+WAUtjZTSoCU+bp6P
TcXBfTt5MZYTmso5zHVpz1gUiLYveGMsEHHN5GqwIeDPulQQmGJ1ll62ql/oepey
KKKejOR9+5GYACdYxDt87UigT9qyt7KGxboUveuLvAAObj89HRFt9iWfKfsfi4Tl
wOrs6EhKWmXE8qtNZlDUJDsnfEw915gMphqPL5pox5V0d6MD2Fb1P0uWyIWUjMgE
ZMm6udx5QgRNCWUOR6kaXs4y7qxmDWZCESgGSHDbIfUzcxH5+ma0XYY7XQEwDYXM
Mfzb8QFaky+JhOwEiNFhMfHMHpNT38/If+fkyN0fmqbIoHD8cwIDGQJmNnhqJ0Q+
FFU+fybKhthy5gT9GDZZfevRB7yZhFw4b1NsaGgHl536QEgSpAq55l+F/Odpp2Zb
zW0mhm7i24v69fnAn9p2pOZrTvDz6g+bZy6BSYt0sDVbVg+/k/Ujqm4LXGrsqbv6
LbS2TDxp2fogF5QbHnWGz5zNPVaEp5Y7ZDDwOE0gGlDCKp9hyHI/qKc77IjqNNmJ
ItQmdVWS6jKzpkjCJL1Q/gLevrXwzvj3KBhCvTr7nYRBibf2rlDuw8oVhSHroyNx
PivNQ4gkOcKrfPexyQvbEgzZBWn1c5sMUzi6K93ARit+MKKrH4677+oBGNaSB++d
tG0HwbJ7qlG1c23fZQj7oc9D3iG6d0/Pv3gS/AiYDuXbuWuobswGYMpZAHtuxwvl
6V0vfoYAWqrHi/72Kv4gD8StzGNXvzOiul1pNWr0Edr+90drdttinH0DjWU4iYah
dzSQAii+vIgg4dk9NrhfiOAFp5OsvAI312wCsKJVzKY33bewMD1ji9iHO6piSa/h
gl23OOZpZiiryRCqtg6JRSOtLGFpdwEJw+u1mmcJHO+Zx1WY6FarsCysYuT4OpO5
efgZw1VcXw74Cg9U+3vI2ZD++cUCVgq6Z/ZXNXu32HAlqWoEf9bSpC55As2PE4zn
LPnCXy4SizsaQJjNCD8sRfuO01d/MKU0cyBOO7TABBU9wZuNGbRB902XM2bUxN3V
PttZyPeNrFVtkOcxHEkKcxaIPmtU7ZBfjfIT1KZ+ToOlynlbYU9BKHKLT8J+tq0Q
mi7xOMb1I2GW/WpOZYrjhlPLWKzufWzyM0wDDhslHyvFwSMclVF0B5wv8fq7LhTM
+FffZ7WUkJXWbL3l/eI/yHGwh5QmVQB2e+yefb+gx1n5XM0NLjPucpxkvXL+ssMr
EKdqlhCE1rM01Nah3le0Mq/EN+9HjycYlkUsBP1DSl32uMDfq4onGKRjJaffmUCV
bGMavJasaq4iTLHbFf8wol4NtyvQUOBoYY1tkEHxyTAk+/f+ogD8s6b9boOytiQL
XACCEJryR8D6RoUFMSDNxI3oYiL+BkAkJ2cnE1gujnQ4jdo8SpJ0/hfcaJA4RY82
Y7tgio7g8PZaqg3wRXEWhTUWAcxcFQJnMV4HpAn4/nswjXSFuszKZm5ArM4NjUrX
HNQSEZBPB+37EedSSXyn1Baznt0oRWCLwSHknT4JgDfGIP2Z+EH8p0SqRo2jBZDE
ejMDJzNNtKejJFYftQ/pK1aOn6CpfIvOzujGQcHgYqr4BDhm+S8euMdyhA7watGw
tLUIMdO4s/Li5Br1q7u9biZdjBVhXQTHP68fCCrd3YTGrv5Kg/TiBrMaryBOCqPD
ZvVlga921bD3YgA7VGjlgIB6kFp7H8INX5QupSeXho+3xOP8wFCfWJffguQtWRuI
Gf1e6UDhr/0/1SB4v2sSmDwuMvtqvjonAeHO2+Exa2gd27tilnp4tdnKqhC7Atx9
pXJl1sQEwzX16pLrPsjxqYpKkNfZ8m62PZbz3uHmnSvy+Hz/KiqzO5ncLcjQOjZP
zpXDO6+94FqZcZYoHSenY92JOlALKSU0zpXuPYvibshNVcq46SObU3VRf4PFBC4i
zIJfYVUlo8iQmBOZPUuDA9xiqzG1+COnAsxHbkjhoFNM8v2q/WGgAR2bSe7XrdWG
k55N4X7yVRqUiG8CZaJzk2xA8rpYaItIvpu7Vjm491mURmLBdPnmRTPleKTqqEUs
b6fXh2Wh1745hkLGfK5tj019h1FUNQnbNISdUEZ0Ewvi2lxHarAUt+11Qu94YWe1
b47uPjcWwvZFlkHtozarH3+buWBjnSxGyxKXXJjeDAjWJFG+dwrItLNWiWEtBq+z
psNUQxpsZ46l2tOOjJ1hcdDgbk7yGLZg1/Pu66pDQjHwF5SQTq713YGz0wDcJrmp
s+iNXZOGNcAI1fpAQxpz0Sb8f+qt6YivAO1r8m1F4wCQwX8/4WmeiiXy46EqEK5G
OXq8WtGZMhlygqbqMaDImfUTzDUSxlY2m0CA2HafBIBvRUH/RpB26MxH1efOYDnA
rufo1NOzsI6+Wj799WdhO/B+txxIw6eDnTi+jtoTEM0NxUnr6cDRSq/rwiHPy0aa
3TqrViqoJwmmM+qUd8J3ldk0JJHCixUNLkvK8QRJ2a4fHBP8xQquviOsYCMWs80d
S33DqBYhVKZiGGJ6m2mTjsFak/Ptv/9YVssWle5NbCxnQSDpwrW3sLh0qS7OmgSi
YYZ05IsZp/EV/5Bp2W5FZOZeAoDsD3lDdhURtp05YsXAWORzqDoLsx+pTXemmAfv
gVGWB0Tx5aVEdIboyx/S5TfpG01NBJ7gBBVjT/+n4uatE6GBZvCNG4MGTFAZCCUb
nXxjkCeY0xV+1hAqXkNkGmbMffHNlbhh0NCuBTBbQyCMzy9bhF/99pQXwNGbEYol
oDe2iXpN1ghPEjqhEX2FZv2OSGtXQIowmWdfrlc8e+npeQdIkdkrb8TYu/6ESN3e
5069FhwPkn9vfnGuQIUp1A8zSwW/YQqrmEbjGXx4jcqGx+dXtgF59IuEWB0OhiDB
WaSo/uSzTRr2DX0ys/Ij8apA392oDgcZO+1uxd5eNw/WJpX3PsXOw61EDRgVMX/S
+KPcArvn379+PpXmzjmFBGHfyjdsaxvjqWTtRxoUYwtadgBmN82qEHzCY8ZSVBbh
RVPYtZxK6FH3wkeaXFIo5Dtn7PCjs4cD+UXd6jv6ab++1DyhxkMQXZTrehz6GzcZ
ba/+4NQ6BE6Y8NhiWaX7OOsfZtW3y/T3UcVq9bd5cA4jtgHlH8NtEuOhkxqtAhaS
kX7QVFWxY6iZfr6naMUX5/Or/QK9ypyFKHZWnt1MZuzOuP/g8e1ngvI6F3qEBBZn
rg9UviiG0Jnq754WHZ/r/pZIfK5i+6Sk1jUC/ziDFKSx9L0qdLb8sV7tXp/meBJz
8aVNs2nfiFPSzkQ6rthRQV1lcTkaEbZHXmcUzkB8xtomEvTvupJmT2dnsoEiyXh+
CTn56e5cYv3vV91EOExUfntAOHVJmoQG/NfdcfIDerOltqMqoWhd2K8sl6ZgpByW
ec9RrpvsKczfOJIuoPquDVQo17j9CE9CDxLYJ7F8/TUQYgR0XGpWnZWzY8HYJRrC
zldDHrvspifSEVLtf7SV2nIHnscMzAZGBYhgkamZZAltijPkL5Y+w334OcXahsyg
ZwjLc7bQon66vN/a0Vm4NYyQxDzcdXlkUcbXQHJYs5mr1RrTl+6SGTLM3LXbYgh4
WIhZLPiZVzg0igv3KYISJm3a8ml7VqTiGNR/e2yiYBBpvYnr12xXaSU+qabIvMR2
Y+GSv0s2Z1nDSCYO3Limq3QFfYc0uoYhmS1WdycMMAj9Gbij73Y8YiqBGaz/dr3d
0tFDp+umFeVyfHh7d41xixImRUhcS6SwSsE4LOAQsjU9BTanqQ9KzqzNnoz2/suh
/8q4fjRt6GV5/KL7P3vj9Wm+3huG6pzjaveGzzX3zlPuR54aD50yGfzricYezNw1
rkbL0Ua7QvTXZzCZB04V2W4SN1pcymQ0KvE2OhRQMhlbiHZn5/XjAMMb372i2FxG
UPkf0UEJsjb5vqTi6Ce4sijxmmN76LX/19zwXMBzO21DPdXT81SUsxZ0bhKb5xx1
h76z6/PK8jseUsbZLPhQl+8o4wqwY8TArM9nWyfSpPSG70Hwxp/lA9cKHl8JhLOw
zah1lv7Yj7xNZZyu8cu3xIknMxj+tZWyFntVsxPXweEjXl4vDOB9oGqGf1pI0BOz
ahlFA0Xsn2ZM31MJYTdUGGqnw3sFpTouS/znu6hXPNViXAzzDlfRvxtHSMdtwunQ
Zl9EC1S6JLCSOPykwgKkHuDErmV/w5myK8ASPBOxwTsimVHbHjxnO5wESjNnx19P
wVM1GumzBu7DxQkuYGv4QbmFwYO7BcpqofzmQBHRYgfbZ8kzOr3bnTvwy12KYYNr
DmlMqpAsflAeUjIqfODHLCO2h/WmcYC1QDJqAFqHUZrI5+78ENc8O9mEbXSlhHsN
gS7sj9R1vmPrydwH1gkNQaHGqQvVmcFkjrUtEP8i6WF9cQmEnNX4xGjOlMn+VMww
neqpEwtXDtvqTpWogIUnw5oQYvYm1xqkszfpYHB2nMMqLyzPv92CxpT1IiovJZpe
m57jfqLtsUe9FSsjnGRx+ZfIolHn4o+eDRFdhNeiCwVi676KYb/8ScWGPEknCu5W
rkTdO1EQAlhpw9EOMnTNBBXpGMY91HUo/PEEFmYnnee1s6IeyPUmvllo6kQtFFN3
bRYhFu3MuHtQv27O0vWfP4ZqR4OFqni/dXr3JCdyt4PDXescnZQRQHtmx1d4fgqT
NSmgPKFvC/aVFmyCMSv/Ce/jdDBQarC2/HhpdDBUSmNUEk7uVEuww0BfvMmX4xxZ
87maB9bPmI1ZIBws2cT75BnhsFsVH85hLPea1Y/HeIQzlA2xhG17lHBEZ4udt0o7
mSvDbfOOKbDYO6Ki6mq+ZQ+O8hjo8KcyUvCBn5FpRlSi9vgQvm72xWibXPmUF3YC
O06UXmxS49TMnnvyewLGSqtMOgpd3hdKFzokjNfQXIpBykiWI29Q384VeC5CAbeV
TI3kEYzgWYLGbd8Fzymu8ytADXZ74FEg5cfjAv84x0yLDo/WzE3PJQESnIwjeVqj
G69xDyDkYKWrqM+833yDrJPRmYUBGF8A3uZbGnnZ/aGe6ZYGXlOt0JGJ4BtmIQvn
qDsiRmlRN7xRkxYKdkdbHiYeXrCTcNtniKkryhXA5BppEDj1/wRfLQiU6sGobZvb
XEW/4qN4sVsPaixXGc3G5r2ctEAnvHxWfFV1ZuJDr0Qx9JykqdJz7NMh3cQyF+pA
vsCMl5gKTVYjeB3KCUdYWtgJcHKJDfq97LtkrABhTs/Acs0o0CG9nArL27xfmfcr
e387bJXPMCGWZv5wUOk7kwq8n0HLvgOm3vLZE1k/+G5nn316YWgekyf5jpGVKB47
i4PAjWr1AnqAqdGNqkm4jXxFHeEMNSvfaxd3RfpbAH2tDORbwC1FUqImTy36Rpj8
TqrCqRCfZb6VjheWTH6hnKIaqCCCugYJUmILscS2+obXMZIO8dA9q5t9+/y5L+S3
T83snezihLX5UlPfHROVyLQcC6kvGSICC5285LYbGiyx7XojqhscXfLHD9ivbc9t
kiLte1UJsvptoPB00FV3cL5pazIuy52tU17kr4Eb2cHPFhSw5HG3mDsWQJ4f7yB6
VtJ6gDgETxZDPFmHBRzWhBNmA1BLDk29P1tud+JfvqPPooXLxXYezUxGU1Tp5FLf
BaIaKyoLbzc4pAL8iNUK86r+xoih95WKNt5HwXX+RwIknmY3ZKhqxtTw3TASBgBs
RLgG5CD1WPR47mOfXc1Ce49tuX9UHlVMcpQ3m1DFbjmP28iK0l/hPcNP1BtiilEm
dkSBphDvuBvlNFizNo36VyNUkTKsDpXL0v7aPQPnzGdEaAS64jb/urejVJTn1bNm
gvpuMsL/n6KcwoqB2mpC8wkf+3wlQA06KY1L97wokOPKIeCx1Cya0uKKgn88VKgA
0i7GvXh9cG1kxXw5+7e9EZxO8nZQX0uoEV6Wp3ezIMg8mXaRiEtkUBqoyEMOaehd
ZELwms81bNkUAO+ukgp3r/0+aFIQH2YpEhOfYwKRNfJBPuFC5WMo7LvVVHJCm2oY
CmHI+L0CxOwHXE/mDwMyijLpljMZbYKyh71nJ4XWyvG2vhtlF8LKREWOkdgLnTkR
1o+VSdO8jpLDSwTR9VSSlJf7H26VVGBfi7W9q4kjJWwRo1bYLq3ObhiTizvO+FU0
KjInhM5AFz0HjCFYmCUt6gnrhfqGDNyqEVKS0gzOHNAROVfnmgpZZYFr3LPqOoXv
FWl9mfzoLtPs4Ib77MJXC1XGO/6KsS8QHslSa9WMX2wtZPGzKGimEhXfagTJvhBz
yzl/zlZoRqjrS56AIcXlzdVWwN73nhN9CahgSJXTsj+C15j4yYb5X3K29gnZrWOI
rLZmA2xLgziJnvScSidh8ihvjZmCMVj6YX4zkc+Kpf5ZuqoXvR5ycsOUYInD69DK
nJx42+9u99zvcICU86jmTF773+tFOkDvOCEcIj00S0vUwCg1ISNTW011O9SuTl8P
u8S8RZxonmssGMpUTovdgn03sEgJqgL3nLNWtFV05ol59bFZKu0dDl5ciuScrDja
7SUgOzT6b/KMy2gzgWwgnTRsZHa76nDwJfCn0IxEKkTMPMDs3SR5cr2seYv+FlkI
oKnW7ON2biRycGMJeAxe1l67w090HLtjl1hgpPOWhFMTQeiJ9T6iHoEkWwJZaZ/7
ezhBJY9YsXWLxjONBjvC66OngHnBxcbwmLMF6XqKSQKYnfQ3rUr4ylJcBY0jxY4g
LWqMzRQ43XLHFmKM/s1dC5Jq48A7A/mhc4NDKWW+ndU/nzlG7etGUm2pJfkDxnfp
qLc0fJJN690gs4odwF7k2a+2ew//fu/xwxmjBjTfwqAnfbHQ1mjYOglFLRKdsfpv
7BaQUOSYIVVmpZg9pqL5wpteD5/wNH6kDeRSx4vD2dSyXn1iyYnPDApY/RNfB0uQ
thUWTCv7O8QFHxNpynaLChmPBBxvcHjSycxBhhSZNTx4UCofulKLulSOCBbBXIfU
+erO7nYf+4JqcniysixveKiCberqTxRepjeb6p8mlawn2R0tS1dz9/O+PkAOCBRT
8riP0ROLPjjXhkRJPmonxIr1upNPqB8O2P39oLVElx2fQDRkNIu2K4vxaI1OwyGH
PGIbhFMJamnC9qFWgdkrF/BjzG8JGl0JF/qjeM7GJukQrRDmqxJrE1qmFZ7GKBWB
k7hcf/7EW8R8Tmyw+vOKZlgLkCbgbVMwzcLcmLDp2sTE5qqvGWo29TYtAajCZ0hu
M1PlKRcPYEjAOljjH9o9z7mJvVMHhFqr8wJqPOt9aSxrq1TJiOAcuSBK+zXHQAx1
JXyiH5nvFgoxfqDRw6aUqQdItGmftzIZcUP4Z8rh2QEFgQiGD8GYJxlBKvKvSeoW
CXrmlAA8wUEtqt51Vy+l5ToeLSV8xiA+mgdJiqK/ps11ZKDI1OkZ2iDKBSSDQki+
gCww/pCcafVu3o1oM9jyW5oRbh7BRMluzWtMahwa8NcPkd24IsY3d5cNr8gpgLNU
KOdIcZ2MNyLgDzwxzwvjTq+JJfV6SfzH0Jpk3DrSC8AS2l27/mDbeP8x0+pXsAy3
c0kVgJDMi2tI5yIVcKgUySkuNrxl/iw2qc9bE2tgWtAIGQsgYt9bNVqWsVtMuvsm
m/b3qM97HmespJ152KqM6m7p6DMw53uyCaKlWi66M8Rg4czs7PWj+FVxVWIvtc2u
8QmEDL71GSbCEn6CFGoZSG7W9ZZYhvHU3J65i8AcUnnL+DhqIjg59WSciSV012Xo
ntmRnzyuzSlQ5zxf/Y8ZcxQFtfQr/4dRfr1xEx0zRCzRjtT2UNxEpLpFYsMqutbu
6Lw0VLKmiefwc7n9YToQOzTQ6Ax/g9dVBfq9adu4vj0/RLGohfCjjVx0HYOLI7Lm
qIHlpDLwoex+Ac3EI0os891L/FwMs0Yw2it+2dwegKadVK9WabhZpNIu9xnx395q
WwMPB3hLH1Z48q5ZaTUR5jJvGhVOAtxZczLIgTtboRt2yR9zLubLcb0agzLg3713
so+jSqBUz6yB2eXZKXQx04ISysO6D6QFXKgXMkWLQbo992WE/OM+uDe98H3YdJga
3qjBE7bs2hm/ywNPtFHMTd35aA3q2n7vsZ8eY5M9p6nietOCW5EzX1DTC7K/n2RB
rm1jLinHfOiTZkEDWcZPms6mOOa8hMdUzyc4xgeZMMoZ3A1uF71KWc9u+3RUVadc
Ql5uUK1exvcsxujSnvo1rHlMq1blQpwCggiY/ftTrewjsaYD91uvC92Kc9iBmLKp
fkCETeFxUGurGh7yN4vuF9lkhBUrPynkVOKb/kczwrrE5E+TPkNgBueFmad0tT+h
z0MwtWMgxocNesZ4avJ4lbPqb0zdbOAwaLw/xeXOqH+y4HFTZAYlOmAsuukako2w
yB+sRf+g39ODzJf9xipgcIq6TelAaeamicGGf6j0amD3l0wUb7rljEai99H77gf+
dK2LFLHkXOvbeL1VuzbCz97+YwSqo02GBurOa513FqvCw8H+rf9K6u95592q4H4Z
BlqXI603XTyBrxF0nMKBlP+l5ChgAqw0Akq/G47ztrEGRaX4VKI9KqtKVivGHIH1
GvKbvL/52E6qU9l9ltBoxj98FagE/+gPBxhCehqaYkhDcPYm30Tdw4HwkTGWUGrB
PkXu/ATW/aSLft8igDLiq8J/Zj36hwI0g8Mv1nY1uMUA/dXYI/+35VhKX0VYpir8
dtIiKjCK2CB9xcrz67qI2u++hZQ3VHRgKYs6JdrC+ZQDD8sR3tfXR5gJgDlrMqfG
oBlSJ6gnkG4yB0p2+muFswamQ+HBbmRV/h6f0BUH0a4vtgTHyFFB4MosQv3Qz+5v
mTNupLm/Xw8ciJpVpR7XET4ZxYMYk95wDGUX61lG0C6tDamtWVv2lDaRMSMcTXt4
MphLvTEchmng3XHo2hOpOYPeNz59JpEAkTqnecspDlGATaqdAS+f0sEqLj3KV9QZ
+XpaykwbW+ovZ4SYLM0vqcWzzt5pUk5E61OKVMMU2eagX45NkfenvaOF3UAlC09F
YIA5VIkwYlZWTffvcLVQmUAOPVqF3NJcaMkuWd8iqKah5Ee9RHeQJntzqsIZgDPg
yTETUYhWMRtM/1Qg+nC+yRC/eiRMsOUqx5SKQKVmr2EdXwEzgu0lICLZNB6ipNEX
HxfrJqF/5ozzPT+If0eSCxwlykKe1VfT9AATJ3aYCX9YiBUiZvK5jfkGYf/GylZt
6GXmbaTOxJlmSRP3wsGpf/zIGgsR02hW+7J86C2DoRyj88AfAGY+OkPOUvOvskXV
3PducuZhOsYC934N21bUK2tYStJLm4BPm+MMHXOxerbf2Kx+SiSTMqbR0hth6gdf
ksAyQt4wmai517684A0IW1oARlpLQmV7AFLehWUFQ5aJlP/nhI5IPnAh7mKBMeZf
kr9NOrpFc93oIav5EjYxJBO9ovM4h+nl7et6co2rnyh6syfSVY+HFlootvtN+xQ0
iGgBeQg2+PupsE5fbzjyaHctJjDEvwDyju4NUZP69Z33pSQLFjLl/sYBiDvcJ20u
UmjGRTfNFaSIAwQs0O+nVoqRn7lF4NjUSypyoFEy93bocK17lmB5vaqz5X8irkzM
BFuj0mV097d17zMQGCw44NjVkizZgm3Mcobl88CXrQn/1Y+VojcxNhCTk4LN0eNo
g54otNo+/X/HOsWAp3p7JSL/rlj2G6qZSTegIfbpCHmXKNDMZgfGR6AmIJ+JJE75
ypJtwLeNPVXDoE/KfczEsHTDn4RkoTmR7qxSurtIO4reeOPZl84lKV8+pLxRing9
Ml+Mo0xqFXFQQeJoFDsmiB45ILB10VbHumjPkGRwSBwmMeBSux43Hg8wG3XbxuQI
mA8fRB1OgyabFNrcmwGZ7DPCotOPykZ/LcPYFjvdJQkHvOoN2dSHC9VPVDbiEC9q
MI/gtT9in0rJfD6Ig2dKb5hw1/j4QaVLWatGwOPYSz89xbjYjipkWH0ZaAOmAPIz
HdIFUKJMjsPqEeDYqRnTz0Z8E1rWeAUXJ2cXjlScKzVIl/s/X5OKPMj9TzmmtyVW
OpJ5UXAfVQd3gZIzfR7ji35utcYrVckcGoUEgOuxx8zN+VRREiGs31SIVh4RaCNF
3MwxyCI8OgVx1noBsigT9zD+eatEAdx+z8g1i7Tz/9dAOX5T5cp2YPj0EBlPo5Xm
MOXpuweka3/uIQA9B+TUUt/oeRiBqn+xqS/ObRDZ38YH23ULjsvatc9qIS+Vsw6I
x4RNvj0cOB4R1vRYp59EKKJtWzUlEFZXyjqFOcKe6p5gvW1zd5SH50bhpZxCmgtL
GLrFRrnJIO/VmMLE3wAYgbevlPzWARK9AAHG9p2af9PXI3AzFRSWbqTidfBK8JFr
xiwje1FISibhRU1SP33IyTgp0tBxRncQS5/DjnSgml7zfFKxKWe1IrrpZArOGj/E
49KxrRLgahyAjQb3XlP8AG+vXGMoy0lZr02r0Uo/QTh9tcsDdetJxRrLR9tf2qx+
Oon8mqfa+aJtXMZa32p2mmIlICCFo6P9V8U1Txrie7DQY5hV8pnaRJnPOULkO1Lm
5uPsNzkNM8YjFJMUL3tDVuQ53ykR8Rg9Hqz6bLlO6t/sdjBMqVzO+Py3FxNRfnbP
6ey6mZOe8poV/dxputeIZMo4IvLIrfqgRh4TkJPh8IKvSrWnXH5vn7ilYDvyg+gn
tuASqN2xLn8Kveukka8DimlQeAoIC0ZF0Onj03Yt5jW4tjy3nyCwbjm6KZxagxI4
puK4mNxJsf0f0aSkxsXw3CZ9W5gqOgLuUqUCKdHuY0rCdygnc+8297IF2T+g0PBt
82IrC3U8bvdG7C7GYpp28FVIR0Q1fWJOvSkgu8EiLXfkKq40PT5rnlbwGMhk0D6F
KR9Sf6yu6KNbZjcsIXn+usixJXCC6my71WDT0xQ7YGXSQ0DnEbSgkYAeYU7aLTtS
zOjgOADxKzUReCd4pso7D13qm5czgj9ncZLVlj5qXgKgp0oBpKEfzjwmPBQuIDaw
Dx+T/Lfnwcv90k4SBA8RznT10AahezOw/UXO5nRE7BtkQUJgSrs8b1CZdBrja5rj
HR6LHpq82khrqYOub9RGtbkz3Kpo3fVcjgpdhYHdtvRXyPzy9sp9zj2h/9Dfl1u0
79xZlMonF3bwpNfc6YYeGCsRKpCz1P8o1VEEjFYDJu+0pTGSz4Ghsvvuj8LQ8xI+
QcGcQmjCZ4KrWr1aKBMZrSzYETyf1G5OAdL2CkbJKP8OkEN0S/5tvBwSngIBuJFI
ctvNFmZ46lcs+Hv+Krg6UKjT1NJEvgqvIyO+xSaxQackoey91JxIoPM67R/LprDQ
MdGCwf1vqWLen6pIhI2xFZ08+vtwKwJdtN5VxHIDEYco65o8ieW1LLxWk/nbmWgU
PXmUplMq9FjoaTi1/EKTU/vWkwgS2V5QYAySutuAC4jRgJlEMDmJNOtv5jDL4rOF
LAVHl0FbvQDetXJGw1S4LTMd+8aM4AWtsbk3sAe97Brfc8y/2uiwmgh9KWi3wBjO
E3tlUaeJw6MPBHntVeIPmoVutHE6cu/tHe7tm3XjArbnUFlF6mFD4BWp/AVpSMKH
m/UTzXlf5KtiMKkewPRvOusDbHITuRvz2ecUTJCh9F0auyYUMgoBLZKgYNi1HCd/
ROEWjhcmlFTlhLXwq2vBrToAclrrHf6OrSEVJ+oi9uHhEfAoZkI7PY/Y8+7qj0V5
glaDKTXMuB8OhQNeUs4QeoXs3NpsgWbRmyNrCxdWj06uc8hT7Fo5OJHdbja9tFS+
m3t0R74G2tyL55bJTTGsNodv64qfdIHWP4EBx/EK72aLUzOs9ROpgyn9KsusRZR7
wMMu1+j5I0m78NOCrUDFqIrF1EJ9nwJi/1XC9I7FEMo+l9f5/55vJIhvInnM0pRI
ljKxD3yXiKh72/vOtxtIrLVYZCcvdjxxqT4FHk0QqsrB/Zn5hWJtnZ8uxotJT2w7
U9rmOLkEVpQy2XE7Aj7JM/e7NtaLDDp01GTQwt4SbuTDiYwjEsw/xKQjQ8w5bUqD
mWSOrWr715nDnBzqJbZ4j+PXDbhhIN3lWddovTwKSraM4HCMzQgOaoGjOsP6yNoH
xbgEBuuRqrHqWLXLlRy+h0RCm82MB8EHsZ9h2erDCPDq/igeYaMhgAs8oT36uCRx
/Ov7yQbjxQ8kyPUXvEY8mNykjGdpzoYeEc/6WecPtoL5hQTffb9sxpQQQcrh/5wE
gC4uiQHL+Beblfsu3YLqeDP4mjKfcNS0SaNHsfUkL+13TQnSgml2ysGj2y5QeZ+n
6l4Pav9TkDtjdIrTOObwfCwioz13ynK86SOFnIofZuvF3lydg6LILHnDfXZMpa9i
C0blInv+EwQGQvM9EbsF8Yv+a34EtEM4TjJpWGRhf9EAV1EPxxYc3ajvIcCx5O21
IBYvyStemK/sNnWSRdxv7rSfSIgH41SGe5tNXSjqiKbkNTWsid9vhMqa9wLMtgHp
gqT0AzhBPFJ5CsK45EyZsmXrsY77dhjJ3irfWIgRkaoLelQAZGfnCgg6iN24q/Jg
HTRhNx0g3in2xWibpmf10/q6ZucCKD7Hn0+vNZrN6k6X5VdP7DcU544HyCfAJbwb
ReeHLTj9hjtTQqMhpdxy2TJzziBicTB/N933BRSyFmJQgkapIyW5c9WMPcNdv8Mm
YkwzSyvZ5q98MGALiD9O4wsv4zbYta6BBtGcjVUAnDwR708UT5I5AwdWEuY7SY3A
jcJ4rm5Q+4iXNuEpqt5n73QwblNFwblZzgnOEi/3jJeSdlfaoxLUd86foB2uMkYr
7REWwuvfuwmV2u55Toy+R/mDcCDjPHF/jonITvRAmF7ywZ/rw2iR+EPUOHXnOyyz
zSKod0NeB9xWnZytp4P6UVKFL5zfw/wZ8xL+d1zefRqzwjgb5mEEf/eirmMsThxK
51RnuXkZ5BV8m92uLmXyqyThXYSlBIGQ+gVhphrdNDyvTY+eqXun8ufE7lBDluQ6
/QP08toWz5lkeheKASFzlz0XXiiqlB9ABbz8G7m7S2dOsCKf2mwg9Rj7Pnbub+lY
FWmuKw+gxpO/hglqAAM89eO2VXqra+7KsIOBlfUnPc8Xp+ddb6g0vDwNuKgDwmRP
/5dvFhlx25SoaF2XhAFzoIhEBm56hW25kff7cigDfPf8JnLiUc8hfNv2h3fVMece
EgzJo5/aZYDX3jEM+bYyNFS1EZ4l0f48ZyqQ6+LnJ1PUOad0NSqFwp8OxH8060+Z
B9mxXAu/qNciYFXhtms+cNYveGXPKoPBuXA7ZeIlJZeCsjLi502nq+zxHGWX1ciX
kJLWOT+9HMJ1N1mVqO3nzmm8x/6PNtQg9Lfhn34cebLgF1DzOJlm6lGZV0zdOk7u
nkkDn4rJaqpifl+vfPr3WxDUqLVbJ869p3vG++L5aHX2GtSmmeKcMd5/GH1/rPKH
EXN0bsnepZpSNu2JjGq2e/SprpX1yF76e/WhOKO2ai3hEs4SPnJV7PazNkynCchm
bnJPfN7Mz4gDNt3rcLPs4s7aLzfuldfk4U5W/upVlAp1m05wPnh9VC4g4EYB+2i2
FNv5fDMdLN+e+mVPsBfcnfTKi3Zu9sr484qkLxtkv+NhIhLG9VE4lasVdVNl+Dso
ngiqk9R8olRGMAc1QQo7RdSAoNvu4P0OeYfHOZ3flizTSY02LZh+3L7uSgsX+h7Y
WyetQ8yApjsWtt2cgSAXVuPjcYqY8DJ4j5FAL8lRUK4lTIDxQ5jtShO/GevCMyGf
5NufBPd6LwnZWh8GqJWkXjFP9Kqypx/xs8QRm3nKLHXdrGv1x+XAnB4U60zMliG1
Jqr8FGF8695wa7dEedcbis+cdC7jKTfure7wijcUiIpN3e8XjmSDbCX7tpm6SmBh
o+x0+qAjumdyZwY4W4wlK85EO9o5w/yLGEzpRk4aJmszWCnOW5CSXmF8KslVAjDG
UK2Fav1A2o4sr7xxlv4YzS7sBPhBwcL+iuWF4Jf2UU8+lKWRBvCEa5MU+Adr/Mt5
dmAgslO2QkjluYms9VN07tqNmBysOin/bakOigQllp2by5lRoo+WoD8XbgpjtD4B
zfiaj3jnTRIxp4ZxfJskf9PA5of18ypZyJrGcelHdTQqFtbDtQ4xSJx5iRUTB/Qp
PY9wt+APE57Wv3zzuKgWszxuTnXhpqaXeoZj16X7C4qamFRsCj1wdNSq1RwigD1w
0qawZZGRWVNP5S6W5Nbr/2uN6Og0dgMHK0TukjvSeWoUZyznu0EbBMooR3uNZmw4
Wx2YPXZNTHWzEPPnFcLMbBQ+JwT+wt9N7sqqwhEEDSupaMyDRE5LfGYEAyT7AxFa
mhoMUes0nJ6T6ylpUgd70tAZ+Zp9EJ5Rkx7AdSB1NuVhayYXmPFZtwMI1AnjVv7P
INCy4QC6QcL6n4XueKkt3bJyQ3EAQ4EbMw7sREE14qM/cvqgaTAXoxFQQUbeBuNF
XGet+PuiKm5w4MGlewuan7YwCVHcA64i8dbNk95cByFNKWwhNV+aTsHzhwWCgDxO
vTMH7NDhNgJM/7T4NKtPTgXEAjSkvlqS2Hu7VQhJr+9lmLXkrkyZRcGjJLhuX3Y1
w5hwAqB6OE1NPQdrmMNjB40TMwA6uLqfyXjhqwfQhQ94GJrrIROPb0fy3XM9TVb4
aLxK3T5TdqlKzbVXt231eLPL/FzolbwTq14nYzuCzMF+B8qMLzRCH8TFUItuUEBV
Ln4f59ZNcFdaX6NBRqd9bDPSbxlqFbk1UEEX0zmvt2SE0ZC42f4rDeQPoNsUzmG0
CVxgszfM37yJDEAxvQq4fJn26KL7e46+eGeg67pSI2kmt4AMt8MCRpq4IjIZzze+
Ey4lPCt5DQN2qKLzxUFNORDS/gD/fBtJlSslNeYFOgQzaScdvOlviPiawcfNKPgr
rv0OMj5//3FQywnnSdDuYLvAfgcrlXzNF7adsyi6c4+0VRRZRJdUDrCXC1X1N80m
prUOfkRkxQihlkuJtdEpsXczoqGLUEV2UBak0++cLG3S+O6txTd4I1VV0C34abWD
/saVZCR57SqSuFJ3jNK9LDifipQIXxAw6cTJPaH3wf9h+IxUpT7D+0oD0mtZXmoe
ljC6FvHVoeKGojnDIjnWipJ9h114FjMw5cTGFdCowsskZA4twea6dyxmbFSjsjJu
qHcH42KNFNUWPQ5wCrQa5JgaoZUsoapwpm5xA7316ioBdf2IMhK34o0cQHOjnoW+
O9ReNVwZcAFEjcOsmy9IQUWobKYqMCyolEuD/ymnDJQlzPkQscmqieiIQh96POY+
c2+RSoPAe4oYDyS9ZinmW8wmZrKZNvG8UK5AtwgoemcZ+IrPejn5xJgwSe+ljFru
rfPU39f0D/QzV8NLRhay+GEyS/KCI3SW+s2HqLaDTPaowij0a3yChxHSzP+oXFPV
lV6h/kswjuareUI3kR9u3KJNTOgr4oO4Wfz+JhV5ZfalTW3M7cg38eWO8/KgF0Gj
x8O8v7wJZNFkfM3JJyDZ9InAa/J6RiZvXfeu6g7xrwd503wl6ijKpSUAkJo3FYZs
7At4CY7wKmFthnuup6edtPy/4yZEiHt84jQuwE237pzLaTsPKEuEv9nxTbMzykMC
vSMLTFA29LJCfriV2JFoayaPZHGePo5TSRbbMZNv0rL39sVVfLMXgRz8YaskzjSL
9EEE907cqoJhXlSEv0jiQCpmxxaxkA7AArUgz1IbHHU+AyLT+dUKq5bBdG2i22MU
aFrmd19IJUfJp0GkPRFOi5G5I2u6WkuHXg2wgYOhP/RKxjgDqFZQv5Hi5J6Xv8zh
ijboVX3/s149lOl2IapB8FVUxXKP41X/8qKW2ZtxrzB/faM2EIB3U5bZHtm1Eudh
Lg0Sv9o3NwHut+riCNdWburfp+y5GWnoluUN1Z3gryfdmbcWnfo/NlNZIGq4yaWv
kOAyhVogPbivVHy46ATE4WURAXPunY3e0UAybi1CwXFRDUa0BhDuHuQJvb2uA+lM
vmw6b/KuE/PJMMBGyBk3B6+d0DFTfG/CNbbNz9WoKt6I9L8co9hUwEkXTsJW6Lyd
jraX4DrENuGpOfv7pR4hiEIC63RbXAl/55ZCChChzwaA9CN92Zo6ra9zpzCIYAyx
ah9PUmYFtq+ON3lPZd4QtZNFNaF3GmfOLfC1WhbbNWFU4E2vgWcKiYsMGmI1RegL
dHsKeUr412TVqgol82a/tCqWTRXrwRTraIj9ezieRV95M5QDvfjLCmXzT6+AHhi6
j0G31H5IlmRUFX17Tto//tiA7OssWmNtOCO19S/Hh/MMDpQ2AlbI/ndNBacWVHMz
M/ebSVHc88Vm/exJHJ2DxtG6KNqOD0SU7HE86iT96V1X/ClEKuBcqMeklxE4vEOT
eebozZcOj5HjBPkAOJQGfxaAP3ppWlKoZFs5NFLCfDVFlMRFjz3pXufyQdTFbC82
y6hlPdUdlKGeOellUzev+MGaDsLpmfwKCL4JGhUtPoSmU2QP+WA+exzDpC7bclkc
B+yV/KLDuVyOoGsYvdGYtDooX8bvvsGhwo+TD/A/g7p7KhL74j9DJCpCQyXFhRsY
282WOHmGrGaXHoOiSgfsm9lKilrVoI2dCHgyIEalzgT3W3JApC1dL57tdXRL2bzs
NjlEpGeSzAkUPzvwvqsOOfbqG9EvhaakryafDSI4OqvwQqvd7WYN9Gbkfwz9+zBd
GIAZbvyGtSvibgfzEIlO3skm5Zlhxgl4x1+KYcEr6RH8pZ2UueIOyG3KsMCfJVPT
4YeQW9UAM/Ds4e8WyhYJ8X+B8r4xwRUiTcmoacCJd78v+0vk7FwG6UkgxDfWWudk
kQeRsaxFygfqfEGpgG3Fj754MNmDLZedVBT15uIO0s9oHRtMZOg35JowpQeoDnAc
OBvZBUoFmxgQn/gIN1Y3AM1HJftKWjHZdYR9USi93kbloYeSAKgSzDbtSAadyF/q
vpXAE0QG51WDwaAnhe6t3R81Wdl62SYi5jmXUz0qZpcVhS57rvBbktnvhoOk0abs
uaG01cFuH1O1ke+uMXCeXY+uIsn5QxNfzAOJoDzLuJG8sYBKW7EkHfam/OjKEgar
9gt2mXsR5QuHcnRoZMAXaTdk72Z/5UoptIyfQTd68HvLboNTOIDUyMd2qLuTMMnV
IT8Am5Lz1Y0PdGTeof5S7lWf8wIsoHiW8H3zGmv7gLF+KIL7lolL/veCneiJCmXt
O+ACtCcVrJyaitL4rOowx56istk6SJ3aSQYwApU4aOQJja1PopKHU1vuBqh795YF
4/RjY+7ZL098a9mwCx3C9aDRRo0Eni06zqcuQis08CMlR9cmPWRl/4WnGj5agmUS
Zw6NTIdzfbm3iDdin9X0U63y3Q9UKdnT/WoqyxmbGgJR2kenyPxfcee5MoiI6vcG
rlqhfl2tnZ+30GXuPGCOgcD+Uv8liQGb9gDp7f8suyWyjFccqGyhbNJqSU7iRiXo
IOctobG1aCfGxw/v/Fs+aL3fKTXz5diGN1sMDJZhRYLGck+kCinSU1BTtquvnGJ9
ct/zdqdXeCgXfl8VP7HzRHjwuzO8LaXtkZPGcQt7l0SHp23MDyPA1QnM1117uPSa
7cPtIujDRz+gbesRk+p/+AMhZK1yFBAvb7LaqpRVzYHTXDvq+fYEfvS1fx8c/vV0
jC7Fk4VpsdDI5iwL1eoQeyCJQ1r3a9UgZoWnGnrfW/y3otfhPEVjTZLg8cvUYWkL
Vl/dkYpZ+wwHVvR67H0apbyezDFDrtAPiKd9tGnXsYGzzQ/kiwbflYKMHJTxQaVY
yS4WoZXKfykkinZKW/cq7KjYw3tW4Uyhbyw52oubwnsTejfdGp3ig+YUM1Lb0Odm
nTwnpy3iXrIAseLi6ORTqrm56cGhXbRQfHk8Pp6RGXQIW995ZvzLJx8zRf01fZCp
M1fhDANy5cnuK/kVtRjhxFFOubdVrSRYQx09C+cK+6uZzq3hDQrwpwYocoLOZk4X
TvHMo+J5r9wp58rgV5rN6o6U7uVC/mnEz+A0J4BQ8btDGYg4ML6gb5kHiP/LuMLT
UwpGxzA2HpFpMPDljujzDAGni0VkpC+1hkMDeQz7NxAfzkwQJE1X8fp6SeYLgGAF
0l63quwGZqLnzLifXcvuypqOCmoBvQsNXLnG/jkr8LCSDa/nkPv90h44kWlsq3KO
Sl527mP1AlgMwBzSru2Bz6jfwvRo+oYNRC9I4/n3Y3262k6Q5LsNblSrIXHn5uCX
4cUksEaX6a2Q83/9yy20gFmDh2q7U57oOYipb4cN9XJdjnVCyv6Ie7h1VjfzOuxI
lIvLShycsjxLLd0Hg7KKL4bEoFByW/qZdGM0r1CVCz+uaskKozY5EBdZir9GkZVu
1cwCAV8iHvZp1AYLu7iN6Z9k92r74cX00fKUkM7ZzPf11r/qxj/Uq0G+yJu5ZtIy
64aP2PY/hjUYIkeBqi4nStPqorfZuSd/Dk535C8/mNVLfR2Sm5M7AIaIMK7QOpSC
iQB6rz+RTWCjljvZMQ8DWNlMUN2MXcDzbTGBefsb2ckOAVOzuKvX9CrHFGG6JDbt
4SkphOOV7NoUisuDcTGJVVmAUoJmgqdrMPQFwKAANeFJ5pFgHTka/dYA9jYfitlo
5TzpKk3r3sT963C0JQCW3t3sYguCRqkQKCHzKuZQY3pPAJKQtGpBwf1AZF9PQSmW
I58JATMbIt3pPWmGQBLEIoBURPE29E8483+8AvRFxVxgNrk9KDaHrTYdV1Qj9qk9
bJTRUEffd24ZLFQ30Ug7gZwUedXTWOVhf8I0sZBGYoMMhMViVUnO6kaalgmBLeyP
f0l3WhXf0CBCzHHPZf7cfAQlx2TJnJzxzvZIb1wNIRDfg777kW5DxI6QfgwtCGkg
YtqcEjr4h6wu/gzBBl7K60S1XaJg87UL0oFC2hbi2tNMyVeCwvnx3M2xud/kix36
4lwCL6RX2bDYBp3Tukt0rZE7B9LD3qNAVlSZqT+j3tFf1eb2ZBLfGVc0BaeY1RGd
JA/80JorQPVjizzvwbOOurjN+aViddolzx4jjulEaepOfva5xDPnFkySnbmU6oGe
psDXT0KtiSF5NAZkMtZMeKtws0Qa66l/gpHw5xA3T89KTJhlkrzYoJ9RULtBY1TJ
sk23r3hXlWLWbiZaTEepcFdvA+LXHmQww1yvi8T4iHG9Vb+L6C8mX5hk6lhyWd+y
oAK58MgiBq6nz/LDIbQsI8sFQMd/q7lJIbUY2PPN9mKqBaHBLwviY+nFu2i4qnt1
lwURV1Bp+n0M3hlU9V3RLn8FTkxXBkfsjhxlkXiVzOt8IeKviRTOVd+GiKOuVZU7
I8Mcv2o9Y+zZqn6FuLV4DupcamgfcejD7+3cZeeSasqYszFW7h7AbHwcghMN/EjB
0/8OHOo1A0bda2sIIXvjcAyOhZJTy9Ou81KCJISf3zac4THHRvvdWk8m+zRRp5U9
G6lEQzhPfOvE+CdcvVC12sfCy/4C8CLazTd81CntoCs7CMAfF+uBBU4HE8qc3l/I
Q6ZTWUxlVSvlH1No2PKmInEXYST72HGnj47frsb8VFM3vNYniolCLiFq1w2rw7/H
pz91/z1aE1307Vw6ILAu3lHMlIuzGQzfvZY9T9r8Cs4lfP8Dkx+zfPWyQsEKlZ4X
KGrtninor0ac3XhrTLLQEOk05YRhK1lMkxfQ/GjL1T+KvoeHFgjWeukNhmANMyFJ
TPJE+r+L4EouyTJL1GjdjqNS/kCAyLmHrIRDwRB64Wbw7nHyNlafTJwlvZViYoNF
mqlV6D9mXfl5eVxenCjpm0/lIofzaYNR03Qb+nNTWXMQpYlucYFmIL9cm+bBib+1
xGmRtladfmskKulAES/qCWW4aTKnPesYRYbFSP+jC5YJe/RDDGZImRX2yxCl1u8n
oRCJc8PLMqm5ncr/38muPNtSzeiiPwbIjT3LiNabwO8hQzhkigmBA/m94SvySLny
Ky1iDbJw+uhzyGTZaE7rCSFynEun1HtZuvSepdLCIhlkQRfh2p+IsbID4B07dUsS
37GOLR+5ncDqRl7bhKtzKT1P5WV3VZaqkXnRH1m5jWUAE/81nPvlb+eiYFwTeRjs
8inJ6SUm7eT14CzzTjSw+54g/djgdUQA5ekuRXNNgpsj9Gu1G7ki9PmjTVoMnVed
3ztvRKQJV9EQjbgL3BUUcCbDr2aamJqMLxiwal4yHFBu0VK4sKf8luUkS6Pavixc
9bE/e1jzivOozHnzzPslOfWt7fAKiu9IZo7gSu+c+qlU+4LP+SODO7JfvqGdKl2C
5aTzNMO0Ry+XGgJoLrXU+0UiMwSmJvgM0601Q1x89aJ68SI6EI/kYrM5KVUcnwJ2
jv2KeyR6cTu6KGmYu7FBAjitW9w4cH6IFC1AJ20/au2Eerw25qQZIwYrkPUX4o8i
uG+Yi9ls5EprmDDkVSvyoW/qxyVdmHiPtTk+cJoqDrlB0pkMPmRbJnox51z4qG2d
D7m1M89nF17fBEALUrfa57bTjuHE6J68aSdSC0Sp4sNTuTAqee88ec8Uzrb2qbuB
D95CNYUz96Qm9wNDeX+5RSDu87SYxao1a1EgynBubV2RAGNJn9oIrtorsXEFu/lE
EH0CelxGzZqESXXFLaWVfP+PpNiKoaKB/HNF0CQR68O2jNg/taNoKHZTM/hkdFqn
lNcLAnQRXKIeaaSgK/gqP/7ibB4nshf3d6rp9fiSW5hdynpFXENXnBbyyp62MyV7
c/ForfMbouzxFiY7nX2ekfLjiY/7h3xOrMn12qBiTjCeb7OGc++k6/K2iuVu5wVP
5gCy3Juv2EGH2Lo8phS7LnyDTQzKvF38dQEF4s2LaopJk/iTWxJXPKuGmrgz/098
bhzMTYO6fpA0bud8ZWIAw1apexTZErDO2w+TZSYwyOGHzzFSrMZOrljz7CbNaJhJ
eSeB5p5FHa6WJ7oTSHOnM0T36NhNQiT/56dohytnBgbPAJPOgwZvt/UWmOJ5L4Qo
kkbgMxXzLk7QEvvC9VskqnfvY4BjYFswYsHkrD5GT5sbw1kNLrO2d05s+Q8EQ5qh
Nmi8Lkf3o2MaN1V7yJE59auRORBb+WXXcqISTsEpwz80PJUnKKmEzYIE9IClS1Ap
qNdc1NuiSOskdCZ+IhHdg9iRTw3mAGedwnzNY6yGA9TrlEu3tuyOcH3cD2ZvEAB8
AzBmOgybzs1Ghl0Rh6UOky4bZd2o7An7OYnUkHRQkCTKn4TLKDg07P54R6bVwTlT
/VPnYf5y263BqPpkKnyEHb+c3S5bqKcUotBMPVAUlnN/7H3Is30dcqWBIgXpN4yU
URfMEugK7/Deo8c9XXVv1z634svkUFGG2e6rBcUVPL7mgMWaDuYld459ZfArQ9Lw
6HwNL963j/zj9sQmgVys3TRl+L7iC0XV96rw6LN2gdGhJ7bbV7Ycn0KLOwsP5okv
4Ppmw5e94YO4uUOhFAhs6u5AII3+kpz/eWKC+a9MkuWTSXPi7zdAmkcrFjIw2vrJ
H7Lz8Iem1Sr/GKHRq4BjREdF3QDD/2NTMG+3ojE0kGudyK2sKg0Ts15y9sWRGAmX
aT0nW4Z1kS+ObhXDqtvIhH3GD+LXois8D79yeqz4lL1jN8xkdlSH7etUy2TeFjKJ
hoJyKxryKbCTuPaYbPAccibvHtz/s8Tcb/xkh8/MX6S915RxiKkyEycRbQ/AZhJh
/VkfDpIp05fpa2LwLPcUkTCZq4mIxjTBaVMvoLdqYk5DGpWvVFV35nr02CPJuGNI
hRQiIp62BjVqHi7QAuWLOBHWKlBF7945IZ1BVmTPMX7Tm5PZxj5Qmq604jCltyXH
TrkoeR5qVFwMcVQKGNFg54G7jhANPhBHi4mtFpEM8Ov/abD8Od6BkwzWk/EPjqnh
f3/k/rpudZUF9ozA/BXz5NNUIlacR3HLXClbykSVxZLBxs5sT638ZA/xvAIXD+YL
H6IyIDGsZb2UfSiid3kViS4vTdUj7VM+ktBfqOyL+7uYilQCN72SxJv76rSbbxAL
3qw/82br9kCXNREBqykW9aygTIAqsi/WIFzg89M1BLlnr6sbLvD1+TC+wSehURR4
nnizUdoMRCQFjH/rJGXiLqYbSSQVoMK7ZJjgbXS9cB105WYRjiGNWXPWNUcdkTrS
RMwaNfDlS1X7W3uA7mHtBjqMoY86CbvX+tL5N4+vWzLZ8IgUlemmZkCG7dMGL/ym
jCFSsyPwnMhF1NuL5UXATsF72pHxkdDFdcPsiOnCvMk8/HtpT8f+9CnqDbIfuGGj
6rPuYrGPA8M7cm8c1AJjpp6iUSa9BWWdy0WxMSDaFxJCL9Xwgra/aTCK8fX5U0p/
WtfHk7NjmVwEipS3Dad5LyWpY2MzPCP819WnKa8ZSJM1McOO4kKTebGnpE+UhibF
PypaybfVm/36Ew4yMu2G6fJPvKRGtgB8SxTBx8cOMmkNZDvqn7opo1zTlk8JhQDg
zZ2mMM03Dz6Rqt1CiijN7JdLZhzpHD8zhCeoayVbN0t2dAtTXLHZ5yko+Qki9BOH
NvmZNtWJ4AqesD5vDDZ5vjCv8Hb1HTdarEK3uz28VCNRXHHbrtpBfbzZhP9K3HL+
q1abk0ApznnVvVFwkzn73rdOge/iUHeQ5ZwkOvuMuDo45fNxOkKxiPYlp8j/iVUY
71h+NPl68P2LCjDz2yX24In/5//+ir+TgthXBKppBtG62ocDstybjVZcW/m/KC+u
MFYdHUbMjuGYWOMAmrs4KJ4N3fA6dV0SHj2RJyfvrPEhsmY9AwvLG4HYPU/vLHYt
OArZW4JMFltKX8et0mYzAjyuMqi1/7TBl3Rweh4ND8QspTash2fGn7AGTpNirVPt
RCffT62I/NluU56TCd1Bw6qwE5ABA/aHH7qbhjL9gYfHxPjxNjDt/9tg+j74p0A9
Y6AKJynUkN4fjxRIh5+g77++6AjU0NIWQs3rUUtI234U/f7ajLbY4WzqnH7vIXs3
aXy3ReOzlhLOWqI0N6BSqi1iyNHASUfKJq0TXldae/zl1PwnTUyhVo8N8rsbEV1s
HeCFhsog+uUtgbT4ttiaH1q7IO+tc2a1a0k1or9BlZ/rjTLikNpNTHiOs403J63J
Ee0o+4ykkH+32IaRy6kUPvcvMBvHo59CVuKoPykqDnUEsfgpdwBquPJWL/Al5e7n
CZ5Y3bi7aB2YaggElIH9XGpgawpc+ysOBYW/SEDHs6ad/jRhj3toMPxLffE7JyXv
ejzjXmQItqJuPr/ZptTFSlVAm6kImConx7MfR3GvgwAAqIlrFkTSDYeJBDyFNSw2
QYtV+adVyloZI5lyMhXmlvD1yAEpGsg6hwUESgtWE/d6dOMfGZn6cTQu07oBENnn
fB1qTuX9akkLzycVoNvHDI0d8Hjr9sobNWgdm6yP2ahqIqv1ySZX8u5QHRiAc5nT
D7TQrgwjkLMVWB3ckFaCT87aY5+K7utZrNu33pgBynTvaxLhyDvqjmDKC2eZqCBY
/4Bpb6ghmMerkwO/LY4QNEcOJaevX7pmpoYWtTMlh635207hhPWeM6PwLpt5JUT+
94sPi+B0qHOd2Bl5uWozaNCP4cA75ba03zjELSXy+QqZgSgqR4Mw+Y9Q35Vim6yT
jsq2CdYnKjvBtcT0gGy2NERFb7dIP7GyoWHfPG5/GJ/TjUjEM0KNzgQRWhcMszBa
WMGpxW/iMQO0a6rni0GpUWHIv62UJmD+Sr7djg7p5X11dE/g9fSCjV8CDgwZ59o4
cTzjj+KhBC/OZd56fye3k+sR5hUbpOqgVQIAEV25VG/DtEe06DsSHlnQeS0HCVYi
THoxJ5p9iD3Lruh7Zn2HwvGMwTyLYfRyeDpSR7NDtxA/IXfHesk/renHq1XH1uqC
FoVsCOewkxg6AYfngKgLlOzjbSVSz0fFtCw6WlMMwGLFHUNsR1tj2+MNobHhgw9O
1iO9bYLE+MhHgyB1/WtKQBdR+WUXHL1DyH/v0geC747Jw/bTM9460iNCs67U1/it
HXHrJ/eRQ9GnB7zfTmTm6vIZF1s5KrAJeglVzvIl5WMvR1a6y04TngSo8q06aUAw
EKpH7ivj4f7gOrW0mavJg5Yt5jHjUonM1uINAirh/fM7qsC9cpnt+UBj494tdrF2
jK9KAm+kaaB+PKypK25/DmYF0qe6s27f4XJaOgkCAF2Jd4zqRlE2bQyb/GdOElol
ymsihM/krDZGP5T+3C7IlVjJSbJhBYBcwwDWJQhgGcSn8ixhGtrXyDc3sizBBK7o
FsABiO03x1o8I8UhSF2Wzy06rZDdsEAydiJaPnGiK3iN0q3ooVECsuGY4pyICIoi
XJFVEmFh4mBPLCwz60QOQVvLb5DnmbWPn8pfQ+qjqCIckOk3blQsfGLDUquPZ4w4
eZ2PcuWJrjISxPCo24Og/mO3nmL6n5oBOenGZtL2CtF5B29OVvJQiOeHkgewNt+D
o7a3GimhO5Q9XHUsa0GvZyoC1Zaa/mo/mlwTwnUU8JJXi8UxxyPPATmpI7pgv7i8
vaLUHw4LRoxk6Sf1JIeMOFvoZb3oxFa/6Ld05QJ0cwtzO/JmnLOdKnYzXKSmdhK8
3NJT+fQb5+3AXbkizFyBIs3zY4xUxsIZTm6BGeTvZR2GG1LLeAlPwsm4Kr+7w1IQ
vENYeNxJYZ+mvnBHtTXXfRufienzrViGLM7QYB5gIquIWrTNx+T8yXdYojV4El21
IHbqb1jMcSBuwpr16itvKvh2oblPMhvV2wOtbVArF8WswsUTOGs3oyusY5jBWN1D
da+9z1HDFYnWSzfHIT8mLy4GhJF6eR88U12MEoFeVt/ZXQlWAd7WeNdaEQ5fRZFA
7SHEACXqfS7+2bB/+qzBjylorFKFC89BrKgtBaTPRJToXyiMqipV0uc+yXjVSNh6
U/6WqFHig8Rg/7QyoxbUz5meRazxGAA3ebLt8a7ja6EFc509YdjGtQOa6uIuTNJ5
JiXb4ibo0ne3w3Fnd0Aa4/ow0Tz0MgVNykqqViYLmwnHw8F3KWZGFqm1EdzDfgrr
HvWBwAdybV3jRYE5iPwv3DP4h4yC34twpjEF1B73ljHa7zIVeEWJQ0c+epWq/jcL
xaecszN20f550cKlKtl0wa2g/QBiuFq0ZA/7wQOlpBUPtwdGjbWiZs7tj26DvDSV
VJMxX+hgorEs8VKVqrs9AdP1U5RbnY1lUs40Aq54SA/qqbw1RwRviQ1wzBrJxcJ0
FvoQxee7IqTw6rZs/QFRyFj45zTa+laeJNo8cqyODQBUFxyhmKnl5LZlw6wV2AZo
cN71Bp3wq4qQldB+4LrwG8oxGSKAudLZeSGCHoNzdyOU4OXdUzDF3OmhbZk7Z5lR
9SxXJ2u4OYVCHJ+H9pBfw+naht2cuPAq0Lj6V12iiBYvMl3sJJ8hxAzFJSLru1uX
b4+FJgbBTp90Ayfmdp46HEzBxaH3sa97br67F4cOaZ+33otaQPNhXxQa2lV7TR7Y
na3zZ1g24nTX0vt9iVmZwogqaAQOANXdWn6ifbWJ6rmY3Pki+wy5pZAFsFeDZzSq
c4GgQKRXr/fQcsZGthsOOS8nul4oyxI7YIMk3phcstgHQEdP+rMIXZbCqR9s8Lgb
L8mRmmdk/DdGTs4Pa/rqsCbrIl23S9fmm6Y39j9suWGz0WSzmWeQ23MW5wV+EGsz
4zeXQxnPoh+rihITt1Mooj2geYYdjnZGvwqV47r7wm3AA+CjPtuXb316ewajGyP8
+nQODIt5uXIPjh32Zu5klYa5W+R4+g0gffuOU3Rj0o0iGthVfB59FsGNo28yAbf/
onkcpCHWCB2v19ZNAERSjRi0sUrf2tQLzCk7X9pYeESw3ctxhIC08KiVbqy3CVd+
+tMYv0dzVFDrih1mbtZuled0pQj4g88TlOwrhCIqyWRDPWWlX0atrGYm46IWaMTi
5UYHuqeaRy1yBhLEeLzCzDx5FLYBGC2lPGIl6RF20qEsErZFtc5ImjvaftY7AApF
O4Isq52ZygzxdB4CpeqISnqsz+iqsVEmyjB3/uymevMOF0T8oPkCNA0JgwSqMGD5
X7ESc63+PZmVb1vZC9IE0smGOZNqIFRd/9CO3cgWgq1Ek5+Cwr4nvFSPoc99I9YG
tTzMW5pCADUID5w+USU30I3smKYJ+eTfNCtch8guGoRQwFucSSeYcHtgJR+Y2E0n
dGQ1435+lswHI+E0S/dASHHvPFZpwjxdImERwuWHZIrugyd9s3UDrvcwymhqXhTf
a2h6Hrx81pcZLCdHaCPF8aY58mxMyGCSBdzn4bcELfGDDfiOn2uY0RYPl24b4Rld
FYDo5E2crpDqTmHWRVzJTnk5mig2oiMNpsilJdYBg6zBLObp9iBetvbEZttRRx3m
PyfDiOZTSLjiNSq7YyOiDpsMZO+1zNZyVC7NxI02q61FPoeJzv9uk58b8XR3NZ7M
o/Yazninw6vwKN8a4zffzXNOyHfT5xRaMwC6gWVrQBY7MQlwKNVR8FW/V3GpaCfm
+Kv9Io3a3bZmkBxJWXnd6uzpb68syR07ydeO4G6Q805QBCzvtiTC+N8EyjqPBTFM
0/7HpuSYxiJuXcIJydRPGQQMp1YLP7UC/aFKDO3eJo3Pu38t0G/wu1SSZB3N/G5B
ix4zlykONBP4+lmtd+R2rOjM8+vHp09UMPGRUwHkYnXHgUn51skpr9oapLYGWOqY
mLLJkD+1d5I6tktCuuebgtSOEXG4qRP38QtUNNoALGO9YpRUn5mRtLbxoFI9WHqP
t4DZ+S7jRFEvSHFyniLqVXmWCs+lZinaCYgP2Ahh7XpJR5dLJ9qGjj+3mhbG3yMT
10XZQrpgBC+ynqqrvLnISZeLQxKlxveS0C+KPeVfx0c5BePNc+ZtSPuZlNz6zrLN
zfmZZg+Cl+Wd3HnBGcW0Jnk+a7WK2ygS5nTbSgifQKEIPfyAwrgHbatTW7nEXGzr
/WasPXVCGidsBYr/+BKkfULTGjXe1GGhP2MLeRogOw77155ywGq0i2gYWwtjSRb6
PZh3ZHNw6M1Fd84fXeuifbrIsvqLpFsiN8MgJncqn0WtKeQP8wLIok4lrB8d8WlK
e3ygCB/mlE3ZfhTg9fOhz3l4AcwUpAFom2mWuwfDgxKNkbsEeDIgQxR0pMAM4vzv
PrxY+Z8l2MwVez3v9YIQPh+OuDxXhTXnCdXGrkOzhJD+0chEVj61onhc/BEqtzrL
LHc7tZB+GMI82AplCTplWkApJzkT5gOMtgQgz37WlR+by63gulYOOIJhpchjL1H6
1/lJKX3V5uoGss8bsRheM1XNWHUno+d9RYNSF04zwI38DZ2eCmtIag4pRDxqr9Ay
QjQ1iegxjAzX3uSDap7KMCJvmHv9q9w1euTftrwJh4RKBW0XgGsEergD6j677Du7
FCd3ABVuHne02VtBzwU71/PJJO2FlIVPGtxgVyLmtbPxxrjkDYhXLkP4JODs/12l
MU74tHOkQhv3oSVf7acI10TN/dHsC3FwC+36lT0hlm65Nphzfk/j3joK97nn/WTR
cr20a0GYgNSrE1ctBSd2QChZKepHHhlLmepjZNU1m5yQHtpO6yef6FQLT8uPJ6XH
PkNOiaRLM4zBpZ5WWt8eIXxNXe/2CmovV5wzINhR43QOub/pYp8hDvVUGHeCTxvn
BZU2b4vljd3JxKl9QBUH2x75HGca37ukaVyDatDh/I4du1FVCzhGTGp8nMk46Ttt
VGWt6jIVULGLdB5oFFub/cLQ28lAyIt8+G/Zj3V8kHfRXEoHIk8k/sfs054TZ94H
AE07lH8ZWRgEs/9SlyCmpdko489tM/FKfzoQ1ZY9UaVhiaTNq0v6QwlQ4Vghge5j
yOt3eAU9bNg/a+Bbvxfvoq8+2WOGG4Y6Jz3ilzJA7k0l4ey+pT7VZCNptgLrCqJr
95P2UNKuMVkvdH3GEG7RMckHdES6UG2eo1yIzz9zHVOTJPwdd7sJSGJP3SxrKIpb
ultmn81dD2EsU1lXmytL0NuFtHvSyFmwsZG4iNOsz7K05T8UPVVEWwKh2hVZcdaE
KOcdL5cqeawQzzRI9syqGCII+SJAcipSqk8DQgQiFsihAcKRYuLITUV1xUCi0Iqs
pQcyKOnX/Qdt3gIWh+tMYZQwv2F+vJ8CxZJML+zQP+aRCXaoUmihzfLdfCU+fZiE
eKDX8Te6UtdS7E5n8BiMf0uJT/nI0JHvshHI2unr/Xwx/Zr8werw7hs0Q571KKio
/h0k+V/IfVOPKvubOnjwcUWKHL/n7NM4R0PhNe0FumLZ1/hJ7JG54FgbNwrcBoGm
Tq+lPghKk0zn5znd3M234mnv1Z0fStUDDmTR02OAejYDFIKG3rM33lGdWeGS0eJ7
Rx8RAEz5n80pVSioXdbplBACwQmL0ymie9VoO+yKfRkgXKvbRJpz9sm9WJMquhA8
BRZJCVeA9QgBDU3Llm4AnFjSWENM6uXp7nmcQgOVrtVmV5pnkGALvyrZFFB8wBqs
8e5G5r8Ryou9KyYTuRwlYZ/9NYqpOHy8NgcoxNtRFC2VMXusKk16n97ZPfFuBCUb
XFGCtc63G/dFCtHkDPPil3RY184wJ+CPhjJB4UyQKKRZjGSPweUCoPDRtQVmuwDE
qFKdr1U+eMRzzWRDiSvqM/m9Xw3pSs2JW9XNu8h+259l/mpM9tWpHhsAuTxmEw4g
tiTY8Ynd656qSoj8ZCxQ2/nH0WtWkV97V3GrJyX6lHlZgVkrp8YZxBt242YfCmnN
fT0h7yDTgkReLsWgKBkDSLLbXsnNLDiIdf2c+WMw0KfXLIaeyKStUwWkBweN+4pQ
1OPwAb7EI8NtCG/yY1JiJa0eImepVXCP11vJAAoYZD2PJJIbxx3Ikh66De0H0K3y
5H8X/lZYLlnHc92TxFVWMv40FgAoj6+874AAKhCIyQduLTO9iXe+91qj+DwbUqPG
NHZPIscVoQxIalaYjkSbN5ZP7ofFIjQ6uZZ2XidqFCk58ApEmHG2fmbOiZ1SLawp
Yx2U1xqzkSELqoUf4/usLwBBDQyvJaU6zjvevd04O0lejJbn45DfmkrRDh3r9gGK
H6d3CVXbkwn9mXBzMrmweRrl5C9sEoYMGSITZolYaIMZztTBa6m8AQPxyUF2IZRw
6XIPzhsM9kcjHUnlqeJeS0iy/DxBgCJGHclwtJrHXF8vexwgEnpE7ASsreXkNNup
bC7x8/Q+nUz9KXTmTGr4ydgxUiQQzOk3dY0FWZ17PwmnvmMd1IEZD60McSrJy1Cj
7E0oyb1OCZKqC+YMI6O/AfGbdFKRc9SmdJTgS/YTGHXVctibVa1mUzVLr9nq+XAl
3kwzsw5u7rcbWQ773uFl1HoZrg7VN1RG58ixhyjOOWZtRFeWGWyEs4DuKLuU9rZA
6Jz1e9mdmhRU3loc64n/wQJaKqggqcFXGbBEQCaTOTHK2bggMdnkKFWTrmvaUZuz
x6dnQprwijtcMFOxTc1JR0zi2jou/VP6B2nq4/CL4SOuh4W4vKyzm8/2lkMrGYad
hkzXBtnx6E6cd5zPJGx1CRTpp4P1+SFWOaysbaNYeYl2AWBP6chBPReRTijwsmuB
XGlkhKCZBXgtdhKE93+AnIjw1NTzS/2Ar0M26encpzbgEzhQIZa9DDjkE/FgfOUe
sdc5pZqwui4QmGrXajHQXSG+mrXB0+hRx1aOpF9VV8Qyn1n51VXrvFGCPgAXV35m
2dgWRHqNoCOy1jk9SwCE19QqwwDKhBONwVPzwPJBYYSNVwRcpd+7TtyfmueWzyBm
MGq/7Df0NLmOhV539hV1MeCXitEbb4l63kKHOSpWzhSNye0zfvm09GsUDchUSGp7
3jWPNh6o/VY8OFDLPxh9sxPGLAeXyp7HYMGY5Cy//kEGX6jvakUfxW2hnVx1Tucr
ZwU77zx/fo6H7lFzYaVnpXuhxYXWvRoAib3QPKWGspOn/elBbCJyV1joGdYRAN1Q
LU9Lr3H2pYwPR+RqmoAemwyNaMUUnV3ykGZzppV5UzQ2d/8zUfWRSSIripT9B1HQ
w+5+7fJIJfVy2dEMuTFKwBI+e0CIAZfj70uz13sXxgN1ub3rwyU465eiSK38VTcI
a93XGNh03ZA0VfZtrghRuheL9av4VeQl7KmxyYAdSjCtRytl8GohtMwZXFUdajQW
PDpWH1fqUqXTf3nVDfd1KW8/do61hrvpX9SoeMmqi4VOlv942+sKOZmm54kPnxna
UchLGh5PgRF3x8ZZQRcnnVPWoOOBDQ4d4K3+BGJwFLJuL0TyXReRudtfDG5QEggN
9aXPfoMq4LiCG/o3WjCdFODxkZVpM7GoAx9+7K35FXZ65Ez27NdmHB8JS+4eNrWe
BuYIOl2VfdzQEc5YSpPnE3xbm84OiVqD+idZs3Lixlq27RRHFTWQ5F64mTURFMov
ltoDt8nSE6at7vfbQ03FHmyH/ysK02ootWO5S5Cb6qt/eOMFJHn5jmoQABlkBWfZ
3txcQvXEiebuXMSb5B30G4d5GI/CtN2F0qm440f9/MLn1gStlqdBbM+kHLidhXJY
Ex4nAqRSvZE/CjbQSPxX1Pc58/9g4JqKuZ75w2ni7QHr6XczpmKSI4dTGMK6kKZ0
vBUYGRQ/f5rN8X5dcLpme3kHH5Lyy5Qbxke4Ojp5O5gKptcBQcbx8w3xsyhFWgoo
OaPd4+/ZW1vcEkIWYIesd2H/D3D0m+EAXPJ4qJZU9xTIi0G5/P1Dm5ylHci4BrUj
BhRIX3X/bqNuVnOBnlUBJW49Cxh6YZqfo+p7gI+Zb9T0lPvWrOJH15biUPBtqltq
8Cq68sRfaH9SfNBTHTDs9EcdFu53+SBasRVllflG4KbU0sqzk9wa0hFG/P8FbiD1
/DWKiBpcAxuJzkReuT9Zjei6sZNouijoFJE8mvfU9ilo57r5oGHINAmAlwcgu06L
fNClRD5BXxq64CY/qsh/RXAG7fXuMEg71xyctYoIfM8a/JDOha2ffBqT7WvVvw7q
nepATAnYdeCwEuB/kUQJPVeJg2HTlLEitbC3MYARik0hlqbn5S/MOOoWip0ziA3V
7ntbC65OlWGg+7eeRxCz35X8ISe/cdbbjGIottmSeRr4x/mVrQlgkgLMrofqnxtn
7SMxF2+1uX0pc8XUvQTsdY2eTb4T5LZT/AKEUoxcJSuSyinFlFyCCylnDd29+WrB
UzmjiAhBJBIso6fZUcNu5KeGg4lFM3rLD3ubxYklBfbFH+IUZh27j+hIuF5re2Df
PKHBTsk8t4EDhHdPkduQ2/XJzS6MmM+IHfeJcXlFOGWK01jrd0X+beAxBYjXZWR1
Qc4D0hCI6pvhvW6wOe8XnGgcEGJMotu/BJwsRKMCcSqKq/DpqIWSPVc71p3aJJRZ
fk6vdzSEGhjDIZ05xtaDK1YOtn9DcG9p3ydMe6K8CT4dRGrYsPU0zvafOQQpzqAb
q5rEPtG8TzGc41PIfyOjphs5Mb0N4x+NL3wYBGua0JhK49K8MMFVhgAGZ6m2svYe
10nU1gc9Nr/AhTp182jG/lHvnHUg2lnDS7qKU29yhn0DDV5Od8nJ5yis2sgwhQL0
EI7wMvneIJjR3GTVUsYlx6IMiFy8VacOT83q2BD9Onj2pJhbqVNyOzI6mytvymWI
6pkG6yEITd3wESNwX9OG7oK8N36ZZbuY3GqUVj36QbJJJwD3ss9Tw6tZVckBb/GZ
8153p4WpUh6cFKodYRPbfWEx+NCtikxfmXRf8Wf4GPtAH5cz67VftDsfFyQ7Nm+P
wWg6s+tQ65D+kAtsUIIKjGF1yfrf+JRws/HfULdtdQ0XBnv88rmxWy2ylgK1opm5
1U8TkIGm/L8PLxHGkDVdJi3Dmr6tEIwAr4eP/xaFzPfUyswhlMmAKfFN7Elotrza
4qYiIpyAQrPhoLJVLX6HbmWGYR/UWn8q26hTrsSufSq5wcqFHb+Uq0jDwBnRp46A
mt6qGwnc4GvGqlubzB6pejWpS19grL2alueDUm3/Ug4TVrOA5EHtsUksr9IGbFS+
22jhxQ2zHY0gMtakKImfCoFZ46ZbUNw90/8GdPQ1NT3z9o8hiapH1j2XygXMY8NL
292pvcaMyYLzOLEiWtigyzBhvpsvMzVvcOmXrsGb6sRKYPpbWIcEWM1yhbuC2X6e
plHjkPMAtRRA6viG3ELEUiPW6I4RDgwJ+2BWhGdWKVqNgHkk3JwKd9/AOAqz2kAB
q36yram5uOngqYuYgQeHsVHfzZKt0Yuiy03z/hXZvhNwZKipZ9xiyjmie5GS+zah
aWKY9ffgNRrkOQI5acZC85R37Wkp6TKk6WsNoL2LkuDj0/UeO6l9cIU91KLu9zMn
ugQFKi96dnqHeZCjKciEzwPN+OYYOuVOS/HU7ORZYXyoX+nsUcCLwIEEzGK33mIr
OS+zgze6KOyUvxhojl3vc8td2KVfbZXEnwfjKHQfrBarDGf+DkjMRwSdYqc1XoCl
8HWPgynofhOY5ZTucajK6lod79ckirRNxDCibgjve3JH0/HMHD+5ZCWyBJkbP3Wt
HojYB3YFnHEPV9WDirHbZzkvH4cH4fKKdibsaFFbLH0TsKxo4pT1kgG86jONLfqW
q3enesTj/JLEiOZ4/2cDiei/xEXE72sRXQ0P2kBHU6pNc3Rnmgs/hFWU9aH5SaqG
qStzME3pWqgmkBmiS9epLMrAOMM+gEWJ2s3Ei82FBGE94jOKLzDvM1i3LWpDOmHU
rJ1LfExkbKKYAqAzb7UhKvmAjc9CIKqif2hchbO/mRjqctq36f3vBydMzeEMCLBA
wd67MbEDnW8DTgpRn+TavgG4IbwHLq/eXHHOwqA+eXSDp7tcWCE73N8n5cCpPoXz
OM/V5uT5xggst+BOXpEwi3A4tWU6cUJtSPvIh3ONGn5wuRqTzqcQl7qk+MwALab2
ABjAIU/Zm7aENueC4JqaWya/DVdf1h+jjtPJy903lP9AuNxYVbDZjmgI9Ot5F4bM
Rj7+sI+vBtd9FkxtZXnGglPeJyhyHG4+lnKsjFM3d2t6wCloEbl+CJtnQNlIgmHX
wTJAxujDcvki8pm5ykZSOFhQKCf42pHmW679fEukmAyKyZsvLm+2hh2tTYY63eGj
AKS2f9zkL8XsuloXvuNL9FFKIZVpFDe3oQzyK7NcPnNxdfps+ZGzs+0r3KfXze2X
Qku4dvFh3oCdPDIt1cI96Hsq5b+7PuNqoNDAZRolhec7OU63zIUfpf8kr6B7xcMG
c6VrGGfbggYBneVHkai+gglyj1zBE32Kqtv2MoMbvrR0l484Z1m3JRSFmRbK7X1n
1wjGd9o80d46Jw3hzkwz9emc8lV3NSjBzC6KUKZ5+n/3zcF5YzGsU1wCfzlrXLdI
w6MYpYpbLeh8R1wlkAC9+El86EEneJ3n6ONZ2yVU8I5JcWPgDHpuuOYykpbjgOBf
5dKKXxBOpBc4HEgE8RpO6qEyAk0a8dDrCSlYUsqfuQlcPaT5dHWolMLo8pOis1yO
oS70eyf8AKmgQMNhyuDfcEj92WFcA11Ic8a8F+YQ8R4S9vjZunnsI78ax/RA90fL
uoUFePmltstvkjyt/IJM/JYS5XZu0USfZ1EnbdaxF3OBakiNJ9ImxHGJGMaTnCkm
mAagTxEPdVbQGYu9g8uokYpPjlBGWSW4oPDco01BmEpl/g+PRP7IHB4sTMlWpHnt
/GhvwVrVz6pfuLtaZk9Q+QP3F94KcSUJxkfJhlaBhoujSrVVwby8lps9RZ9MTSPe
pUKDAPggPm+NYteiv2lqmV0wrLQy0MS2l3rgM7rCk9oVxGZVrG/e2Ruw5V0b7/Y5
JTKF0HpelYRyc7bE7Fb2ccvm/gvI9sJjLUEcXpXNkEyjsUle8ZxLAUabKFoj9MH3
9XkpeyztYCjojDD2NKbRfiAkhwsDL8CYdOiS1wKxx3hnPBnP/ZLUym4dBTfC6fG1
Auo1PNRXGE8Bi1zVhwm1XjdyKgvL5KY81dPgsbTzpHHngjRQNyesDwSL4bCw8DqA
JJec/AjcvgEG8vJFJmZYpGia3h1thTy8ZePd8qbm23MFemz9NyR1lVKtdrfBB2ex
FRJOk/pxF/d9SUoInL0Jv4u1YEHfT5qJ5et6o/uylJuERA5F1EMtxSfOX8SXGRRO
idpM0FMDFMl8p8s6Na2BNtryH6qX+Elcn7qBMGSB9wIBGNYUErrqt9Ylk4zjsZ0I
r8gG0uiao9kmlUbU8AuXKtO00UVzdw4ZAtRXHlShaBItMyyk5dHDdM5bekqXegAo
AfQad73e67COUmn3tyuOzUtpurr8SRlTasnRS0/wFUuAjgOJRESDHGjk1im7AnBG
/iXb5SP4xuifyyKhmUHQquG068i9mJPp/NONY4Udxui0sa5mKt+gTZy2Hh3+eLYA
2Kui8tnSN5Pl7AeSnjSF/tNBuupxlvwAcVkVQXfOxpw8bWka7sLPMKxb1e8AuPwY
TiNCvYL0zoT71uLEWDEL5xex3bt83Zd7vjTnxp2/wUl0+naRsed7dbCtU8WuViJK
ef4eR3n9yChg0f17+7TcifUXBwlUMlkYhzterkUVd2rwnCSvGA7HV5IBVGKkMATz
2b/IXqnR6ZAgzGatxiFoNHyQyDi4c1igz/cx0ETx6tOlgFk0MeWD9g0Zk0Ai1Jfg
rx6UqSLPy7Vu2bNfCQ0/w4SHdSmSUOy+YeMiudbPmU9T+2ZlcC5L37ZmLdl88lcS
vmw4tqO6ok6UhIacRISSx9aw51yCjNWHbEzRSyhH6dAM/hGWOuXetSjvS+E1y69Y
jXMciHmmErlYwKWtWmmL2w8J1yEBhogJgoQwXi9CNgkKd91iE1RWTYIAiwqD1a22
T3prFjWewCcldUjizaVqyg5KKNASo9DiCFBksDXIrPSQLsVbU+Tx6RCbHcKGnHyl
N0OqweQRy3dKTgYfgHp+W5qlAUotebN4qbmN8iX/u8011gvJ9OMgJbzm/GxlES2s
EBKhhw1D/CnwG/5xFIRvX4ZksSAsbdzabZ2Dx7uDZVD6CCOsJdDNZNdtISMctQ9Y
XjlIVBXPOd/Ar3NRmAAreoneF1TddGLw6MOuTpZV5vo2avo1xaL/e/CbXeDWXPBa
YagFY9akFPmc8Cvc3/+T5x9YKElNGUZxuK3N6Tm/vI9jyu/1rac2ge8bpR+ASnAr
6sUA1xTTDC4EtM9S8SAjJ9uA88VmcNN5IJ0enGngdmDEg2FhsMJR1gEGdNhrpqio
ph+px07ELWTlJkzhdkqPT8dDdvAVhO5HTRy9H0J4fgnxyk1GtG2t9rye1eRz+8gY
lffzhEsq3ZOPpxvIpH6EysFgt+XxemLwEXPUoQBI0kZwLb3AReHOBibd5vWSICiE
k2NBcHB/18XsIFq/GWOPo1di+JiXmGO3Q6tm/jTPQ5XMBjU0jkvVaB4rW+clhtyX
e6oQ5gouluryt7N3JP73FnN0qgIx686ekQYvppo1J98vFjR6cm9Emsl67e2BTAfz
XJawk7Jmxe4CuG3HLMRpntTAi1xmBhDe29fCaEeCGjdr1As/TTtXkMvj9nFoMFUw
S5Hni/frXRXqQ2kVnSw5WAlRaOKqGE71ObgWMbuN+GLIPukWolbf5PiCZCmdaopo
NPsydTMyVspPVeAcq5jjPSXpKX46oxmFjLykqp/c2WxI9SoDWlyMMgks+qU66eTP
0VYvpDFmHE5UEnUpsFWYerOcHZTlSpcKt6LWoBTn7iC5uL3b9lGkQy2ODAeKiwKZ
7drSFF9a0Dw+xb7ExfQcygKGlep1pEwJsFAIYrqjF0HsWzb1y7+0zW+b5IcHM0f9
chPyfc4nTp705gN3TCFJmrZFCViw3cKXlLBLdmDMI5a4rwC6gBYReeG73QeqTTFV
yPNvRcKVJ39rkc2lfD/eJrgeA8utFudnSXA8siR2ZmbI0HK+p/nAELWIv9NL9+2y
h0FUo8xYx3R3sEvdns8/bhMlhNPH1PLtxRDshPiWsjoxyqhV6EjFi959f0oD3Y6H
/N3BDPfD/xBKTw4uuRm7GkYCR4uZDp1z4/ZC03KGA3V1rBIUylZEGZLWxQHdB51P
gsW1cSCX9nLbcuwCrmXM1mL6HorusLfxo5pT8Igt18Oh4S1trVfqffg1LjTaK0Us
sxqdcXX8IjqYGjpnC5iZlNWJdsG7hIONzCo1KEYldz7Hovmeg9ITMPS/cH9AWs0D
LXlBKIFR6FXk62TYWmKBdVEH9ZB+WA+7jJoIoFnbewiXryzfLjPqShLlh89OMZDO
v0r3j5O5cSj0zLxlPmekQt02bTp85xaw7zCwTAUN0NORKrZ8rRwyHJXB92X3o2OW
uRgXObDkAE4fl2KD875PzUQpLBJ+0MDljvNWxR/IS2w6uc+V+orIDHTvVMsLa2cp
XKlpkP0E/elenC8cmorQjAvdCgZZubtI5OAR/sc8QlXNHPn5GqHHwrE8I2K4I2Kj
9e7tu2l+3gbEX5d/Dr8rvQSPt/7gkVBj8UaHXY+ouDAM06Avyn3KCKYyu50v97TG
58C5vM3w5gzNA1qaA57Hi1zgiPg/Q8o0OkruI49TKfgvPF3VIRXCAzuh0H0qR1ut
Wp7csuw9TbQKfs4eTYv/bj39t9DE8So5B+Qkd/RQsrys/wUZe0oGM01dVZKS22pd
EBtb+WjOSWklmyL8G3KhsNnO1xGJf9xaDLUxJpJO2/gKE4IA6VpUJF3bewSL4a7I
Rl4cuhMhwbZ8HTVjmTkbJwgrp7/LdBlv2batkwBCiGhGvPLzViGOQu2C72Ez3+KW
AdWK0eLaw7YWjcYhvB6Dn6N8iU3OBmdMtvRvKWWoSD7rzb45KSjGUrOh4G8lY9hp
UEf2nyhQ+Am29ItxEedHjh2Kwt6eTeCKAejOh8xpaNd9N6dEk8sOCJ5Cd3AHk6MI
ppI5TvB+t+gTIwBkyDQg56N4FW2xpkVANQRrR2O4zBBjffZIziiqzDk7hbj53EKH
KcfDvFCKSbbNVpdJTXluCA0WP1BY4XJMkA5nkbO6RNKANvfoLSiW02GxxuztTDbZ
gYvxBjHKM0cTn/QqR9yh48f0bF+BvJl9oXprME+RM/BdYDgN/lHc9I2aksfPXh8N
0d1JDJ26XCKfvhgr3L7urlyJE8SwJqwgjdv2ew3QrPzvuT/VXPzzCcEp3oH80oeV
VWhkFNshKDPTWsOi/eoa9uTUPrFtntuxFXwbExaD6+eT42D4BIz4j8o9j0EqWM9b
exuSd7E+G8IINuapMh/w/RgxWyeAySnYgWwppbVuFYt4dBuxW94mHdFy+4QR3seT
NRaVcU4GBdD2J08pUAViQfOQvsRcLqb9Zcdrsik5lcdecGnQFQVGrkh17pJP7j3p
+3BCW7Y03Dt6wbOQPmo4TqFDC9m19qPFZdBOV//kBqtQGqe/aVX+Est7V80hZf3C
HsengCe3H2xitPVHR/DnQBHEJHH5BtaFMhTT8MfguyiSSOGAbVsGtFiQjHvR7eHJ
sgGgUuSiijUT0CoEyHh9+NVwWLFaVcYRMWXJuoSTr9jwUVKGVld/w1F8UQ9d7+gi
kxmmaC3ywlYDKGiRqp22Cr9VTTBF+CvlZPqriFbIb5qTDhoBW60qKqsH8YfFm5Rl
Gm+e51YtNv8ZIZuF4TVXdgweLHA78TlWeABtCjz0HNhReBILYPkWi7emJj2GduGI
07UJ+P0ICiT6B9SvK4bY278pzpJmnpRkzmOvea7vntuXSzgdVbd8JAqeDH8uKFad
bL6/bSjBLqqWWywLIz8G9y3TEGSAfMx/8V9XhBkS5pIdB9nbWeTczJVmZf8kn8lT
7vJs1ERtRYQ9UUpW6yRwtQpUpBwxxIQBy/gWdVCsrhBDJiHdG9DpPn31yfcpaU9j
DZ1lQdcbKUrLL2UNW5ChxCVA+On1RUSq7XP4lH+wbQmEVeO5H5oiraKdosARRDUc
ydIvzbLsM9dQHrRSdeTZR7+tOUAcoSCHwFqMgJ7WvYe1EpXmUHQb2KWdeTSvmKf6
lDbOPpfoxE9G2MutoFlI2xHBewR0KQuIB6bNCOAJ/0n/86a2d7oRbJwKbTrOFniI
uZBFyS5yW6hd5aUc6rji5VRHlxhhcMs0dqEuxUFNqZFFxtl0kCwLaK1xHI7Rck8I
mS7I/9Np6/c8xxqll4ynagaiQgRKrVQdHhgUV9Vz8JodQIxDgJaXe4O0O48Wmxcg
isfN2SV1SS5UI6YfvKFl7tYgDvoRPj5Ex1aCoMOIFxIoYkIYV41YGLvLxrnalLjF
vgY1UBHPhqMySgXI1BdWyDHSq+cBiSBhZoBStegMBjLbRx7WPxu0eHWwJT/Dglp4
TKPr+iydc23pJuXP6x3rfwwJR8fazx7HIDhkgRBnAdMNmzgNFCcEWvnCHhxTDE64
IjgaZVAi+htY+YzE422db2DloThJOvj+XG1p+SGx/r7W2CVKEyKci6cy3BCwBa5g
jDVKc9VsFwXFnSExF+LmZifxy03CUUPvgYQNybSKRtnhTUkTz+2tvsyjWW7+QQBK
jI0oI07w+PK0z7Ek1whmjW8V1LHqx4W4zq2dET6wsbfghrtr3F5LHaUGlqU0Kvx6
qGeeWCRzK1qf+AhPebZo+P62PDSH/y038P8j5CfazYSE3x+qqs7yoCOxbnn69X94
FhquYA4MDH0Ygn/u45r+CSKwXdIHKPKkokTDjM5Dq7riVyA8p+Qgp5aXmkYkOrSB
lbyY1ENs7zDPsNHG9BpToExwlAQol/ejac3fRHSggILynwReMp2OdDheW0HlynZA
TWS2hAjYURnDo5DmJoL0QO3L09y8WQkOzz+kx/pbBdqgVr0grIKhIkQuZi0RMp++
TvVAJX+xqLJq7sSAVuyPMVkwkoxVewiNGHNHaEZKhx750FiCY851qH3HpEbtQZn/
b/KHAkfnhRVMVD5T8DWFRvdn9vXa4ofqpnSnTFjsYLAoUpCR+XdnoLHe61aMhb76
4w74HgPRqauc6CoJm7Ux9/zQrR5NUjLvk690ddrnGu5yiMRxbw52PBefifq4IQqo
mz0vdK4bH4dIHisFmoij6Rlo9BqFEYNcGcl6lLFRCzeqHXiKmA1pBYUAqGLNoNdA
wzaZk8LdkmqpSYscfCX0W4xvfGqalenjPaIY9zFuscXdVVQmJPByrgIjezOeLQre
DnjA7eDtECnfePOVpEgGvGWcCSXXNZ8SXNLpvb/P0PSc4vP0P0qmOE2cR+Q5SN/q
jQc4MMZWIAC25A2+UcXu8Qj+Cnbhv/Bwd8YwZ8dKyof2OMMVsV7yUCcegmBWGFQh
XeOgBoP27+1AnMY8rXBUg9ZzSjiG6oqmdGflvkHEpOtIXr+PZNQzR3hrpf9+gJDz
TVj5ltXrH2y5IhRJTZQKMrlzKU42J0EDN3ni7r36breYqIYPLKMCfBfRRwl+5xUm
rzqWUN9IS6Dmt259j64OpUb/FjJtNmX0xygu8vc60EFiQ0Ng4fAqvxyO1qpb9/aO
8O7K1NmFpX7GG+HBxJQXSoIX3XajDIgKU2KelDvTnyPo8gUlJlSVWw1mCwhoV5Gz
w0FN+9VpFugiK+nljzaka7HEkzJhJJUs7E69WSwa/soScJl4i1wBk8ZuAOx2AJaV
Iq5JTZtt5H0XxQiewq5QK3G+v+UuxVkDgXz3JCSKHDpFvho9PIARV9AMipaRG+T7
12hLQjD5w4/D99i+cflzAtoWk+76UsZhJ9d8Pr2I6DQh261OUeOrzaz2W6pP2SSn
vLMqfnze/ZisSLYbmMfWDcTuzfFliIIX5DXT9xIkqlJTLl6kySL0wIZMY42NXl5a
s7U07aLAX710BiNb4bMIhTgHZYhkuAW8OKobVrc2DSXZxx1QxoogxH7JmvnwEeUj
9/rj5PcPCvu3RwGVG57jBe90OwY6JnhYAdlAAOXKHK4cF1T45aHt1d8JqKvyMrkh
rFTHgfE6Kz/WEJTlvbS4KjMiaWnjVRR+7JH/yoP+blsKYLQb346b+RT5zro1K3Jv
QFMeubkchOL0LzNvTaya/MFU15yA+rNWs7Fe4vmCs79/pxTyeQ6fZZ4Mawyhfgo8
IOWksRRSJ+yAfuWV5kj0aNVjTp7uSolrf2FifLab+5m590B53jNOqi4YM3cnNX9i
2eIbKumHARgcb+gIMZ5WvGLMOeD8a4VmOu8A0LpVeJx9zRbSr1I+kK/E6NPJ26A/
59qOQYSR6vUHpX+SIpxoPCxFjoT8CgDZ0+7CEfLujhsxyW01dFKdlDyn4IKQgjfF
aeGjPuiJtmYMNArdBx3Ilk+egndCZt0ErGANhiUfoMbdJZBW8N44eD/ZfMBq0BDf
dSN1znn2mdUWK27OfVntSMnrft6+KDYXMOACALpcsdfvpjluw9JD8DeykqoZooSm
Iw7Ihc7PEPCw9ASObo9FdKgcI30OksFx3uOU3tJkTMl2GJbUk1WHrWm12OSDU8dd
mF5Tag276onoGhOYgoybbdtL7Xzt43GCTunZrFMzIPI+7H2/bTCxkplI6/Gs0pyz
ShM9q/ahdTRaMvDRzFdSDV2ifYIIzuYtuxUVausON3SzhkW6Mqe+PLN4zSsD9Ycv
Nw0ZAyip0B5X/IODcYJlKtv8SxeWxxUnTZF5ijuymrk2PR9FsTUIwKt8f9JZ3SYB
W6Gnn4iU8AfhZ/l1b+ut2rbZJSgqGKW31oyB6O+UjwBrG5K9rMpovuIno65xMtj0
NSdGodkTQ6Qj8H1uNou9Dxo1F3T43BKzca/u4UAvJ4bmajn9rCLVOPFdwdhJP1ow
kkVRthw5YEcLPsxrSyKohClCN53QTDZUwVaCKjark9OR+gvzfxn3ASrJ6babDFh2
s7TFNReHFQqPFvVqqonkrEKWNlQrByWPFkaykMsm/97jRq8eCgPysR6guPOqYbRs
Xt5VgWe1vCgNLt+TkI22VjuobsqhXHZ4Mc+0YPM8GTjOKX60PEZKuqVs9vVC6S85
/51j7/Sb2bV583Zn3PR0PPOt8PIerp9i2z+f6HqxfCXK0P8Rtt8kIoyFA8XpvC/3
fQvlTbK6KNAFwZKRw7VD5nBnfiUbGQo/sENBtVkgSo82cd6VXbbD04j4WMErgueB
5DfX02jaTbc8+1CnKIepErbyasEv49egNH9dD4RG2QXCQvlEL/Nw0rvwHYXFBY4J
mQe4QCLVFe3eEX9gDR1uJx5wl2Lmo7VybzIm3UsRUF93lLIvUUKUZ7gfQYhLFQve
aohDshdcFSsP3X4qD2lZsHtgWdzDcR4FSIkEya/DNYrycvmY1jBoGdvM43A87YnV
B+OO9yKRo/zxQJuRC2OoH5aGOv0WRCrHPcL03guaVZ6qyAoicTH4DP7ovwgkvA8o
A81br5G/m9QmyhJXqLx9hvs7Ozc+rjwlOx36PsPgs+a2ANtkQc+VhKVNw2Z+cmG6
i459s7l5WcyR4v62gwjG2miCLENtclXC4mi0nqcZeeOlR8ZxbIyM4LPAXoCroNo0
RdF5FvaA5QpR7sR2nZ9cbWNXDRGyZRGMk12ol7hcCOPgADo0mvSAUMazb8hjGelh
ZGYWbHDSx1XrKFdgOt/gOYiNEpC74+47FOAjgMkUbPJ/72pXlrSqGl1Ov4DWges5
P72iV6Ahf3otah6n2Ry4nDS7Qb8aOTZURNncl7+KigCWbGmYCxw9+QtdVcCz1KNs
Ewf5wY/XxFDb8HelVqzd5ypBBasq84cV/ASAHXdTvXn7tPiGUZFK32M2rpYxKxOl
1+NE2F4uY5KkPV2ouCzGwHV+QDjdHVhr/X8RwbyHEXvKCSAq9GoIL6Q7lmuVMh1K
haTdBOPvxESNGCBCDuhIKlcJgJGMXOM69NofpoHeN7FEhAgcbWxnOdnDEADEa4jc
9/z+K8YMGvxXtXJDY5Jo6I/eXPRR20o0kE+t8Zx8uzOMfbdYlwXK40OYNywm0vIm
gZAbdxT+slC1cvu4gGI8JSP/BJ1APxuvFNcnTxGdFvPe3WElY1TpT/q5uiBGk4XL
GDi7/Em1I7J9elIYWBktLCPhXKTCaKvWmhJu0vwCBE5CkPlsxizXWwXnX530d6b9
eHl8VwiHm2ehNC70d5AxZICcR6NMhy0QcknWeMW4xSD8u2AnUpi0epQ7yen/yIhA
27E6ychuPpxnusBb+/Am4ew6FxHXjMn9FOAEihgBRQAsXEv9FjIn3rOJvAXFWAm3
ufWWBu5Cl7VRqzww5GMNaZwUIp1A0S/2vl9GiTYfJDvCTp9EFElrUZ5GHmbzccI6
5KAkdFGNvR1YjuEP1EkqUwFTlbapyxKj6P4J+a+D6j6eKtxn3behJXeSRYVq6/2G
NinS+DKOe7FEpPICfMthMxyXvOyUcJN/KPWrKd/GmCe+SDtWQT8E00+7fAB3IWr3
LrOPsC1G6yvOjibTOa/nmxt9eCZ/RlSz87E4qUXZSdRV0kupc4lLI89xd0nkn/ED
L7Empu8lAnbNNeWmgBbaH+FaJTvLa2JE4lHTgpKbrNsUBIzMgGMhdpQT6ZdjTaIX
yXJaBAxDYNsfux+PM8Rq3aV88eqygt0gbA0h6i6VuXKp7wBG0Cpcm/R2AHo1TB6g
Q4qhUYwMrH20f65hRVqQVfjdZX6Sm8ax+XLoW9VmSD/lCSq+mrd1M7xT4Ky0kF8u
qxUojoCCVC6DzLrCLKoM2HDl3cw2PAyd9F5Dv+xT0GF19VhGtu8QurZqkgQmmiJj
XMuEYaVp8RYwjT+7x5e1bCAmF22nWrQ+A7TDCr2TSafl8aRg/3O4LtbztLGXUUuV
pbsI24mEhYOauOsQsjaQqAJuZx3w7jJupcbJF/qDqlgDU6CjUyp5b+BMIJ+BtGrY
3y24he64OAiRTdKQbCZV7UEZEvFTb9aqkzSBbI9a2wpRpHOjMsQ3vLVTh+/97XTQ
P1TnVKza0B35SQZNkDmt4ZLHofsCjApgfyUpOD/1uw1g4TDrp+1yzvCFr95ebtcn
37V+hNGTPqgiJC28fxbZFRSa3MlOuzaZWwULOFZ1s0CrZoZ4IvXKnh95bErTKT4m
obKv8jlqaNKa1GXMsqkhz+wqOYJZBPZM9gbcv1D1I1gBy2kVZhbwaxKDbw/IsC/B
9mnsk6dpGpqsUmfRRa97bmTxG+h3DyTIZNVqHOJ0RYgf+WhFyMTcc/TCeY2iyXGr
oV0gNSyMcDPM+3q0r+73LOtOsBa4qRzaHTQdD/M2UhtGAFlfVfmnDpMQrhjqjw80
hMLg2yP+4bK5V/cvM3hPgTF8Ldoq9zbb/NmC/IZKPjns5Bjl1DAH7zaVQvh7763f
dew+g1rU7e0CA1237Y/yZ9pA+XfOuowvzC3tJy2HzZf2zKaJL0QjeCU/8dK/wwqI
TZ+N9WKIMJqbnETm/4N2v/AOslj/avYESe6AjR9HtFbAqL1bppS8T9vYbCHUcok5
Ts7AedpupPWlpQz9qB2JVUEo3tPG+htPCKle2GA6QVRdQucczWPoyNES1oKyAU15
bKkqzyabA1q7bvo1GU378tunrcYmRBm+aDV7ueUcd531HoWKUy4+CGjb78ifxQ2L
SDfn59z+KPWOItqLgv2C3uUv4BT70yVrIUodN5hozHDRyIfB5ny8L4FvEA1eFp7k
Bu1Wrb1T/QsLAgmZDeu1rAu87KlX1dYUIQn5v5vQ7mYZZLq+Wmz0Ceflk2HHDW2e
t7JPyr9MlG/+I6oiw9AEMMGVw5VT1ZC8zPc9LD8DebfFUJccO1pg460J4M67In6H
2+YZ4XSutIUvQv4a1lgCDWpvHrJGwfslFgP9Qte8DG+frK3uk/PEMw5mPe9SOWcc
87NE+ODnoTQ+iOrCYw5XNOeld2lKPNMIeRm5z6EzvJyP40gEn3bmiHTLWgCttPwd
x3S2mGUzI9wQmzCUKuJTPQpbsX8kUuPYogAHxbZriJH76nwi3r5tbOmJv33ReNg6
8q+3IsdVAg4Dos6O5XPgaB+vgcMwBBg9Ak/SYuqIkfztzYCbL1Csuw21gsnpKCA9
paADs7OUieRUN844GVvzuFmlI9/Xsbc8XSYuuPHdJ68RFdz30vbtNWTeCirJlK/9
c5ZbSjp8UwwlY6i8gBd5f9YkHPkNHyocQREgWCY2vodz8p7LxuaPaiebp9lIQFfb
9bUx3MFCMu4S94N3hqITPZXrNWHXXurgnDff9Pif4xEFk4/QdIsC6Qx41SwtQ6BV
jU/yBnfdU0+DxxCy15mtDA8Vaq4+yfnwFTtsJRpbjxvDlVqC5A0P7UvS6r2vTm2Y
MmM/HGsl5xolCLWX405e4f/WCrdRW536m6C414x6JJrVtL81xri6CdNj6UN4dRBU
wXtqJc0oNAKlGL5Qid3oI74oita2bHUfxgminmhRtj4XGhPe9K8bUsqItCs94hhF
Iu02RRF4oluTRfjZObyYYCMEUoIwbHtX5HC+4OUA0Pbam59NajqmeZyzwo0GGzIe
+YYh/ps7B1GuG+OTu1k/a9rT0BW8HPCs5oHmE3fj3HS2WpKhI19Mnwl5B/Af45kz
i63wFfGzi3tbxjsDuoN+cIPuxuVd1GGWwfKd3tFB3HdIgLBk5lPrO7DGwfpkjcV4
tk/zrHVnse2tS2MhjIPsPJO+dnoI9Kn5TI2eu9K7muBC3ESHAIjfoTNMvBC0KSaJ
VDRRgEoowWT11bTY5vkvSCH2n1iW859mTUIkGxpG1EoRPRUaTjSqh5xKLH0gqrqP
CmPe4K7F/A6T2O+zjqy4EKtmUPvDbGtPVoAtIf0UQ60SWKCm2ssYF6F8CxwGrdyy
QI1mXceUkrORHO5SwasxtH1GekYFxFxXGTGcIODqdA6a10KbuuAyw49xRVmvISD3
SmUpEC/THu94RxOI/3VkRQsaooTQzVMYTLt1llkmgSxV1C7seXrewNq4sKK9cTwW
LOYEyd1/WLi3Kc20hl7+Txhn1HymCIZSuZF2haSFY7CYw04upZnYPN3atkTndgQf
wJweynS30E87TfiOaJHTecv4Dw10ywbfmOLVB7Jjn2FCCUqTuocEIpv2vgbTapd5
ebU17pZsCyGuITIUZKksiWWcrDijzz48njmkIQqPCA5Zm/m5PTdzd0ahN2a/nn2/
hQ37Sxt82pjvDVZ4ZlhAmFj4zDhL9cRAR77Kp0uyRVpFVYdUe2nKNARXiF81bFuE
jVOux3vb1Ij+UVJMZh6dxnei/h3/sUnvxAEPZ+rF/cIbnc5NKmmItPk3X4W+ZzZm
I7erDmOqP4M7/LjcUhGvMt+dO6FYnWPnfF/PeSBkO2HR/06TBQ9g5yiznDWl0lWR
vuc5jZR/ppHedngcrc+xVWSxmEez/bCgq+sE1EFw096vQFotl5QMk1wnEgg1ix4k
NBM1g9y/reei3qOt1tA86Q2vzwFCQhI0Mif3KbVOkt/T7mbwMhwNvgUigb+CEL2M
Avb8bZIyEcB9qcjVMidzHp0YjhieSRMTkNI8OMYprFVFBwetgGavjb+y4tDhU6IM
4cQKcaHbISeiZjpYfwFyX9HY846JjFknlha8nNn970N9VP40Nj8pTOuH7xE5bvnE
kYmhawHCNXi4ySR8kEkA70xhyS6Ov7HoEaN5f+SJ7omXdWrQ56iH1hB61iv0KoqC
Z5/6DgQAeOKuYJMLRCMsWl3z8zlqE567IXZ9ueKW/LoYC53pjTLZzD/tL1nTVb8P
oEv6j+sqppJwuHPsPYuJQpBYANR4yhVP33iRLj7EkjysxT92pSrELwgPVIgAlXkB
ezJUoQIWhduovHyI7foMPBLUMua0TBzcZzL3p24ic9SZQ7glng6+YKhh1S13WKC0
cbg7230GkvaXyzAjuMqHKU0HnRRwtd0RE2ap4iz2FkPUu0jIoOg7hcbib5nkY7fP
1EYTCp8ykLxZJkX6zO2NgNwR816T5avDN3tWuuTiAaDVGk1cVqYTfBSGZOK+DZoz
M8hMZ8pL9Jk9WiiEIfeHNIvw/52LlgSueF4wE5ba2yzP3/rsJaB1YB+pXK4PBtiW
VPE6DeYqJ1vURY8NWEXZ08s0C52luyjHiM29vdqyyGWOwtgeUC3k1N0vEhAhqieB
h5dpcTmxhYOY5ka7yro6YlfVc0iLSdTyw7vCVZgcnW8xyLKkZpNOS6jeFpFmoVRX
MgFKsgO8tquaLOAToB2Z9gzMJIVQE0uhg+NaK4IrUz33P2otHZQB8NGu7BbPo3FH
ITsPF+hM0My0AB/86rP21rCIjzeYHJkKNgjE0/uzMuWsx0jyId8bs86mNEhosmUa
5lYAFEkNCE91uH46LeDt5QK0w24hVDB6wGh7kfQOOhpCm0YE2nUz9Dr00KkIHqAg
rU58lbZBUjzKpxpO18krVPckg+UQUeZKWQGIG7HjV4sizGg9RgxPgv6dCFPsn3/d
qarl7WH/yTRb3rCFjOBKogY7DBnx9xDJksje0DE3l1ojvChEsG39bkuKoOI/qFNV
5KY2nTWaJ+Q13jJzktAum8wu5LMramIq8+RPUsYXyR2tTL7lLoE0s7OOzQygU8Es
G+upGuIC2aEw8MuFd7rjmMkPXSc9YoHa+/tO++Mv38FMnRPMgF2XR6pyoFoFWbTp
JXU393PS/O4L5fm+ZQtgFHr1u33Ay3a5pz0uySnxZhhK2+qaCLiMgAvCHNZuZfZo
6cChXnebHIfifqMDvNBoRg+IUfDbgpESDF8sbUDwq6YGfwblWZvwQAZf+44elfZJ
i3K+JPzIJqYyX4H8wx3L8OiG50vohEDfPzzZx7nfYHBwL5/uGl4vSCih1XG5Vb8g
PtDumHUATCs039cQgsY2cH81kfx1qEhYzibMXneiRFWR6p3pV6cZixVMj8frGs5n
duHfF2p/dEDd2NExQnrFljteao4IGJ44qKqsZxw3PYStUzLyL1htOPYCIIs43liw
Wxz37THZOC95J+r9cztoEMhgFV8DWXT07+XPv6GUTGt3AbpjDrGWHYo7voNxOla/
t+BjKaug5GfjMydFVeqlDbAz7hKtonIhYvfgN8WmYvMA603tiMN2TdqG/bmtkPSM
F+emwy68qtjD1beFbcKRMPVQ+I1lbFmwEUNZXhk7u7UHh95KOnIOD3IqadDiuSjs
aDl5OYFLt3grP0k7Z3drSBLxgYtbjeDS+wmFCXIvCcjPcXsMg5HhukqIudoP/kP2
i5lTGhIzIvsz8iZ0zZHz15+GWl0RJ0fKSRVQm7y/PceBnnLzxs/W+/4Hkkd3C6LW
77aqD0PVl1n0cDo2bPhfiCJeoBVF6C/8tRbbhSFDAXP9o1acx/MpMm9cBewI+geP
N4sK1D/EMo36uAr9KqMZOGvAoK6xthG+Uqn7/0yPmhUn19u3X1OjNPUSKbyZ7axY
oAlOAcN1h+Eq7xtfBs1HiSPIj7annyssxmYmGmzVGx//1qvSs0xiDhgpLWBCe2Kf
cXGkQyyNYmBHbqfvJb+nx+m+4v/ApqGPztnUDo6DxC1D7yzEIw7DR+wAH8gVMtKW
iBxBa/Gi5nhVvMkQYrdO7H9Y3/Tl6WtzbcCPwZQSOJ5xkNnSx9zX0RnMTqc0A65M
c0T++yM/5c8OMlrib/EJpooNuC8i+DZcu8aRZAP+K6V5tSHsefhNJ3A0A/XtCB1t
BJLhZGLqjWwmT5z9VEyl1J7n0AzYnpDCHBDwjZ3zBzg3TlcQV1c7BYJEFkJZxbfu
F7VZcynw6E7RQmtXlaje8bMYL6FvTMSzHjupCYwpfqaF0Jmc82kdrSXpkh6qZWk4
f9US47npFDKvqJxQHRwZyLKosP4CJNjFtG6lokrHm/ouhaCwuQCKOuyXwRUDQjYz
hCye0MqEDc6IScHUAtXi3pDBdLF7DLIsOrO8SeOl5A27bOWyARdeH1wTswdIG5xL
xY50qHtDfd7kCHkb5HWBdngNXZKV8jkl8gdwEYJYtMFwUwuKB9E9vdJ8iBm4tvE6
UTNa24189Vkwf4JbCfPpbH+BwL7g/fXc+YL+u55hdEblTcoZwqUk5I6e39L+8ehO
qjXal6qC93U59UNwCD0Abz7tEBTRrpr+D5kbb57pYr8ROQDbx9sxy45gBeST1tfy
7Nem2x89gVk7iMp0au8iEkoabResAdmzDJYm2qgSsZ43qPMRrQlVlSAzRme2Gghj
RFa4pqfxo5lJnIDplKJks/+bBYYbd4/qwRe0N6rew05LfCuyEuOeAeq1/pKqHI+Q
gl2Gql/CGxq+FqdTg9pD1CVobZXcLBpdqIIEJAoSqCYsQ41KK0vdfL4L7CyTZ4tw
dpS7rxxI1JKBrcYgTBQYWdWD/STslnUfyVKBs8xDtQhkLwa2JsL2QfhRDGT3/P8K
/VDBcEQBcw50Jh4LPNb7IxVDlwQ5e6tv0Un/8a79VOBXZCOHBrkI+2X0hY+/BtOw
SHPVL2VvYrpR+3JlmC5TMRBV4tgDxKBZv4QsTkmTismNu/K7wv/ps0IT9zbvld4c
`protect END_PROTECTED
