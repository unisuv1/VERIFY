`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jKElefbhlAjAWx7I+zgUf4N8zeHyziJ0Q0f/mtgHJPLriG8JiWSDX8xnvPtQEZw0
LCKvZj6QcW7J9zm0CvLiO4T0Wt9yzI3ozuTjyg6fJiZfwS48TBfzdq1bAASIyCu+
3R50EJzH4p3fAw3wf87ibE3Cesd4SU25EMdT8y9YmlMILMnFHGWLj3x5tU9qWbl4
VSi6ZENu9VAtmGMtHlEdWnqYI8x8xK1/OEjEVSyCrboflgTDTt6ZYHwRonNhIve+
/vhFu8LZIah+ZLlIVYgXxROn9KtXrQCMeeAHbRzDstLa6zVVXqHdBcJ7YHm+sfOm
U4l+JoRqBr7B0rKWABWp5gR6v+C9bCMnuICmGWi+BEHtPGh0bWu5RgUYo33pj81H
hvYUj3jnWbcB2kH/YhQUTrzKHPgGiJkMy2GTVDLEwl/03OKOqEYKL34O2qmUnT1o
k0QGlDePigfEKuI3PzEoiGy0K6nO1eqh2xBAR2wx/DEw/5DSaHappGWtwN3ZwsS7
zlmCU9Fnr9qJ3/JckQdWHQy4STWiiToNTTuyh3+GOs5Fd17qkQ9InJ7oXpl/FlA8
lrMDK5v8yFljGFHJELub/XpUb9zjxM7sov24NLzHUiQUfkPc0BRRaqIrih5EBHyI
5P6AHnuo727juVNb5qKmlTEwlsVoj4g5tI03kNp39VgJmuyh7o2bWHim6aN4XGVy
RK7Y/Ykb0tDhnAriIM3LhLHRtMhVeGMxinU778PuICB+JuMkX/BcNlTmh5Pdt/59
cFHU/EwqVl0Zup6bAL4Za+FxrdpcU0B9/9mBh0kSqCQVInRdmVmTc45uxPsdtprw
OcnhqCs7SE5RcswexJo1rNlv9yHvy0Kv5nZahnNataL9B6TPYEZgYByWtlAkanmN
nLmsuHMywov6jMfz1+sut14PMdpPQpMAvHy6/jJoOfBG1x+MvFeZtgmkNL5cdKe9
sdmMFIGfmkvdRKHHgP2pNJmEuPi2PlJiaGXMpOe/RVXzWrl3mgZqO5RzQmElKjUh
Fu27/7JM/Xqu3PkjKhNVKfY/irPqbJtTEV47Kijic2Qf4fbuj9QlFLuBqfFY1PKQ
RoHaglsyIUncPWqfcPOpTxJYLXL5N3+9AescQJxqHTjBcAju62bTaHCBfqNjoSeo
d5x7elmJDPyO/Wgqo6crOadXDqHX2pgehnCeo5itnFqSSQYhJRQgFMQ87Qvbdg0O
Gl5r/7APNlltjRv4ewr1NWPtyEplK7YZaocaS55DDM8UUV/Cn1O9Wq/NmEjlA5LR
pmH0ac9D/ylp1H300vcturX64vWZ6lDw2dZf9axWh7TUhSu/5KrFTczBp/2ew+Ou
/VXqPIAZtmP5REf61yT5q84V7hjFscLieGoreREfqOD+uV0Y/GK3f382mKxG453h
EzuG0SVuXgUDg8AgihL9Qd8Jq3OtL7eEugseAppHIYWQu6JP4K3fpOSWLaZCKQaO
EuuAJaioUI8De4kUMlxrTII2UgtAsigI0mY6AJ/cq7Q2C4dwGE0xerDYcxAOpwM3
ZmnXMAZCy9LiKjxq4wZ2ZSbDllGRx1BabmsgTlSZdD9nPa0c03//kRIkuw1PkGDV
Rp66emakgRvSAvYcDiFlFiQJ6Ss5LIfmjlo+pmtSpo59UnU3SAwQtow8LONkFuY4
qiL2i2mTtH7eCe6fCowZyxjT40W+7kn2hscOvj0Iw/7bY1Urdp/DqGOJgAq4pPGU
IVh0ATG4pp5ImxpZ2WvpcibeggZCWpl0UcNGS+NxMNXPAyTP4JKN0P1picc4sHZm
hU4ZhNU3hmTNO4KGg6lZYrxpeWJoIuA7jto5SBD6VVIB4bUe3NRUxY8ULs09AL4y
6ErSz+qhPOWbzVAKRtB6cfIuq46YPB0x8othAFYG6xjwQSVgjUYqB06lrNSzFOgN
f3AWZehMzqNvhY3KmyF2ncHVI9s1Y7D6djZrTfrNV3SvS4Q/JFtW5uMpIcjTOyGs
AB6SW0bWnFD2DxQ3U6mIi0kLfLfp67WaG5yj7lqgrJWuNO64vz1IcrynmxGQlhtn
VgoVkBY29pIDi0J5tPOMB+pqdxRVn6u/aQhi9n59z6RY0WXE2Pb0atpJOzOqr8w8
5st3z8S+mTQ0VNHH+P6lAOEwyIArOEpg404KsXmclaZ18ikL203CsydvMZm7cHeG
OSBgd3/Kc7sRtNLNmP9bqPDdXV5uSFnxbW3T5SgfCDP6emvxdpgqg8w9ijOjPgmr
ma2yV5ayq0oA+tOhUGfEd2L4FtWor2iPxt4agMw83A0aQrCml1M83Vzzt2ufCIVI
5MJkKNFZDKeTPukYSAZPkdo5/dpiaqjwFv+T18/CPFYnFG+Rl4CwvSaClEI1NS1f
D3RhWRAOP8B+BQw0L2scNDmwegEd40R/nxAGC52MOyeW2f9rNUXgf6hbnTbdFkvu
Uj7Uuaew1t2v/zLu+zn8P5+GmHVp7Tfm07xAsPqpPPCA/gjPokRJOTnHwi3TeXG+
eseRndq8isrEhY2UNEIYO45xbBN3aVYSbSf2FWP5bE9IVKsG5y1/4M5Gl/99AvnH
z7j/d9CMFRTzD/VJvf6IRfJJlSBTFuXej7dWkzQ5OmQ=
`protect END_PROTECTED
