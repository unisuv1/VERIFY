`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fOcQ1PohIDBhvD93593niuNng/BpXHnih1nn7uJfCr/ueeh5k9Cp+QcLw4DXxewv
/nLAG112JqrxXkI7O+Ksw03BCvjiohbv7hapXgbE2VYvdFAFd1SeeRN1ZDmHfChk
w2gdHzmwouxdU/gRnodPxsX94VlmzbWPYXlybgWoOlsUzfiXciyAuDXc1m1EpbUd
lgzQzaV/lVF6oWLrxU5Z4W1Tod/KU8+WgUYHT8fW4fjMmICkq09Fo7Q/KJ9Wdk6h
AJ9hIa7CdtR6qn9sBOqxkgRSksJqEZE7I01hox0FnPqvdpvZtscuFonBpYbeuJUc
6CZfvF03T/Ym/pN7+HJ3KTO9Kou2kk6DnczvM2pCq2tUJYA7FEldCr1Y/Ua8Ut67
Us2N8RzM3q5kKkDrMkI/slhMNA93J27L8S7PnIW4KVGFGmiT9tINMjylcdybS+C7
bZduD5Ho+71VRgvhrTFCSwLm5uQxxi64m2OEfdf2SMFn9D5T8zmM3cEeIhOOyRSU
+AcaeQA/P8CGPSMBJvlLlJst52DndiSE0nADUJmaR8J7XoesGSbAJtj+UBYhPhQN
p8+juGiiUiwmR5NUTUnyDymlklXoWTY1s/JIxqmqmRRiDXHJ+WcmUoBpM1g/ncIo
rE7GVankWkdVoZlXa3qBzabAt5mbF7NgwhG4Gq6wNLWCYQKs+HIcHuX74wQpw7ps
dpA1D8OA5snaRH35JWuqgSdOAlDw4qICniJ413iDaAfg/z8yfPC3WHLwbM2tm8YG
LSc3deG98aMUXG4by83VKQFUf9EnTBviNZ9pGmcyU1ipFh+UFDfWLCX2b/fD8CXN
ZzbfANuP/dIhrgBSn5cllPlk2BVvKXP4QoW0+YlHqAdJ4sZPBe/11Pda8/U2M5gy
mIWFddaO47tPV2oIGT2RJvIODWe5KnyMeYe4s1CoOYUrnDkw+u3/zxJGhO3yCxVg
YoJ4MdXLZIfI8A5p1HtyWV1MDx0KLP7S0Y1C7UlBfMx5JkwtgrCbPqPxHau16wQe
Y6oiBcNDG/LY//aCxAQZZWLdK01XoAo1Bimhv4iM9poZ9GcqnpQ1zibfV3D2o8xg
Wvz+TgxurDVCMFTCoG9G+NXs3yUnmmxRmXu5Q9ydadGvwTO1B33PeCOGUOV+H0zZ
lqL48FLL/8O9is/Pqj8/hsVfIfAqJLvi7KeUHDgztMmJsEiIA1IMPr4ANiAJh1o9
maVh/sKH8sFZs7LSX75OZMH8qxTumGFSoapuEDfchHa/CccGJtEs8UOOoQO2X5Bs
`protect END_PROTECTED
