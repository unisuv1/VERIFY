`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
x3/nTDqrAXDAqhB+hC8eDYhJ2G3LhxRCY4ICOWj5u9RQ3OwkpiVWQHOjvOLSVYYE
lb08VL8F1GvrZczeDNyoRZezs9GzdXf4WYOSsbIln5emftB/YBJO1jAJ0LyysUjC
UKyhkh+Z4mJY+dTBXj38mGU3hRqTQY67Tanh+VbxDDi+Y0mklae/6ZuEGX12aax0
/XxP2l3nZ6NU7cZ4DTQ9Fg==
`protect END_PROTECTED
