`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zepcXH7Jhbkbg9gg+zlp7kTSVEARZN5xTOMC3iuvWtks+ufjp4wzIxlfCQI1i/vv
3TQEglZiL51znYn12qjnZpK91PHZFoNe2x3C3ZW+3UHY2o1cqU/T0CBGdRANXU8C
DOk/46HL45QJnl9DrdPct9mq57Yyd3Rf5N9LjowNY7mF0FxFATSbUZN4ng5+3Fp/
GxezihVT9u/SIZcoXdMheTBL5plJsKaXuD7DV+bL9ZZr9UW6KHr6bwMawpnKLLjg
iOaXFbjk52+XkVjF5kfv0snOwvYUZDK4WyVBxXVDMFcpDTaRdX8ZuhL61jSY/1U1
6nw748A9HKx4AewyKDtn96jR61GpaSL6cwTdw5Oz/PckbiMYxwVHX3BWoHAQBya/
7NXgPRNggC+h0nNcSsTRmLbm/mbja202hQ1BN9z5jgnAxmBmCqaShQQGQNKkT6sr
44U1DKfuSq7lKg5uoPclVF8gekOHCgd19M9pJbn8t+TfHdnVLSyR7zQlbx0Fm6d1
YtI8UZZ71FTS/ksSUGFoZg6YbenepqQBYVioY2uNphbW+Nwa70Ul8thTWFddwk1l
Kfz0OUyRCwlZPylcXEo601/J2B4O3fySUpJpgzP7x81RlI6msVz6ucdW8aBqlMWY
YUhRXTY4jqr9+GBswFRXo2j4KIY+qa75s0kDc99C/3uE6jeg/x/COWPAT8ZuG4D4
lH5hC88OrRxqIB7uhQmuwbpP9PM8ih1Vd9I46gtGu/VKxTttP61nQsp923+xtPyu
cX0mMpegZeQmYyNobck7aiuIHihmDVHUQCmL3WjYK7gP6QvGe86iE4/kKcLr0hBJ
JDO+0a0i+nmg/KTKeeptIUmtyg0H2kf2f0hsmFTWzKxHT+YZsja4jV8T3Yj0lvgU
03uDxhr9Wwf3dKQ61zL6db7uF93W7jN/RA65vfpB5Wb7B8DsyO7B8JwoWoBVAiyb
bsbW6p2Lhj9fjaUdKWfravvOSG0G2g9bgMz7DE6XFZiewy/Ff9s6SUABK/IA2ydQ
mt9kmr8d2bwglNMQLpMwCs8g0MH6pwOxzSw8BvtQa8jid3eAQgCRQ6av1aq3lD08
gOByHxlYLGfXio1WMmuGys3qUKApubO0gPyhrAlpOCYwm7xBJVzdMee4ZXYHqKa0
zq12xifOyBY8ajLkrxBRMubcUp6BHrQZJpmMiB7jJ284+D3AgZJIn2tYnCH4YNhb
NV/RDOl8wtvjacqTkje0bO+W1oipREHxA3m/u5ZZLENWU+ikhgqmcmQO+WbsRywr
XS/WlH3CK2QSY0xpXi5XW6WBG1iZ7M7xdy/Xgr4mzC9Raayo+HGQbHYT493JNMR2
l1kN8ZvPvfWC9tiOcDvjfWJyh3V0CpAK4fuwMeq0yfTyAg/gpomJChLgxpGY6QTr
GS/prFp5O2dnkXYWkxjKBoxi98KJ6Y0v6U85vzm2zpQz8FENYwDaNAppTlHYw6IZ
mMOwDDIsfd4p497oGsXpFFzC0GfOm9u0PSSY0/xkquB9iODQQLG7VIxABA9gVjF0
BwFApKjuwkK3mU6DhDl4VC4/cVh1f2TP/+rHj7PEVG7QPBuga09TrhnwWJjPOr7u
hKKQZQuBkwXHlKA22M4P3upEuXQ4SnJ5lKSASdoR+jf56XqDteVunyirPrYX7qL7
eet+RGI2K6/1EJjhTndWkzXJXvYIixJYPVg7ghIsJOOpUMJPmcXLojl2kRmiCu1a
NvXmrYYf6hcsNo5yhfllig++AuBgA8aGFDIOvMK05pf15wgIvwZq5OoVYOCmdbrk
d3xWUd9ihSfF7KMGdGaP5evrxSqTWW91FTJCOofsodrgsJTBZGvKn00D9aEfbSB/
dIP8OXHEtaCTRpnNkIO7xVTVoST+jx/7Cy/Dq15c/JKGssZW8JsAghVWTlC/2KUP
QJMTZEzm8+SpT0PxNEaRmvSJEJbkAXINTmbaeCNqe1UwMPG4mwQa+gxBrLE6Zm/z
TfB7JyY3dnQLyB05JUokR3OKCJQEsfL9k7S5b5CXjbBt7vQqcMZ238pVEbxtaiu2
E20w8TuTKI+McNEXoDp+cZaE4D61Ix8ACN7Hxt2N8CnMAHnurG6TwieKIgrDuqX3
v9lKR8TBNRCXMmIZH0x//91l1lm8k6k8NYJhX0rz41UylcMiuWWZn9k7JdhUeLCm
GZURtLLlfXen16fuLFryss6mbzYKfMK97119tzO/OAzzfqTlBkKIFO3YIctSV1Rl
nMXpiW0phLHR7qe18fOMkqKDmnvdB65mZwqWm1THDTXWDibXe1pTPW3RRrU3FErh
Hxk01YIlUgjDJ63enf67QeeRX+uI/JHW7FWJ5Yi3TWk7nr8htfgkC9uaOrvnRMgG
5TS22WPqHqtsGN6X9eetaTM70PAAq7OHSNWN78mhToJm7wnS3JBz0+vuVpLbyOkd
LRt3SYplehcB3RCZ+9yHX5zu4uNdKEm77vH8EmJy/rVrxow+O0ybznw/f2+Nv+rW
ku6hTpbDdkA2zlX1KTrYr+nNdm+bpkaypSgEgofmIajsM01xk6aNxEVotBngzVNN
vBgjNBBSK4WNZ61zVq1tFJcWri4CB2wnxUKbLPpxnstPG0ugAos9TA6iCFp0OLXK
sBK4DN+ilzrk9CakMbQrOM8GX0CW0dDx/QG+W31QH2RgpgXcVkO4A7p2DuxYDtkf
bSRpTJkOfTZLHtotNNXUMyeydDn/UXUzhTQtu61jS96yprUsnu5ToYvMdjvT5T6E
AGcFTHG8mPKhteq82rPjxsLjoL3U5jAsn6KUa3HGhpQabpV9L1dkeq3BpQVLBuTq
3S/URN9K4HgM4+7VJSg3eU9h1x/gpOZ8poyr6Sg1pYMQxDOtNv7rc4J8lpNsDAW8
E+eOEkg34PCxdm3vJWnNrfHTuByOJkxSE1JAGctcPwqfd3LJYNCyxyvM8TzEma+h
Sgr+cc44nCsCs81cJbzNvNz2sl/TotInjAxCsJEeNp9elb05T2GOZViI1j6fjckO
hFGSidfKl/3Yr0gVVb1fMeSJydfzwgJkw5XL//PzKZiF5nZU90UjtpSJ1iegsM3c
32Y4yheyvy4Ru0xiiITfLBB/96wVB1dAwCIVaKsO87Xh8aCk5u5EC1VEMeq2WnBX
0H7X0APi5NlhH2ux/+fCkwfmoynsY5H/Qkg+JFgIGo4wcZUeZn+x3Gqc0z59prM7
FdWl2NNDjyWSgJUDNKmewD0w/8mW85OvgIyCdKaJTh9No7XChRQM0Qr0joBI0RZz
hHNz3SxKJGLgzCCYdBbVYmZrm1wI3Yf0aIcb/H5mzDCkgXFVDytOBDBs2VDL1y+V
18jj/rl8OUvfC6PybMNDG7VHg4BvA72MqxJHRBe080/0jbCJYmpKYKWtoP4UzeWc
m8ijPdzWR6Jb1HNP8eu+7aZOdtqokkkiH4ES48pO7ZVaLcTenxamZJ+TgBS9Bx2p
N8/fheQvG3k7Mf5EuGr6nEuat9kdlmSEk/DQT5EjfMsbuS2sdPbTRXAQhvQpUhNn
EHRaKA4/scNAXcxL3yFH33GMhPJUPEfZ9DceNAhD4CzF9iZpmaghyCq0R8hSiMAX
RlfVAQZF36KnLxlY2J+XlekSd5iQcJq6zTerxk/PU0PLrntwGZC/ZF2ZnCZpAoi/
5N3aGz4OjYwnbmvp+WZC7GNpOfSpoh0fcb23XLYQv3TuHXaep3heSoc8h6ritQjd
epJcEIZ65MkVR/MvKQKnH2kPzF8utrBcN97OoQac3ns/dX+Qe7fY0Iw2E1LQHDUk
yWFr1YLHzTNmcB7gtc6jEQ5LJSM8Vzdaf+qIzFJG/aUedfHtGMhG5osWG9/TRJda
Obzm8Q8wgXCR4yRYKyZyn9R/g+le/lIkEmm6wfnhEOcuzTxYJElQQR3JmCBNd8m/
+B7E6oiqxXlhoZWpE4Ljev6cUWeVMS2yW5h/jOfAUEIeyIpl0hq8KRz12dHaTyVT
swRXOdhy6qlW9kBHqQCArQEOAh1U9OXHIwzQyzKUeGnL5HQb4DLuTvJAIRrTNKTc
YBixz6t67YsWFm7iR9CV3j7iXnpMExI68bjund+nM/FwV1ViJtxqucq13KrNLlTe
RSanynnUjTJRdwSrMRLognzC2X7RWcP/1n6sFX70UIQRb1DjkYsjA/kc0jXjc3uL
ExhwUT6fYGoIblMcBNImBToFDLE67wuod19tJxiOzzH3k7POt/d5QjYmHbmF21FN
hEHk9KJPuElGs24xskUvzCjv7AtK0x5/RImv/3m5s7nAg0WPTl4MSER5iR8KykXL
o7TvxkasYGY0QOdrUL6hHL+iPdZV8WYF88QzgIedLqiV3OyMgNFfbgiyVeiKfFD9
a+QeXnu3ehyqsQNXmf+9dtIfzCQ5ThvbQeLIZX+gsA9vI53I3fHRaD5RM9f45agk
AvpKnANxKySD+BN+mDKeU9C6qiPDwAPyvatnmsvAqPdrbEQxIzCr6nt4IsNwfVw9
ZUuz2ZanULDU0vFHyyd7ZhGjmnYm9gHQXD2Sp7zIZnpF7ho6R3DTh0A0EyW5DkOL
TLgsdS9bonswmMQNo7FS6e5AzdwzuoMTw9/R8KKrKpvoMhd/G8iklB//BDMziu7e
WOwB76YcCO2jzpytHEBa/u8+OpS3QI/SPKQXnVc1rnwOA5Jnj0zSn6mak8M16T3l
Sn8rBeDS3+Jt+U40bY23YAfG/alkw3sScS4c21QDYWkjlCp+Xk9jV8wKxzrYNZos
VnKAqS3SgTYkyoWeR0aXJJ2YfcN2qdLHfUnq5JVUOorwo3LstUxgfi+BLng1rFe6
kTxAtopE5AEqTDijNKDukQTUVXMlN/1wYQpMTjikVjw8Z6pDago8cxEwvBkMV8VO
XVf4Rwm2dI1UHKHcsAP6GYBIIKJTQt7CaPKE/gIj8XFKaliTdKqqvQpj9HAlzQS8
9SMcFRMmVwz3cSA/m7m9kMjfs16Qis7QViLfso+2nQOJalVhDjjnWvzRmI7UR29J
nrCkpmvTCn/4+CgiWcNbDy+BC4Z77p8qU8sqjmxGYAheCDRFnXRFFpDkW1sRg0rH
PUkN5XuaKIagjQAx6WL6x96GWRr+12M2lYSBOYqBrA+oLVjafaHwWtWEvCaZ/38N
CvYt3kKGs5xS1Qfcm32it1szgg/d1p4KM/6PHgE3fR02xvGOoOwwXpRKalvcan5h
eqpJb0ss6WlRC3OxdkrY21zsSPhaQ0pfVypBcwjeQxUwIw6VtJQxWbsctUAx0OvS
CbWjT6upUqZB3GOpo/g4ImFuT59k7QdDVm+mV6jrCrzZk7M1xRXQOuIXlGtaR6Ap
U7M0DCSitQ83vp1N4CZzfxxZX8v3Dov71/eGvzbhpNhupFQno4kCuoeyALWKLFfJ
Sf9c0nm7xcghkmJRqhpN1jmgwX+ODq+OYdfJDZXZfy2+qmrXiUd9uzG0EpQOczUd
UR66+LASbB7trOfzy+JBfi6cxHeBdF2hIgfw+EJOGw/Lbr1Hyi1/SiTWyMVZmi0W
2bOPgVScFIULgg41TQBRQvg9HJMlCDMIAqD3wq5M3X1KfZUt8zsBsCKyLR1LsK8Q
/ZwW/uggnD2Mthk8bgcsjlkIlhGSuxSABrkorm84g9QSKeXdE+zFfTwMxOWW0i73
yFERRdFg7cPklEZ+qCVC5DkqNHHjh8rvWiSWWuMbLFIZ59Wn01AshU9IX3eqr7w0
iU+m2/HFnhGyU6Unkj8/BC+opo/wLTdrAXMIFHcaEHiRrj4ElF0upDADQQ8d68XA
GWilNJHHb2tkD2b/E4FmsQ93gkvh8ce8hsB2He4RRdBMBGDXi/Juk5LQULYYAPGJ
JKv0KErng1pDrZw61s+CnfARJ6nys9PW6FtZQQeHxklM//2q1PrCrss8b3DaDpYD
CmCPYaWQvnnYmBNpLm6p7MsiTfG0NAr9Lf0sqP2sHoagCW5XvUyWaMjyRIac2+NO
76bxljKzs5UipzNUcDC9Hw624oSnxlaItYsR4CXLGJyeahc9isTZLpH9c+7tVReB
dahq5kwbbzU8vsv01Wis4LbcpsdP3U+pw60sUqqdCOFxpxO26TpxB3iD4Rw2srcW
iZYVyeqS+TEjU43sBgn0i2AMPYiXTXzEWyFWO97SZBOZEO5bdRdKYWIMDkjYpFy9
sSH9UQrA0QzbLZ4ym9hNwrj9Qa9rZ0XJGky3R2JvhZxA4NhxqIF8hnD403gQOSpD
TqEInIrLQVyB7hB8LHcRbgbfxq4E+UVtNQ2tgn7vSi27KQkNwSqwgSO5kZx8Xfcf
yCl1w/BvkA/3qUMtZNmMo/LM9MsWy7fhrfEmS6p9SdEPa/MRWEfTqtHIKrXt3Pkp
GaRU56f1qsOFg8QS3F4cdskV7f9CfC2D/QEoZYww5MPN7fahKp5iwUEuCl10jpXe
YPYCQEirITCu0kzfHAMOWN+8K89Hdfy5YetiAB+nPOQYPHIY4FUFfqB08r1kXj6z
tRa/U1w7s3A1p53oyroYpSzG9ogMuw13EZhn31/Lx+qIM1Pep7jXPz/yuu+6QFBt
DtYo7pMkw/VUP01K1F8AGkQa0cjJgrKw38f3r9m9XlkKUS11dRcI+0/b6vveW99t
8Xh9mo1tYEbtw+4xDAuSAbr4CXWOfJr+Hr3WRvrFhEaaJll3HrMoklGytAJuPSPw
Ve7U8Lq0Opxj14sCEnamWVr3CCXa67dsLs35ovKO0HHn0/09sUPfrnCtvml3/z/L
/vQLBFp6CnTaB5E5isYajAQ6lh/29Nq57u3JMs4NPYUnnME/ApyK+YuU/8OW5M26
mqeeizt5Y78JqVM5Oj9uuZNQeO1SClsAsAWDVMOz/GztVGi2ZgWA42f0r+7cxwq7
eFpN+Q3uqZo20Ri6NqBrpxLcggge/w3TTTlEFmVkl5IwthfPtWUSUn984DeCBnZS
ZLg5rWNHX4Y7nllUNV6Buud6reZ06vRCLNRhopoaDzPk9qPwkzSlnuW8e5X5bAQG
vClv2XIhk+fAhxFx0IpgVblmmv1Mx95AsGbpgdOsvrYl1nJIHRzXvMIFx4/QcLQB
xEZ+hfJOgrabuisBHlKjFrGs/dOGHcYRTxpz+l3MtDNHJ2MaxBbDu4hn7cbXvO0N
imiB/6N3KnPYlBXrzV7DijpfoA6YkWNNXkWQxzXfHyfrcedUdAHC0D0UVc5xd20R
0GG231+VZSFlkbubnaydtLDDMz2uFsnrvPwGYCpkdizhy0YLrDXW80XiR8GJAPs1
EPsQCOlofKtQod0obY0AZ133CF2XLPeoWfqLqbOZA5Pa1M1ICCqJ83ZTTJ2dF9HO
QXME+81M71/hKhAqcoO2vw3pQ2FwIGa0Tqj3O7SN8KSpQOA7bbDhOC505NMbBOkq
OQxIG8dXkn3XE1c8QfE9vMU6m3KnpdycFebrDK6Qy04a+CcypGT0JkUezT8y6iZV
SQFiDmVBuJsKGpOZuWYvSt9ThcPHmbZtla4GWYxkHj0+ki8Clo4NoWFqddeLGXTk
9seCg1Yd2qAPKdEaK5EmMUf9wdHP71yiQSi9ye6V1gdQ9djUAdn6oJqv3XTUNDNn
GNm2n2zJ3awJjtZA0SAOEpuX1g8ys9selt3nT02y7GMS2waY1uU0fjk1Ovk24lb6
okfP09uiEiFqh9WsTPr8NN/K+78VYZibX2n4vuz6K44WDo7Nisu1Hg6qVmI0wx6M
V0u7fJlW7FA7a9MBRv+szudD/etwpu5g8rt/lXshcyOOmc83/pIyd1L/BYOPiwf6
uOXYnrccbS3gXXpCbIqhdxBK/nO+awNxAC1stCP+OA8YTG2aMlsLujvue98YOA8Z
4x43GPgnoO0crkDV86Gt2t0n73z/flV6Xhsrm0he7VKFJEpr/GYwdH08whpNxsRp
MzLSfQ5sxQmA8AhuvTrEo3KO+n3y576iEnQn3GX3Hvns4lShJc9L9JEGIWcRyaE9
p5bfcr2VmPz62QhrjTP4xskYgULoxwYpfiC8TKhbpb5iIsL5XJvnXjghueJS1vS+
VkeJgRVpcNDRplVOwwQg0KEA2u7o8C46QY1iXxjNltzTqL3RrpKEpoAirzfzkQwf
ZhX/KYTyFKk/horG1x/fR9u0Q3VUCIbFdd/UQRkLExPPETrMN2gKjpT9XsKrRl8e
6zz4/urilFIjdZG+ZebDITa9mTut7D67LKpLcT5HbvccZrBM4ga+47my6DMn3g2L
8mqXm/BkKVLiIjIRWmbIcUHhwU6cJqcpRiLAR4R2muqIMxn00Vt7C7zGW+b01QIP
NrU+o4l+KC9AyoEIax6a+JGFjIx16O5Rh5JCA0KKN68amUhQTlHw0Sem7gBQqPAB
h2sf8w0k2qwIbi8sQG9Pd9fgGYt25x5ZBDoo8jLCNcPZ8CMwGrZvhf4vWhCbWmXN
3Cxdak+y1yslWEp+2remt+FlQ6POPqB9AnIR0hsUgHXxEDRaPy1Fc7bYxqXgZibP
L5wbJaIoAEPspGmOSjkzafTGDZs60FY3v/r/pne9ntAUo/JwREog4suGBCM2kx4l
EgMMiDz2ixKcyfpViJvRpqY3Gmo6ZncSmxYoDX/TtC7n7Yx7GASFZ+V5PXGycNIY
CNNJUzWwjeraz5PhHqrm09n0j8EKKhrYiTHZ/QQHGkYvwVFSNwZm+UGidoqZjJL4
UVSC0hQlN0RWJEA/iDwjKvJibiQ6zO8FUPqVlWaCGaHgvZc8gGyYmi5L72wqwu+m
E+Xaw/m682fQfM/hfyystoeZMyRVLCCs2Qxsk0F1G+VRDJX/9D/si1X/CjdDOQGq
lPbzoQ2T+U4FzymdHa1EvAzVVL+xPfOfJe6DLOHg/2zYJpiQXm3+CWdGgbMUC2kI
IO+7sW9flJwPyp1xLL6G3+UNRdmqDCwCsa57/Kqc6iU4zKNf2B+XSoqc3T+Hobaa
cy7R4dqs0f7tUcjdNdgXG3vIAFc4raBcX3QG+bA7J037jvsJns2wUC6O2bNVrNrt
ylmfKwN8sEFiaeLbBh+rGbVFjnuFqjGLTXyJFj7UAS56iz8YYUlYYERLaVcNYMCj
kFT22ifMrFQvsqkE9ICMl9qwUqvZAs+D0NdPesX3L6289/6vSoFouHPfNhQoEG44
xijRFG8ganbocmPv8ZKb8x48CtGJmZ8LsRhfVl66ITE9Ay1LmWeEf/0QikxNqzFk
KldnKIPEXTzlldRl39VdePQ35iObtZKA87tRTyIO7OGBt20foMDWF8WANoMTTnEi
aEn2fgRN77D7obKXzraAUwIDbQUwVs7sdSheJd2ez7tzOwAmQFmb9w3Jdbo+fp1v
MQl40FgHkzwEpvbIUeY9wbGUOAGO5zwCOjet6daHckI1HQbQ8dRX9DErvuX7lrtA
RZhDi+27pR7NP+EqNOv0FjnUrKjzHd8GLaIZAxVCVFBbNVR3l928IXKM186RDsBv
Mks5zR2iNLXFZ82AJvvZNkfcWGIDcI9jNVZXgN93TXYFzP/yXX86wtVvTmHmqhRM
glp+iFMhZPsFAP4Zh735tvgEuQ/FrIh9BnVRtFy2vdxg1SmUCEScf9UWAzc/1KNN
k/YZFkpMO9XZKjcd2XfDz0gFHUr2ysoYSGNOcoeotmUgzsJsDOHtFlpRqIhS7XZ0
genSTP1dYZGBmouciLWWCJ7nEa5gVKXlJI+Wf+UjBdzU1IKL5f0P6DPKYp4iruNG
v1lPbZWoqy8Fvp+2Ho+2awSmQemfvcW8YnLHrw7+aV/O4GT0e8/2jkxzTPSCYAKs
bKBKr9E2l5i4KbpgRCjleBYRhv29Q3o2MPqYsIq9x2tmcm/mipAFOfFiNpywIfDF
YUkjjqjWHfkuJF4eXq6YYXcDcAOAq1uHiMG+sDfpEyyQ06cAZzBi0fg7Y1ff8ILc
lxgVVzYHTW5ot9HGpVhbGDoGlqAudCScXT9Dxmyw3fa9GaXoJdbKDhia1QPzF6vy
oYwVrPVs8AQnTjgvMHjj7up4uwiNytphpIez6wbW5PvXKQx1OD29zdre4Pa6d1/x
LYuwOb0bjFi6BD43Im8THOH4T7dtNvBflbrW1++OtNUGrAFQPOFe54YzmoXMitMK
1hrnWMPghHuDbxQuxH13MM4rNVKi45qFznWMPexiwRcZSWE4b8xMVdapvJa9bxIx
gGfKIT1pHft5lsB6gpOidcERzLi4e9ecFxrquLmT9w5f/SGR31jkh0W/UmWWz/ev
6wQPFGfat/72SMw2vYn7VkTzsOVNqQtCzgc4flxhkBa6e4cxyuWht9yGmuacqavh
Y3ADSiQ6er8UDwhQWIMto5AZnuof1vHnP5danp5x26pSXtciMyYSwK8FcDlRsqNL
GlXNaxT6hUTTRYo3DVBbt2SqqofWS4gc0TRwfiNPSbxTdthiUH0xVGIyViNXE/+T
X8BheyyZI04VIqwJln1BOrzL0Ox4XeOX7HgdDEH6UqkXet2fpOoZ2YA3cJuJvbPU
feDvFRA7bUCuTKvfzM45VoY9DsoW9UbIbBvNQqmxKPvaGEI2KDhLLerd0rNJ4Yx8
oUSlVJioYntn2HCT+UGNTSKnnChreFyOwoJfjpqfHQXV6RSx6yk09Q9TBrR09WXI
IqsW4KZwFiwFd9ZcembH7ZopyfEKs1FsjjndEuELczmE1Kcbb11LHr72sv1bsxNO
GsYS1oKkUCVl3yG5ILtscOVVnZDDKN54cipdWtwW/+Ien9e4MVAZTyPyGezMbHb7
JOKYKm8T4f7fnM6wNLLISehqWNRdmBJxBoTmAfnktPe76SavcTX5z9g1D32Wpd4e
hLD5Zqbgxd34cTCeMrB2zkHz1LuIA6LWwx6nAXlAxdj5z8EFFHMlCkjV55R/LBk4
LkI7XjvyRMO1mNLIwIfXUCWLYABPJ5Rnsb2h/7EChfjHCrEcTP6ItMrusdXx3KDL
O02FTnB9rzS1c3v2WpBb0MehYHnYb3KpHFRT/HG2Yr7lDUJhsGuqBh+8urYLJPRu
LDxQZGV3/i++eVoz8xC2FUVcFcls5K3/gO+zF1k3ObbtiJcZuh3GQkfyk7z+gb7b
N891qRQQEEaoSKbmdSymMMfC5AM6MHQ4EsAsNeIvPDkxG2WoHVLlJKrxu3Mi3UUQ
xJs5Q4k2w2sHWboGsluAuCRhbe+9tLUoRikGyaS8A9f35HJJy3S5FdV+2bFwEuGq
QTOXyOP356VgtacdV0c1OcFQqsS5SmRdHUqkd94uX6aQouFHW8Ej4VvRR0djO9aj
7CawUpJi/PGQXi1k3ooQbamHV0WrGBo5Pwt8NOfOimVn8AFhUsR8qglOIP33aTGt
2wN5/wLPvfEkvhQbfxffkPO9su8xVKmREhvTL37ZjDrC6HLTro1pIJT5tjKMH2W3
xrCfP0HNllA8hDgtry9xH+orTg3mkMg3fqZs+2JCue8+fDVxLjjXYILM1H/c3SX/
T4RpzlFdbi7hiVZD/XkYug4+Ynh6k9ngwQK5fNKseNwrbhwvQV/q3UnoIdjgJGlU
EF+rDWXPucAjupKe/M1FjsYgEdQrt2a1py8qstcUtqugWQdMI5Zy5rVhLycdwvCS
XcJtWs/K5Ma93PKGB6SeQCMJZovXoWN6CYUYY37VI5YUdHeZfAfIG/MR5lNyOeQ6
0qZ2qtnvzYPueYrUQkxynft9ZhCjPaSieHqQfTTgH6NQTVnMCnf9HdO3JDkLr5pO
9l+jazs1gJOoSY0iMv+2rwIDMJveV7COXZT39YqNzvkJcnU7/FYMVgc1fv7PMJd/
2u9KyRfqzIBJ9rHtTJ+KnJjiGWO1xyWY4RCw+BNomRNJYtK7h4ecJOytxgx+Ehnm
w2uhbppfcSq6QuJi1AWOq/mhzzXf38Dxi75vMrIBGYHB21mPN7N/CW7HPZ0Fw2xj
swGPHVejOx6Cn/ZOKHc0YS4kjkt+XkQt8yKxzN5fQVYsZ5uM2NHrHAS2Gi2ddG0d
kcfK9FTdFC46UIsK0yy/hJO6pyawPJt9+LOusp9FHbRRQT68smDbNqrZc+Zp42Di
KF7iwYinndWjL/O+6UPAjFrR68SWA//HWroG/JlVZhaq7OyKuv/Pd0tNzuW7f6X0
03DA3kGHmNeUyGJOewJE462EPqrzenTNoiAVe0//h/Oa5KLDZ9IehMz5stIPvllW
7QAsNjrQggqSPPbdkZ/N6YwYVDwZcwm3QTLD85c8rGiefYXvkeR4xdMFKrNkUmCm
szkSyR+T6YoqYFjKxjuPTiPXlk7IEyz5WPJwqC9KVmIbWvDbWrBM+ccDaa4C0oWt
+laMWeDLUBKRnleyYZP2d4c43s85bbEkp/BXOeRFE6I1UPpWGljJ4U8xMuYlxFIf
ZtMtfxZzeErNBsn+zigzwzdHxULtWRySAL1hyDWUZh6kLphsPvWHxULMvgYeSyoE
lyb/oWiq/sJbDtr9FWdqUtfH7o64AIccv5/S0UsrX02GAX23brNHC5AkoLgCVNlZ
Fauqks0RrqMtG8c4F2U4G14Piv5gcPtl3jse9RIeKhdbzIcke0rF4JMfvB4CZuMh
xPWmnWUiEmZcLw0w8NByarhA02O8phNWPaoFPKbnp3Y=
`protect END_PROTECTED
