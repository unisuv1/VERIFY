`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9e5O1Fg101VUvqfEx3PmQ8pk3H9W5x9E2UHZyNdkLzykZp1ol7aSG1YroR5y5r1M
sIticcU6EH8sWjIx0vOR23faqGXZXDB/SMNeM3TBI6YbQeSz48sJ7bZ9ZbfqrMpa
/ciufuaKbhXgKLKx8PnhPFm3H5rlK2Idjw0GV9+ngV8gE/0+8X7l4VEU5uQst7Pk
SZYzv7rkp2DblIujveD7oLpX8YuIkQOq0WtPVzc11jte1JaNRIMJFzDbIZu/ECdo
3N7okOS4X8EtcmqoEbGd//wC7lc/QhAL5tJ+ZX5bftofhYXsOclx0kvvZENNak3C
D8YJYEeDSNggUa23/l/thT4jtJkPNiaFrbxY6+SApx72MUSOcdAOpkkVsGITQlHO
7oCOykTo5w+l7W+YtYy3jmB6QEW//XF8DKxSc90t7JlNBpMsNqQBhP8MWreZ3jgU
ZQ0ZjfkNCMNPXv8yq4X3hJlAPiSXqHS78VKoFo+mPeRwhWfeMigYXekVxl62sNZT
B27EN1D1FYrziQQILobWEjVR4DTIhSdGU9PpI4dSwI4ntuaL6emufWifOgTrCGnV
WjAL/jhua0ZxKc3mhMeJj8uon8Er4rx18+9BERylM7vAbWtxSBn4+M9cFOju22Yj
SVPsjXxJWJny6R1DNPUfXU//E5YopP2SuxR6WhfcFI47jI03EjG+J/lMEwxXzqCi
ZTHgc+s8PSIw4DBaxVMhc4vpeo0jZe57NuJq3P7b9SYvBw1EwqYwNNcdUZCpuzCV
obzTOVkO+NBjcWHNpGs4EkAHwfKy/NSahQq3H+0KGVmZmcILCsDTghnQvqelufNj
fUh1iRyO6YzuZ5n4lAqFJApPKFONwVQDVzVyv/l4yaA+aoAacPPRRE1RPTFY1dZG
+cvXZ1K7ynPvKpAHJp2wcfTKoTbq8yoi2u7hN05Kc7CD54v94jhfaggn63wtZpDF
xDNOe2oWFZisNEmXou/DrSsL+N6ylUpD19YUKcaBw9Q88Rz7mB6PivfVNzPYbkKj
IWZVGQ4z6yCc4brMndDMAmmMDfxJIh6+Br6ByhxPwIporQvK2OU8fhvHB8ixBWeT
mNHdGEVAZtoZiQOi5zcNAmSlUhlQutpZoPLgHekg7DZl2+IP24zt/QiQqSqvmAOO
xFYf9lmAmDHCcuksbSDPFbN272yXgUW0Z7lEa9Z7a7cFQywdAoobliBTNe+Z03pX
2dU3tf+6VgJwWc+VcF42vFXZYBfqYO66WyLkze7zLm66dSaysSA/RSvMiFL1JKZl
WoCMbg8XP5CN/CqSkN/CRaqO+166k8Q1BTiiVRs6BpVK1azaV9ze4L6XidVKa9K8
buZJYaSSLZlMSwX9FVWyaEyeEvPm/c1wI9fntClvuPwJbRDw9SD/0NlCY7n9m3SY
mpkA3z/oKwho4/dr9zqx33dB3d+bPai0yTNawnH1+6Y3o73yhXjt/Z9vBt8p/GQB
OY5z9Na3by4/17ePnVOSYRC+wZzEPijHVpRqNd0zgj6Wsl7jsGyHka3pHUxfca0r
2yfFZsIo6MBeioAe2ZGY12qyQTATiFoKPgUbYUcvxGhXZ5cATLIt0yxE2OPYKPyl
8cmnUgRSothhbcTA2LWyICc9XL0O5jc1pXmWcrPVa7u9Dy6NRcDNqxIR3u/z5Rrc
ho+L3IoPzewnGNYaerwYzNDQm2ngFWToCXPTngDwVD23rc4xYDFoztzvgmQxgTri
6opvzf3yDO6u6LPqoYhDVQ4irlpSl42v3r4Ae1w/4eX0w/izgsKs3Kl2TcDBzDoo
i8d7VxneI/uk7NEp0LpXCbi8ITE8pK2BJObqCEGIwmXSpJ4QRdbGtq2mR0l+d1HB
M6oXk07NeJAya8vTcO+sx6L5zhWTzckfcq79ALoVvuRY2xacRFl9bwJpAKJsAKXO
oGG+2Xo1MrJwAb2IJPTMQze++Wnq8+UkaQyLfQ4h05Rv+6XgvxLhfeRotY2xoW/X
eFEjQLCMTXC7bYbO6Sh6AWe/9x+LWeYOonshoruPoPbUB867N/G28J6yrLzjGdkj
I6j23ST3gb/RCHvfbHnQoSF7+CbHeYQTdzlcvFLMdt7DIHmq/gWE4N37XfFGv9wL
iupvdyGNqUKn4krtL/bK8DS1W4P/vKUdfe5P+aJ0W1+phNFC6bR7XeDx0zNm/Lkc
y4qW375l0Kt8MCTIrNIszC3mF62U8tCKivqLMgvwFXwHwCi9XKhW8MP9681/1K96
Hn3iVJ0vhzeI6ibjOfzJRz0521Kjz+c8bPdbcxpmsLiEPPG+zWcigE6NUZTPFEGD
7dHsgUU+pKAJgFIXWTxHa6Ui3L2fiuVOo41iyMN3+0Z6vpxojPVfc4Fn2bPio0si
KojzBRw/Qg9ET5kfqpPgPpTHKVyAGuxxKosZAdOUTzcDEDBk27HftnO+dcXlqG4q
+Si5J9ZJ44zq7Vt4zXZKQpwPxZxiqqTktXl33/+Hw3KfRe5XDdWxNFdKkx6B8VbX
WveyWMxh9keY1PK8hjAKvRz6R8Zd+92u/G5luC8Ub+77xB1TbTHVVcBomXG8cxUZ
ZA5LdPfeOscDESnOpZhd0H8+znpOcPRW8ywD0qj6O0hhG4+2wZYBg9MP1Hgbi02G
dbyeEnZXEGU+fyiK8JHEk7o5QgbpqFzyk5PDXbgg/4l5Cw1CqR+cf3I3SIOwcgy2
sBBHAFvV1kml84uQBnUHomul7XUNaYVlB/KrAGMZn0I4zVHy2tw8iCCmpa9mvgq/
Xe5kWTS847JrUAGTzp5eitZ0+TYB7MpShNwdXMmOPCUZx3hwl0VplzgKYTUMFe8K
Xe4INB7UGG71Uxd/3LzXuaWN0QcpF1PZlnk2Rp8V6uE2JrmH8VGQeb7Tb+YOCEml
BLyy8p515DBiriWEcIdPkl9/v5nVzgQ4LAp6j7wOmZvCPzcOOckjSRt7+zNvMeuZ
olqzSzNIijl1CWUnl7/VmLh9TxI+MYqjA+OICmbRFayZhk/ojy50iwqC6HT5g64q
kzQXXsm1LM0a8TNlaFFrKprjNQtqnSnd/7D9a0YQtvzGmZzaftA9PRizA5YPE7Dx
A07x+ytQ65irMHiqcMDr1W6z6SPU0Eiw4oBLMLwaSg/XD3wm9zMOpUT8jUPCCPaX
LClKf5kE5VUDj6YFofKYuUwIsX+3z6lguSVb1aI07WH1o0KJaqPkzddrErRaPYKS
X2DLtHjVDt7SJ9+I1nAwMOqwHSFnKXdFPdY3oJsFWQgJL9lNkuaVk1v31tnH6Pdb
fpYQW1hnhPk6jlNZDd70PqENHVLh3RjVlLGl7eZd1RQqyPaJtHHzkY9wlssEzClq
eY+zOpesgdIDqgk1pYjVLop/h7uYepqRrO0tpaAe7uO2Vxu1TxsuIY7dT0ut2ejN
qeirTMyX1K7xRdqwQ2ooYxL6NvPX1V2ZlLvGRFVj7EQEWJFojLMuNgV6BrxNtplv
9H3gvftPZmoBAqknZSXkJ46lYN+tkS2GoavqsRR56kpaLAEGkCUAmvvk1zt/wvfb
lC+fMlnKPznnfVM7s6/obII8i5ALp152kStXakG5FC6Tn8r8N9ZRILWUXkp70y2Y
+qD46mnL1GVTRKb9dfvpH4HLLfy2Pv44HYTkOg4rueMUuRfDHEHiMoDsev3MLFr5
X/GbGpPwwaTe2O1Md95Apv05xnYP9yQZzcTbcuCCX+dQ8gp+umf1/RGPmkknpdoq
/oeR1k9GCdvZrEZET8OIkX8SA/PazDcAWOEhANAlqqMhAIw2WJUAgFAv6a3xpb1T
WFSx0Rm7nm7Ecvfltr5En+uOP2/yWj3q8svmT9ObDr+uGSCjqtb0qiMFuoZVcDUU
Eruv1LTEdh9eAli9HXFwkT+xphAMe6MY9sXq3fq79yOP62n9zvt42XkDcGcI0rhB
kf+tqgOWwzN+4zlmiy9B9wMsGrQyH4jxw/hJ4Yvdi2KoMKf9xCKmZTy6qJMuhWek
jK3w70fCipBG6xnaBq67F2u6dQTJ/LMwK5m7X6f6xWr/s3lsk1MoCtnADNNWMrkh
fX2sWTTiVR9zB20RXkp1zTzHc6aaIeZp75l4C0B5rFKjK2aPCt1pL7ZCTeRqSov1
RLN9NF/8HpEJyBoI+oi/1W1VioFhO0TfPgbQWaGqAywg2Of3tM6ZWUXDOlLsL3Wk
/t/vBybTXoTC0BSDUYuSQQZgUmNR2CUH7Ep07qULB/K1Z4haL6nxCVO5MdoYTl8U
AEIXGdyRkIoVTouTVBV+vD7LF9fLvqo/2HptHzCPGdiKlKW61yypmuQY602ciztP
kEOkNHtWzusZfYoaS2Yp/UDmkR0EQMoRxrIZTjss9osQy9fN3RODHxlsW96YfoMr
RCLI0n1t+tLMcR6b5nGUUMtoL0z9VbSkBfEDjRby3IZ7WLJNnfZa08WARnKghB2O
1vAEqGeVanbN/eHh11xLjoHFgZgpNVqPhV2X/faa9gNfr9ixiNOFIrNbiQsi9zMD
kXpQq3fsOf70nxqosESsLFtGgLVPAvCDtDWh4dRBW3l5LrzED7cuzfEFFuSJ/yFj
lM9bdQrGNy9/+n/KjGO02URUxREMzcdXlaxpJFVG4SmAPmrsyshE2NEpmnzwR4Ro
h0lzATbAPF5EM3k11YOnhdiXzc3qdtr0hP4EYL/4AH0BciIMWQpR0tRLGvZMByVI
GU6g6ApenszJ4YNDTHUdG5SpxDm0On9FWjDcnnIyt5bYJ9cmies67H6vyGEER5i6
jT/Y9GPk3a9J6S9o9IyCOad/NAMsI+P2Lr9zrkIiWT+JAP9VUP5mncmLkn/NQffL
c/eHRDj7gIMPtnUjaGrGy8R3jshvPgMdFlc0zKMSEsKGZ6pjYI1Pw/FagKNE3gL/
DsxTU/64GG1AtdDyjjlgw+2L/GAfovPPnciSWRJGDMK/m+shwlYronYHGmSjCqay
QMoliZvTfev4w1KCOx/i8TrW8TnmLflKqv8fgY4WWw/bPgCcjxggzZA72dteUSsS
jnkQJtjWOMFXSIMivkPZfQZOQeLVJ8OJ0k0OjZsDU3S0JqkvrGACZFWmoNxKkkrx
GD9+6skr9sm41sUsP3fBaxmhA+SM+YYXC8SBbHs43Nb1fAYGFat42+oxuErBDwdQ
EHjZ8vE2zd8FZhuqCRX3ef4AYCsHvof3z+mlnTiv0PlnYUn6OySLfn0fdOl1x2fG
DaQdAh0Z9z+Fmbj/F85cscLXNPFPfCfNuASWZoAW+f+wwyzyvxK+PfCYW8a0dsor
Icigkm3KXHdM8dJEq1jq5C9zjQEBJdKtxwGYe25LdRnsNsTElQxBLYo0zFizVbUJ
dVvLSIyWRnZXHM+m/RJElhAA9hjikmL+tccRVJH7Ns892xTbNC0zLKVSFG111fiU
0fW+iwqGLBtvfF97/vgmbyBm08g8N7HNbV5yg8LaDF5DN8RIrtH5OcmDIz0GGvDa
31NFpAr7CuW0vUG5eQWaG5sAbN38csUGGfom2A5ECi46+NFx846kStPxWmLcdBTU
vm1Q5XYV7n+FK0hAfPQfTHWSWL1jjjkqTNX2K7GfIuydnCZZqXjt78sIux//7Kbk
E0unPTWl3YAKfOpVujGcS8CDHu1LtOKw3EmSjt8IYtdmfrafWZotZU6wFobWQzNY
ooVtHVXud4tnaCx7ngHYTzqrvgBocOUY/LdDJSvq5qofIcwocy2Bsxo8qdgZ07fH
mmKl81vWdeSRl/z/kdOrLlEKjdizvsZ/ANtW7zzwBfLvpvTBCfZVxfTJa1uIOq74
kymn8ryiOZJ7wUJmva2gAMIFR7wfjb4DNQ2KNSF6ln0Do2zJFMQJVTEcYso44w+x
QN6Ypg4i1s5zhSF9kLUs2yvGFdifPngyex1gW3Ps0x6j6Bll5GioeF2KoSRAMtO8
BGg9doAmEyQKLiaB5LpL8DE3836DOARe4hrq26Q94EFKLZAiRFMCU6HR5iHIAng7
ZDwZjQRju7Y/m97q7GzP+MbpW5hXsbxVq3tMKnZY91AQ73ggXY10K1m+N0xMkIM7
54IKrcAEctrWmB5FfPx/hUwXVFFLuk6t8adxf8bfxYqebz6IPc/FxTUVbwWYV9fE
D9OBSdLTSzSGtQ10oDEVTE0oPSPKhj7Pasr/sMLmf4CHIrZeMYmKbh7Nh5/TRXaH
jcKL89SWVpSQxxzsb0MYgWSdU75P3rCR+EcAMt4WMaqimWdKlkWo/QspRJaWBfOF
u/WSxaQA9S3dTOPcAFgN/ZlSYja4YvegnZ6PGyaxV9kmQJ0NpNDegDxYIM2ZE5S8
jUs4MjdE8Q21iWSmMki2aAB9JgCTKs4UA3GWcTDHvDJXXNhudv8vLjl5K3IkQnIv
U/I+bFfMAmqEFK3iak7eV37rIxDWiO5qPF+hmmUHLjSxi/AVKBWh0NxC7B2JAa0B
5RKu4zlLaKrcKJ+gRrm1ROcOyWEGBp1ae1wzim2IL3+ti6r0nm4UTL90zdhLDUDy
2/yPkI5EDdJRdcJjlpsbEGXicOg04PYtG1lFw28MN0kJVH7LejZlOc0p2Vvuzgb/
NMwpVunuyQVce/k1d3/1etPf5/EKCiX3dpLhb9+gOUpBQ9XU4OjBYuWgI/JAZ4yG
W7q+X+Cv/uLHhI9SjRhiTrxgUR9ZMWpjlaxs54dSxApUx4R9zx9QeAaSNgYgIazj
toZ3ne06pbtR5PB1lFmb7IrIi/znVjGcTZ5tQ0mCJnCt8unKcGHNWB8plUy5lkql
12I5EIP2ynqZIHNQWrZvSL95GC0SNL46GHPBo2cQ2TG+WWl+Mw+U5ZVB2K2XhOsF
HrruWr3qf0z1Nu/nUc1FuHjqmGP1aoZlKs9GpD3vYdQoUUFh/lwb+TUOU1kJmhLs
Z5noXKSRp05XSsxF9U2mOkBDzG/9kkTl02wk6edviHEf5dd+y1zTtvTmG0bi3u5b
XIEl9DMWwOouuEIbrpaDfj5O/BXLmGnoHxDeigIAUVdmoRgi2Fn1HASPNz8tPAz9
Su4kgAPGRDfbmb5t3XAZP3X+dbOkLVoBbJfFcCGOi2wl9pfRyCphJ+JoqCSRhLYn
unADdORN8/ikXTk4nPXId9Pzh262mfEIr+yGR3LoOr8op4T2vZrtZQywOV9UyoGD
/huDZCb1lGSIAgPbFgYGwL89Nis3pBDhn9n0RXM+LZxXBk3m8Kbmu40GsnyDVCWy
ARv6VyrUmg2Wb065DS/6ee2WaXd/pq3DfOL/mFf1ljhCTIEcHMcv/WVGKGv2oif5
PqC8wgX20hOxV+Dk9cBcJ/PD+WD7MN+yBGHPTmP2l0Zu3qLwXd6tZ1e3bj4jGX6O
sw/ErtRkqDIPGDbdHDFeVTrZ0ZiX6a/s+y79hZzyQ+cqHbVLq88ntD37ZGAFgPoX
LwCK3iva58YbYv/YhxLYOw3Yv0M1keKHkoeugypvd9BfqPvhb5/y5qjRdi5i5hIk
KIQb52GxGE33OTI3RTDYg23rzDg12pAYGcKioSUQSFeg6TcQG6Y24tkE69yBuyIo
rOalVHGNtJTnXzJVxja8H2XVoN137F8rtlctB+k3UXoU7GliR3O6GnlEGEgTC1cW
Le1HJtBPVvlQeL0ecili7sUj8tCbKxb2ow1A3vkYp6YZd1510uRKvQYqKzoEJfhn
HhMffpYtLJK8On9s1v9R2FR72OcjiCZMP7mbnq9AD8mR5RfFEjA6K3lDF6oNXY00
agJc9W916+WKufPqPhFAtbKbEIVpo6Dad0gD3QpkJzwOF9tvgXvCufHuY5HAsEsg
25G7QxTCym3hD2zOvapUMfODOEci6Pz69LXE7gMmLaCJEajE+c+BsGAcu1MfHIEP
2dhjR3iqlS2NpqdZx9mdisZ7azkEnlYGtuwjMtZw7Xg40szi0q/HbE/64ViYoVB+
aIYYvnsYQwAJVMBM2BbyBQ26/0zqC9nhYRvJUEv4IWekDpm/bcUxSkggfIj6th1w
Qrl95czpyDc1IDHkycrR2a2CSDuDA7NLf4pMUXNZr2KofMAVDmrpTcZ98v5p/Er2
5sobM1NiT1AHXXlLcpoXmSgM3soYqA7UAE7/ACXeQa77BcG4AnaBWVXm3VXtvTb0
zrJqLmGja9TgqIh+s2dIh3VneJ5Maawa9kGei6OFt8c0WC13V1u5yPMfRFoBl1A1
zrrNWpwMLM5ENiGigxSX0EleDT8A4L97fA37r0RHVaNQF9bBAZxeMUuV91Rr5e6G
ZJwclEjDUfKEkdzjiCnN2Mnt24Yfe+VZH/SZ28JR9K7LQMPdvqbpvchAdhBB1Yiz
M8oWIuvKO+NvH57otDi/30rpCKqPm2NRJaLPBs4CRtkk/tGKRLstUe2JpcIkLoSM
4kUqD4Ns1D6C/kG4KG1k0ZAfgqzGZS8ORzYI2b76kJpXACIO07eUfWYY9o+ZDbRx
t6+R7EJjtcaBa2FP8Q07CbaL4JGBiI5B24+HORdI/Fs2Kn05mx8Ghx5oq2vGiQVn
lRykgjWKiZoUPx88TCqEN+hj0QnItCC470osjwrbcC5Q2rhF4B7SBzXlgmSU0gHY
Cnz0jqtyrcSBf1GUQ4iUyaBzHyDSgFbX4NvXVcOCtZRQGtyRh9HBM4EiUJJ/p2iW
+kjIskJHcVByF1UTNgM5IuUykxPUPqQW/RRi0qesXU/ZGlLRVsoE+h70Nfz4rWy0
J5hzFap6O4ZDXQQH7JwqkTYxM6j8z89n+moRqgcMLWTo/8+mRKsKeBRVoo2Ot2MU
wZ+JwyVvCHhmHGDVB77UDBa4qziyxXLWmq6VsAjNaDVzDw6pLSiV6n1DDmGfjTGo
b1kqd2nb9bjhleODwi6oO/zqTSrVdtpD0pl7jIsyAcvCHZiZpMqU2oSqvIfdwhNY
CJSRQioHCez4OwcZmNl/6bi2/k5MOHwPMTwtrTJmmgdMIW6xAlETWk6ReVRVj5Gj
DFhCdxBJy2QRbnE1syvhm8/Rp82yfQk0qmSizgZ49Cj8Hsnl0TnumRM0/7KJq7rx
4GP08H0cTCmj+E9X/fMz6LZG1uwRfLKQvHO1iOZ9AuMe1QFOwOXf/QC1kIuO9w4G
CZqTk78Sl5iLEmvOM1324mYbyD81BTqqXaVhJtJ6JNfL6jquJ9ie1WZObI/1DcSN
IVehLHOLE3Zvl1cEgS/TdlfpT9Meex9q1zucKh2H6ch50MgKSWq3HRnT4dVi3Atm
cscd6jfMGZFIGrJnYkFxeCmfeWdn2Ko5+2JmFGeCW+jbua/5s1NqmnUfjYXcfjWB
IKg5QzriqXC1AkRzIOeGTt3tzZoP2AF9rNeEf0PXYfpigGwLwaBZMxzF1+A7PFSs
A8rwnYVRk9keB0IOCH1cCGSLYnJ1oWzQjmutAAGO7vsGn3Ko+1xz3gHEJqyUM2jX
6CZdE7GnEUeZb8gFHJ/PnZdS8mQigq0pFiS5a5QETa/BQKNSrIi4Y4O9mlT4rgYX
acrcCay3kjotJLDSD0cwbo/4j2QpeJ1IndyToX57H94/Ep+zA27HKfS9Xvy08QNW
oYiPmJjezZlVko1rrHdEaQsdpCQk866xlp3v8HlaDk4NrsXvTLHhmtBjuq736Dqo
Dx3jgJgEz2V3fDkkFNUj7dY8naIDd8YaawyV3h05xNzuIjt54ShUSwgSRLH3YL5V
LM//j5zUPxgZqbNhNuWChK+oUe99qAC5kyXTDbkKdQOn53dke37/9557LS3Eq79B
OQLebIiKIx5NRcTiqCgL4MF4cy+c7SKVsrwiKmbXQ/XB7Ucs/ghzFo1ALQhl3TO4
1By6ipFdBejv2wYUckoEBb2OoTmdg5G9s4iL+IFHJETbIrME1f13xDezNZIKyfwh
qSGAyPjNmOfYp3qAJfqOcoc10tgjKGsGmFtNQ6+qDKavt0f3fxeP55KF6LYkDB+p
wOLrDRcEqkqoST26J6sCphqdb4V7ZpHpoBaPJYyHEJB5CKQCnXmijczG0EISmXlr
zcV0NtZIyII0VW/Zsa6dsEhQnk7x/MWKhK4iCLUggxPOUDxnbgO+I1BB0aAw7E61
2W/ACEv7oBY6xvXXj0n+7OXzEk/GADn0f2t0WbCs0N/kRBKbvaThe2hwQzEMEGwv
I78LSh4sxrGJ1jDMVuqzlu9FAYflDwxRRB/VI1qtxj+yg1yZp0AGeDxIJTaueFft
ZFpPtsN2vlnhycR3MO4XFq9+m6AGNVL50fFD448HHqnTahwHmNzs6HfHoalxs2E+
ItWssdgF0zPdS062wegiyevnNGn/PlY+mDM/QOBfb8sDPBHIuU3K5bhLLbm+aMkN
0vtInQE6oELzxufZgwrCcI9epPN1TxpWrHnpuGUUJW5a42FQKYMcWyFhCqkHzrsc
38ADX5iPoffE8D+WJvx1yE+F9cvMZxDtu6Vda4kz8Zb4qpEu+DRz3+diQ4L95VTK
0/qdQwhwfcdTHlN6sAt6IxQkW0eV/hF6LrCejqsprlF/cQqHzKcMgx+CfJlzXATN
f+mR4FSZHWDpR/5wjhsFj9u+nQiYBpeJ1ndWNaV5EHZhN+otTFd+D4guMPgSi3Fp
kBAlj8dsTHBamqfzK7YfnLZvgjdo+O8KEQ5/m35Gyo11+/QZmjSVRNBr6kntEQXd
60wBzgNAvt2YaVZbcxFbimwim1X1V6lehEwd3NC/c13Rbx+OdZ4x5HLUzTbwBQtT
+8OcPbLpwYUUcZvwoVMua3VviX91m9mQwCQejHre95ZWzGq/9om6OAPw36MlOGta
tBMrRi9KOuEucV4ce8JpMNpRMzWXJkwysUK7agewmXPN61DN/8VbTrKsh5wkjRp8
cHgSJHFqh2nVowoTMHFDmgRdoKzbkb+Sm53ndUviiar9TXVPsJYRgULXYvUkuXhZ
Z15ltaRXMUjF2NihXGXYfAkVGSkce2kALc0pX9hugoyQ+FXa6WddCJZ/zux7sczR
+SloDynbR1UssvcqKildNWYLUQOUHqIfi08kzDx53RWY5j+IL4lfdWIruggzoTOt
qQV7q7uHimFJDCWoE8nUXkvnQs70Q18w4MkM8cup1LBM+fbv9chohhoLDHDZYnXw
QXFhgRltU4IkNG2vf3Ig8z8SOHLN1F5oL3Fv3xyu1rBDv3srA5qWvSg5u1j+kttd
/JptWmhRqVe4Z38WTVHx+EI17NFz272ymQWVUUsLLc04PhBdeRkbF5ZlzXs4cbS8
e6tyCxEtrEB17PeIGsGAyk/H5tOY2kw1zDM2UEXEErnpFbuqqGTtWym4OGfVQb66
IOh0VmV4gEDi2SxAwsjkIcNtuhtu0XyBOGjHQiu17ZKod3qiSLv9UqWvxU+pCBAP
jlYJQZ8UMR3onrCI2gTWJS9thxj9NRKR20pPjw29TYuiUEexdxFh4q4LSs7MFVBU
Id6gqGVUZ+ONxvK9ahTASlOUukvsJqoxTekvF/CuQwaAzGqbRUPZEClMfyJdhqBt
y7F+DyDQOvrOD90U/u4WE+KjNxrPnH3AuL4SCUgRgvU2aCXb/rAtS+cWg8fEa/JU
Jawq66ISqvnrUyTQ64/BTzqgkhIWNVPp0w4IXPI79s4XjvSVm9BPjl5qEzQnM+Tz
m2R1YCtK1PZM7Q5H8gggfBpMWz272kShFn1Alfo0yjVZGeagSbtu/OvATX2HDnCE
TOqx3Bqam1oyS5QYfyApuLkFBx+usvPE7MxtdbPkzIzcMrYeuMNRe3iGUseYhNdI
c1/QeQEaPLBALzKBTceeQU5bOIahgd+0IDA857xVWq8MLs0PvfHz/lmnwgq6+rNy
vXht8SJEt03Q9WLUyPyXNBiU3rlv28XpNGBoz8rt1TboV8stGZgYotBQJqxlwAQT
htC3KBVk4wGc3kQqaxu4m9sbq409/p/rmSMOR3MhJjeIP6lwB6v0cPgKXgavkGEC
z0DHd4N4H8ChrM8hS11PR1F93JBaJhD1+Bs8nkNcQylXoOZYmO4uziBhy9mnySZF
95J0CIKxF9xwqjbXc6zd9Cxzf7ADnawbEvvwKbUNHD6GTjkTJzAADBcebfZYGSmX
0UOtHDezO96t1YBwTLYnTQG2DTULiPT1asOOzsJQiLOq+ywOCE+ftREI0Lw/pn8P
70PlY6pHsD7DBkC7y9tXQ6AkMTELNVUWbfM2TIj0wBot64KY5FEtqEoRSYXI/19F
TuySqW4lKZRLeCdwWPxHyLVMKqSVRwJuhK18OejoQDrIl/DeoqlRVFCAeFtS2IEq
mbsqs6eGW9crS59NKGD6fgk+pFPo0Tb9PmrqPZaWsypAlH0kj+yafVQabFWGyr9k
Qh9ePL3NzXAxxb67ECCfS0NIgUM5R8bsTELvmL9wShEhO5yvNEM2r0iH4AV4jTjw
JJLeRGLCwh21NPtOjBOqZjraNZykvRzfEram+KPYLuwPcugsaXaLkCUWeFkZsKuH
+mCKpjUh1404EkqumA8uCle4qoi13L4cUC0w3pntsz4U8/2jAfD4Pqpd2aZnr/Ok
52FICsoVAocRLpiosvYLCZx+9ZGcNdGCZ7cDWwz+gFipARKMI4OR7RARUz+TM2uh
eSVbPgcryEb4zBklj/1RxUfCU7fVNCtLzf2l3yVDUDE=
`protect END_PROTECTED
