library verilog;
use verilog.vl_types.all;
entity vry_divider is
    port(
        sclk            : in     vl_logic;
        rst_n           : in     vl_logic
    );
end vry_divider;
