LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY SENSOR_ENCODER IS
	PORT
	(
		nRST				: in std_logic;
		clk					: in std_logic;

		gen_en_sensor		: in std_logic;
		
		sensor_cycle		: in std_logic_vector(63 downto 0);
		encoder_1of4		: in std_logic_vector(15 downto 0);
		default_out			: in std_logic;
		sensor_valid_time	: in std_logic_vector(31 downto 0);
			
		gen_dy				: out std_logic;
		gen_encoder_A		: out std_logic;
		gen_encoder_B		: out std_logic;
			
		SPR_XRawCoor		: in std_logic_vector(63 downto 0)
		
	);
END ENTITY;
	
ARCHITECTURE BEHV OF SENSOR_ENCODER	IS

	signal gen_dy_cnt			: std_logic_vector(31 downto 0);  
	signal gen_encoder_cnt		: std_logic_vector(15 downto 0);		
	signal Pre_SPR_XRawCoor		: std_logic_vector(63 downto 0) := (others => '0');	
	signal trigger				: std_logic := '0';
	
BEGIN
--Sensor From TIME
--	process(clk, nRST)
--	begin
--		if(nRST = '0') then
--			gen_dy_cnt			<= (others => '0');
--		elsif(clk'event and clk = '1') then
--			if(gen_dy_cnt < x"7A120") then											   -- edge is 100us 
--				gen_dy_cnt 	<= gen_dy_cnt + 1;
--				gen_dy		<= not default_out; 
--			elsif(gen_dy_cnt >= x"7A120" and gen_dy_cnt < sensor_cycle) then	
--				gen_dy_cnt 	<= gen_dy_cnt + 1;
--				gen_dy		<= default_out; 		
--			else			
--				gen_dy_cnt 	<= (others => '0');
--				gen_dy		<= default_out; 
--			end if;	
--		end if;
--	end process;

--Sensor From Encoder
	process(clk, gen_en_sensor, nRST,default_out)
	begin
		if(clk'event and clk = '1') then
			if(nRST = '0') then
				gen_dy_cnt			<= (others => '0');
				Pre_SPR_XRawCoor 	<= SPR_XRawCoor;
				trigger				<= '0';
				gen_dy 				<= default_out;	
			else	
				if(SPR_XRawCoor - Pre_SPR_XRawCoor >= sensor_cycle) then
					Pre_SPR_XRawCoor	<= SPR_XRawCoor;
					trigger				<=  '1';
				end if;
			
				if(trigger = '1') then
					if(gen_dy_cnt < sensor_valid_time) then											   -- edge is 100us 
						gen_dy_cnt 	<= gen_dy_cnt + '1';
						gen_dy		<= not default_out; 
					else
						gen_dy_cnt 	<= (others => '0');
						gen_dy		<= default_out; 
						trigger		<= '0';
					end if;	
				
				end if;
			end if;
		end if;
	end process;

	process(clk, nRST)
	begin
		if(clk'event and clk = '1') then
			if(nRST = '0') then
				gen_encoder_A 		<= '0';
				gen_encoder_B 		<= '0';
				gen_encoder_cnt	<= (others => '0');
			else
				if(gen_encoder_cnt < encoder_1of4) then
					gen_encoder_cnt	<= gen_encoder_cnt + 1;
					gen_encoder_B		<= '1';
					gen_encoder_A		<= '0';
				elsif(gen_encoder_cnt >= encoder_1of4 and gen_encoder_cnt < encoder_1of4(14 downto 0) & '0') then
					gen_encoder_cnt	<= gen_encoder_cnt + 1;
					gen_encoder_B		<= '1';
					gen_encoder_A		<= '1';
				elsif(gen_encoder_cnt >= encoder_1of4(14 downto 0) & '0' and gen_encoder_cnt < encoder_1of4(14 downto 0) & '0' + encoder_1of4) then
					gen_encoder_cnt	<= gen_encoder_cnt + 1;
					gen_encoder_B		<= '0';
					gen_encoder_A		<= '1';
				elsif(gen_encoder_cnt >= encoder_1of4(14 downto 0) & '0' + encoder_1of4 and gen_encoder_cnt < encoder_1of4(13 downto 0) & '0' & '0') then
					gen_encoder_cnt	<= gen_encoder_cnt + 1;
					gen_encoder_B		<= '0';
					gen_encoder_A		<= '0';
				else
					gen_encoder_cnt	<= (others => '0');
					gen_encoder_B		<= '1';
					gen_encoder_A		<= '0';
				end if;
			end if;
		end if;
	end process;
	
END BEHV;