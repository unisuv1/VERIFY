`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LL/HTAJ1jH1ggv0TVuV3t6LGucjwv627eiTM84F390oGDM34bJnDxf8iHbtaYxRg
5TDT/owsw0ds+loDtH6/3DqOJbDwUfCNciIzPiDTACq+bXeFNNCi9SFwQLZWTSIh
JYhpT4I2ptzJhmqS52wR2vNDSoo6/Sg3PEL0sl4fFb5AcTrzLMwTLnmkfnvTn+iN
elQImVAgFHp9C4yO8ObBjVORurqhgRh8ZSOzguavu8Kcx+/kWjUMAPqQjCeRW7Fn
TDNEI4glbbnnaeYBVv122V4K9eArcw0hY9RGYokLRYDcVNQknbc3kNyabaB26k3O
j6rz+8ewAuU4ilqzrOAN/eBwBPcPzdh+jxv0ETqUxrPut4xTCS/Bh7sUOsCl+2t9
33MzMlay2F6SVVzJn+Si7fAGe1Ee4szztZw7iv5i5EiuF+gXy2y5TUDXMwtHRD4j
JN9n5SwrXAaZDjEFN4NpAkXC0ZI+VGzBw26s1bS6AZdql+zr9ZkijqSriSdce2Dc
pQw22KuFdndSCYWSaPMKoeGofy438rxKfKIuzKq0yKXPp+dPENRECMxnGhDtWnRR
dURjihU8WKiTBIF+cLL5DcGlWeL7tIulEGUK1DkPuGRjrxMJRreOB6sosRfGa2Ik
rnpSchtSXYtynL4jnA+PEufgC61xmUsK0JKQIcBk9vWDcyEqbgUnDMoQVuGnCDwi
rWcoO8UqFS8b8mLtZCQyvfD02vM4yn9X3w5wKg7XbKgWoj80jE6br0khzXlmJA8/
GkLcPHToiQgBhhTLhr5bOKK9Ibsmh1TcjneiawNcGAhBTDPuV28R+zO3mnlGXJro
BH2Cz5l8zfTBxUp7hYPK8YC4SsUB3RlhHBKPtsdyE+wBI4gqyT8MWkq8z/t01tmx
cfJMxcv42RpYu/UrEgrtC/2Eobd96s/Wf1xv0kMyP4IklvVeT4B1Ocdz8vDuKz3d
AcVis6NYnHkzakVk0LirgZp4X2cG9gwSvg1HUVE5PZ0TX2B3nFHy38DFhjQowSGI
fpZQCWFEzCals5YGV5+QOwuW4Wz0YI/BvMnYEz1xzfrPgbRyUip5E9nwfYRGDKcH
0bv1T2hpykjfii9q5z59AsirQARkHqSzClQetGsRoP0i22XfjEnKqGQseGWuX3kr
3VgFEcRsOVqKHWA70RFQ5jgMmnLvfCUbEQkzz57w0NBvEhjrBq/A9IIOnh54sOw6
lVXL+Hj/s3d9lqb+8qQ3mebUnTCQ3ol17QDB3JG+bGibEeToJ58N/WPdIdL3A08m
`protect END_PROTECTED
