`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Sq08fkn2PVULTrTSwGkJuXfSFQXP3IabscpexJJpMFd+7ZTzwXbZaEQbOCYIeVbv
inDFh3Tk7nBFgpkgBwVuw2CPnVqphmWlgcFScy76txm6SNPxf2Lt4ODu6BYo+UYB
mTJdBKQdq/ZADlCK6c/qyS2dl97K0zYHsPdPlMa1cmVC8dPsxvTkfU2apW/RzPul
BfA+ml9MeqLu3VLBEt0UYzyJZfSZtMyyaFeRwZm5x1NvrPcxcR/r9tarDVzU4Qox
wKQw0vZVBxzl3gt/+tauB2jmBXiS63KwoKa9WsRZHDOx+fWVzqXiIeeTaoUUXsCV
wD7Uq7nKsC65E3MeGxDnMSAfDJOSRM0OvnFLzmqrlBu0rNpY9DsxN9EPhzFlQydM
3P93b74JxQ9cFQMYjGzqzifDIe6JMZCNG0SkI0AwuKpROQrgdnwAtGgZAliLM2Rn
zQeK3ITLQcouIH/54/QoU4ruBbNmvdkSbnZ/7LV7+CddjceYWhZvTGPdXztDBGQa
PMHm7ojzGAnJrVKqBnEs3pL1KRT7c7mRv87dWBBi2wU4ZVfeQeDTaUeDF82t7hqh
Fn+eXBpGgc9I8ANIYRjU7PfdEbL42jqqDLoYWsRcyFc0IG7a9q1bjxdWaKdsVgH8
wkeX86cq4QjfQ1zdqB1aqsp+RmpM6iPIhNokxG4yHomcRfx8DTV5dhfUA0KVAU+x
HVx4ybp3CfkhQfIGVP1K3KZpJnM4BGvnP3jJopLTSiczrqJcIZxw8grZHreP7IS+
FLdZ43QBBW5SRtJdKKFUGoCjftYTqcK+rIGlaG/eAtRDJH5u8YnyKn2JHs94TJ1/
nlENAj5PBjkx9rdCKzIpUjrv7ElmBEAnnc90FkgO4+0GcMfKjJVd2EmOdMda0xEV
DPUNwTVyPJ6qAVLoIvar/SoejkbKucvPKbXpk4z5UpBplytxg5xptXk3vctTlng/
ogTE20w8SyBE0/J5x3mZGUMURiMMMTJdSRYWRvIv3BsHs8OjiY2H8XWwvtF3RKpK
DuwRH2jyc7/ffg/smMATh/P/iE1Lu1lO9//OGY1JTnOLpk5PsqdmH66kG8ytUwrZ
Ga5Q7/gqFEJPGUPr1qfdkeJ+ISGDGgOrvwuzphUhV1c58YDNWTxGI8a6PLVbHkC7
dJdqvLKKtq1gYEPKuhTP/+KCZdopjiWCMQMlITRhagbbO9LOAwnTt0pwLh9RPcY/
IN5JoKZbKS2v8nTQsWLjm0hbjGIYk1cjPS35ZX5VtOTMgyq12iSuSPoRWk5TON6U
5kDSm7Tjy3CNZzx2HgEQh/MRcvSEPQCTG1lJU0eRiptz1jooNp/VVM4gL85potwH
+lGPaCo4mOTWnzJPcE2CYKBLG5g7J4U54v13oxBRuHBe4QQN/D9dozCU5OoMGNjV
wa6xKOockg5sHpKWbhGDMzt7qu2XeGcq9vhpk721atuv/OrG8GG1uSVhGG9OvdaF
ANRMm6rInCYGWXAqZorKMjcuHcCIvTuy0JIgr7x36KDZoxR7ysquXHZXZPhOndp9
odpW1CSjVAvdtC+OyvM2HNNvnc4wlrAfXfhjxAo2PiQET5CB7GPyo0cTav6XdqyR
tKucqWOk6vpDAu9ufx7KzWyTtxmee4/gHfqa1OZ7sCugEC6fZzJBvjkKPr1Q3TE4
9MCYpzisB6n8x/w/P9KBsLN8u58T0fSnh4ayF7iv6b0Tn6sn4BsOioLlEpMMDpQT
/Z3HI6WXXmwNfPZM2MnEp2tnWmzjuqWrmwGzawqCH0/YlO6Twjz5kWmeyEu0Haqf
Uzxra2D91sORCbGQNSExodap5EgJxSwrrEu1VbtKuGEyQ/yKlPZs3iiWW+BoTS+h
1djc6QBoYkW5KdVMBRwAKzGUEd6T9D6KGrSGNr5XrTSOtiMMQ1c41YrzXjxS6aSz
27MnBmtbkKl1171niBwKzWr0EaMr5ItCNxAGAZG/IoI9/tLPcvZxUnK00SblsMKf
gvIOrs0gGG2e0SwSZqnWzldH56k9f6BIJOAspJU6IT+HFqea7dWAzlw/GoWuVgDL
mWq579Vt1DTjoet0HN6DYDTbnC2XsHUgBnqqqdfmL+8/gw3TqSZ/bISUcVQlvt9S
Xt1MdmBcfB07kWlYPaWIH17bcDnU1TDYx6JeQheKNlyCgXxoAWtI0eEgwpEG9UU/
yKRoevm+wIDMg3leBE/KFjSugNxbIA6JeDR4rWAhA/cvesSfyD2y/VzoqY9AQ615
/w55hbEC/us9pHOrYSzmiei2Z3cBADOQFt9ivjgDfYYGnbos/a8WyBGncLsILsOz
H6w5fuTeaB7spYjiipJ/TidcWh8ly8RChM1zMB8T5n9oPNlO/wMyEFVuMxkN+/CM
1ipSnrqiIH5KM/2oym4VL9Y27/fijGjyQO5oEqhrGxueHCglL9xFhq5IBr29L8CQ
cDe0XC6pDz9aCgJ/olVgTPj5nw+b4f8yeBClPjRbhwP4LyfUzCYCzzcxqlTW2F+o
iPC7HgDqyHim/jDCEyhL961ZcuKbv9uHTGnlAjsvCypNRWVo6tTGSxrmJIe5otfW
Sr8u9jBTWTVg+JGiJ1m/Kl2KhvamVo3jFO03JHxskU/sAwkA1CjdwW14ifKxZ5qE
mME7Uiv1vdpinRcL7qEcpwtnV64gA8IDLEIMbNHaXndz93jQjlmrl59GX+Q8NhAy
1tkN47lD8Xp9XoEQ+BdMNCLa8LTVHIGxoHMx9hxYxdLXrKRJdr0eqVxdSuC6PIq5
RtJKoaCpQP3ML2BuFzxQHLNHLMBBEEF5J6UmU8QHtDipX/PQXpzDE8KyLAkCyEbE
hCrkEuRaVTQZeqoQje9gPqbSNKkg95MifwncljD4DaShJS/0NsdodaPb/EHKe6Fy
5XqGrZ+/wHAxfk4Wo17R5P9aGkqcIbJ5CEWPnVjfHQx0pIWnobKMicYQUYDVyIAr
nfELaBYIjCdhoIEJNb4reFJAv4azDcAmlZfuaHqm+yLExqc4dISZPmHRjoPoDe8S
gkbkaKLm0msEUHe4aZbAm0SFMCGZL2ceTN8Iu293/OdgRyfiBXgB3GrsHgBfGji8
jkswTfQuFl2Hk4YGtrD2ywk91TH+WY48OYV1yBVGqmdkMvhImFuNi5X8Xw9jynJo
ZpggZJLulQL0teoAok2glNi6GFNYHec1BAnG+442tXJN/bWm4F6ww6sqwKJszQbH
WKujMIgWa4VKxNRzVA4sTs8QWPsQ/OM0nhcKPAGLOfrjChRXWZeNWg/IgFa5pROd
FAdxO+zsZZRjd6cDLe25v0sfXBhfDtDYrS59Kr9u6OZX1PjXTi5cAr3AqtHCzev1
Q3S37cxEEsWCSt4Nx9s5Rhej75BprRNZSIfoMtRb578rhVik2pbfqAlS/IPzpbSZ
ONfvfeeLhH50O9uP5IdgU0lG8xP0KDTH+OgLzbXcBGDXP7t6MPWf5zTQ5Bjb/MOX
tGP46iqIXoQ/1xPr+72V4Y4bNET5ZazuR5WOcZ5fYKnqAObBOmO+BPB3DbT1CGpx
WYKZzRLgvSs0p5SQRrVsPqCgvBGJp32/Awy9evwvLcUwNVuYAi/NoXH6YTgIlYXw
0/2/zEeRM2IzhJP2xm97Oen1zkeiX7I+oi9Z4pNQRg3Ycm02RruO8RzLVABLuyEH
yDT9vuZtSSWLZ7moeINYPWfsCINMy2pJ3O5PYJETnqGfUQ+TVFcri0Y/o2G45t5p
bMOuDxlS9d/25PAwpY1hFtecDUc2jUVIprV8fHjXU8AkjeQzWxzHpyfEydWoLilH
GumTG4CIPAee3/jTFUNcXpkMwh5qRJmlaBN1GPb2ea90wCUzHFGH2csnzA6aetj7
fbBsCcQqkqOGQRotjx8bkWdtHbSDi4ocIetohyBtFSxUEoeharXAwDQSNR1Xc0za
rLeVMqc/0coLPjW9ywVfm0SujPLTxrm0J5v+SjrTm6H8BVKoy3qlQ2Mv0zqJySb7
xwCZB3efPazr+MQOq8xEqEMO9UaRUwBiP5UiNAxyfPe3WpJiQbIqPdZpzJuhACih
ATfy8FVirzDzOfcXIdbzEM1Jv0fo6mt3A0iinPvH6Cgi+GVc1osyHXhfXJ4HpErj
Dz5BEkGjhZKEaKEKIj6ZsZTlPfuY+b444FOpAjgl4S/fDTokOm/fGl+3SA+xaVfq
n2lx6WpcTW9xNB3e8y0scbTOpPtkFIAV+6oNrgSiQCUx8PQ8CgyL6YT1FqnAi7/j
VOoZ3WBtoDSDH61ZyDq0OFtuiJL7V7pZWBNOULtpXBATy1O2Q1iaTWVHUax+qfT8
l8CJ6j6QWMX66tD72r7LDEsQkXkRFFNpOIvwcloD6lGVBUAH0+D3J7KUh+iJ4CUe
BELbclLEoSuEcKha5nMhMA==
`protect END_PROTECTED
