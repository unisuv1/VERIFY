library verilog;
use verilog.vl_types.all;
entity tb_vry_vhdl is
end tb_vry_vhdl;
