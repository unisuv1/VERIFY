`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
n1in3aXUfXCbIi333vCRQqmE6/yowgxrargBpB0LfEST0Q+cW91rGcjMwGPuzgli
+eCq7v1KsID+fmWCcbEfylEdRaJ/3o+2zinMw/BucMxGgtEiuNiRJBxHrUI5gt2r
wKqSeQLTFJnn7Dm3K6hu/W3uIi4Uv/683eBhxKoYrkZPXFSHI0Aoe+9TEUFA7rjs
s63mJYuW1nwOPXqmU29ICYU7cpQhGxbHKFXw9TaVlbBlVCvEsC3spAnBVrdDa865
aAagKQCDkazaoQCVWq3Dbl7A7dlZu5S6GnvfGB5KkZXIM+fg6zEX8NBOYDEregQx
O9dNWsrPVaDZCiAIjkoASOSe4reeqRxWi8Oui1dM9TMx6sIHHy7JUY3CV/AZUYn9
YdWaWzqFeONVJ8MzZpFsAyUXl7x0+vaQHBK+o9Tr9ZO2Y+mlPTc6/wbVQYpiV/we
YdSwJ/z9kWvS+YtmhTVF2CIiCVbeJg5xVZuuRKwS+1yAGv7B2rgVaoTlGu+FkYoq
EnmjWjpWS93xzWS9QrOyHGRg+KhK65rUnYActXqLQfQfCoLBvzWIq51XnRkx4J7z
kswsXe7RiK987tFMcFRR5hyL2wWRxMu7muOlCgTZCr3iNwpKPutsFoB9kHbG7bJp
hs1VeJOYQxVZWf2LfHfw4aOZdLrzfs/8iBPoMgHq1FNwKKc584bEeNcQJpNHZPEh
XyDNv85hF4a3o++jiZ69kWfHKJp+57WCtntitsaJyRy9OUr3jge3lgl1YCSQdIEw
13A8B9fwyKlrcww5zlBFLEuublfOHhRRlzuZ0JFdZ3jhBPgXkCMGVMKltW/56S5P
hMJFDBF47LNob8lEWU+N/te7MeglPpbZLtV6nC9hPB4Q52K+mciQ2mI/lQGmbt4E
p+TlGgDdg9KaW9OjJRXPYqwFjSxuflnK31lGKKhrUF04PEJ+fg+gupwS1GjfsaSb
j/QURcYVoBqFA2EggtZq8+PQrLPaBn5UwdxRPX0SufGts6XbjvThuH5jB7f/MfLb
KqHB+/fit90S+hS43viGTdrPTMYmL3LtQyvGdWMxRzeKVOnZz5VUpH7IW7inAGCv
XoA8rIzpXXiM8mNXBvH+mvlhloiLv5fNxXKf+yK3gKbFIzjrItRYUnVDAsg+cJ5+
vesGoyWkdDSHW1XjC62WP22gyPVpdeGNjc3nmAj4CRPZ1XRt6Hy8h+TrrlPNxQbJ
3fmQEGAQ06dneZJFtDau+0shhKo21VxEP39h9ITaz98lQ2rast4EKfSEU/hg2759
6tsAnJowMHqeqzU7r9rh0CsqF+Uf4LlhDNmm07iHWoH0/IW4U1q6VcA2LzT5wH3V
hKlnccQczA3PsUFZfsrigEwhKHgKvNyk5G+6tVu4zqf0kkuQhNAhx5kabU6FE29Q
G9CIcPqKlSDXX1TlWKFvlDEMX6fdwlf8r0LdvEc+xht6TkJSrf3DiU44CqrfPGeP
qL3WSk2bDnM6fALJq7whMmsJgs4ZwVakfmAgXV1e1pqK39tTCuITKwz5I83ikMf3
a1cMkeMhtl+DqKBvltsT/rGAFvzGfhtal42sX+xHTmyRlp67m+G8cYdMbfMDKne8
xt6Ncji6oc3VnK7i6fkyl4qLAEtdSm7wTke+zXuY3euCva2G2GTQk0UP8tRpBJzL
zluZWrY1J7e+nGARxsAYZYdfQjdjkkREt41Dl5NSpWwGbcANrRuN+GHrVj/1cXOR
gnKIE8yn1PwE8yOzdPoohL5n+Wvr8eLi0tqoEmNj1yTxVd1nTvrluc6zSZwLTZZg
5k48fgqHhrjddw3FI5KKkxuAsxEQIUZzBQm3yb8k3QfNsPKfEVvnbVW0KLobhUsv
YWTDlTECgeT771j4uZZkqQQjkVTWvHg/V5q25ORMvYn1MH9KTOUDLxUm8ghW1jN7
eUXD2YfVda9wBCjojs6niemeZ+2aS0bhxIAv5IfLCHy7JarEy1iiggy1r4zVjzJy
+XA8o/ic2qqwRAd455tP9bkxHhu6b6i11eEqC4e4lr5EhZbc/IHGonM0cFCmOPzW
lBXYDhlD5UWYHugry0QGo61q9N19HKH8fcDN9Gf5TOxLEzRwH2f6d0dD9Z0LF1ff
9XXdXqNbDg/tiBjR07ONcDpBwGGe4Ro5Bbn52ewc73eXnXp+tl18R86C01e3lqRQ
e9Go9H5w1PMP7inGfn6TnmsyCT517FjnYXSlM2ySkoIsOo5t97fEv1rRAaKWEgco
cVuuPA5fJluZAzSr/VpuB307j7DHwuooYXy8xaZyg9wEbQ0rK0EZN6rKiXsijH4H
5aRS98LdbPs5Rrl+h2XvwCQOyzKZwRsnlwa0dXHGfjDs5gYJAcDHYmymAKUq9bR4
Y8kkklMLhAF+lzJcU/f8muPJ1KdKp1/KHcLpE+LFP2PemFkeMxNbq1GjN9Xadil7
0Fcy+c2R06rMURbyKv4Mv6tfYsiLEnJF1b/XEOKbGHYe6iZEYC7UAehZJupxbKvV
Xn+dOZgWZN+DUlMDrP6+aE+SgAcDq7HyYR9iU6aBMyWFPj5w3ozYHT+kdT7ErCBy
dBaffrP9mh/JqjARXQnBYV8Lcei47WWY04AC+sUxvNJWKenEZoGWZDxroGfPCpsO
5lnPiW+et/5tIqrr1Q0vxsTlbn/Z+6gBU5cu6XJ/912H/Txk6vyLd5jLU4dsWbC+
svAjqJFEjjbtXemMWsrwlbx90XpKNkQjdQEl9dp4Czq6vp9Gc1A2kdFyOJo5NMtZ
LIGqRjRndU/CaQgaJgcOq5K9H0IoGA7Ilq0tqTm31cv0XaeUNF20iEqdYDMZ3H/k
/dOgMPew35atEih36HzuyimgGnNDju22Ujk3d8Ga6S5sDreE42E7iV1OcwfbhRjt
7k8h9u4wIEB98h0V42WSQyb6GXihUK301ka94RiUcBIliDOJvgJ7xym6lB8HjQYu
8gBeWcGRwZrA2ks+qKPsX8vwxjLZl2ynwbJneCr5DgL/qbEyEXUMEyCX3xIphiKU
ce4e6iGj7qENFOj9c9FU8bMrXA7LXc0BeqCxSJzRrJR5znL/XOa9GZz4vyLd1rX+
TczCAIRAAT3TFARjuCzhfFyhIv3v7OzIP1yh1tAyO/HWFZzoPfrY3WSRjZze150t
vfoLGzfRYi+lxQFKqPv3Y3HIiwessGjKyuYwoiX7iCra05E61+vr6L/mHLR2jc/h
m8sHbu83elfNHnjWb8rEAcj0HPSQ8p679we1g5eBh8VE7aoY6tFUxTlBg3xoBCET
CCI2Wt/6oLmvXZgBeSAsEbtwik84cmcb+dn3kH/CAMeKFM68wiXXA+ykZgArMMW2
bGvnmCLYPDMpOrrjSBNI/o0C/D8IzQMbGSQNwB9DYvR0GbeGLkx+aW+7+pHVWkEU
XaFGPDeexOtLZrg0cnOjsykPdmqiS4d8Jx+vwO9pKhm/I4E98x4cd32Sf/UJtAA9
j8R8qURMpGO81BUMbwg2zNtdpjQtDuenHyPYAs8GblwifJrlD0vAuk1GpRbn7Usv
YmnjfVtHqBmMIPqbFdRlPM3bZhROZ8Jkg83q+fzzzJsFYcNlVbsH7s9EyGJ3ry2o
VRIcLUnz5vxjkEcYwQPqfDkCouHqGBp8+H9XKRPAls7cYlhrVGP3+DyLH+Hn3WTm
Xrq3mhUWmWfsGJOgLbUTWNiZF0XKioq26B8QDxjH+m1I1AZqNPAfXN54w3pS+LPs
MVA7asZs4xj6cUopW+P4KPlJHXpp6uEtEF2lOtjzNUEc5jw5MUxl+x9BEWd6Ypia
An3FmmpWutia5EkT7QjnO3ly2SxaWkL8r8zpHDqvYJiBRLtcVehPD8jKsAn4hdZN
zE1PKavpuHRKKGKdzl5COWp8RE4+3bR3+fxqy0jZrEhaDgFUOL37eGTNvKIXiuyp
ZxXxeImRCU0zeagLPmcyczOpKhVsYVsfPCEkvWdsux8V8GCPfkHn0ar2eftFtq3c
tmwTIxKYny5zNWpyl61nBW6ys/uZ1U5rpdEDdElOQL2PsNp3+P3vKs89TwuC7+fo
xO1WbVaI1qt/550HEXak6/MKCBGj6sLZ2uQ8LW4sseyz78ju7yYJKZ3gu6oTfg3q
1RcI3tgocNR3iJ0L/rV/jQ6O7sO/KgItUrlZj13NxCHzuZ0qG4aOSxSYywg8MbdB
lDK1AjXVQ0hqYsq9AnLbArCY78b7bGXiut9Tu9BJWvb1KNNBeSfQbmPsqpGnQ8uR
51sFcffPuKu6RFH6/aqA+3Ng5EHB0N35zSBGmvABfAKyNxbih82xX5D4vDyb6hXT
DgJ5Nwu2aYulqX/ekMV9NmH69pZDDYTqLzjVmmdRvyoHvU781NPgIRF6U71E+GLa
IPRxguJhRcYvy6DS5LSoRj1acUNC0UfWUb17DJQdhVs=
`protect END_PROTECTED
