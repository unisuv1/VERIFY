`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
coq4C/CymSej3HEZrRh7/psBeKYs1+MOFMDSdKcYZhqeu0xBF3doc/HQk4nKx3k/
/18LtBcbKo8sMvk+XbxRhGEmm8n/gm7ZVkKLIL4nEcwQhq8OiBPB3WAkZOlOUkW0
r08URmuBuHBhryLuMwEJvw8pmSz42Y/Q24gaUj6rC6qDfbgLNBQogKbGcsk8s7Fo
`protect END_PROTECTED
