`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pH2JiPbadY1/Rw1H6TcQxfr0uzzPPvq6izp52fS33d6Vh+YGuTIsd42WyrDX7kfJ
SL+f3+zzA7FvA5zcmVbajL55HD7mOLqIchEKAdPU0wICl2eR+djfWJiQA/gGJChy
rW4FgNqnmHMs04UCT7YeONFqGswy+DRHXdH2CIfXZmiH/0N4p/8WjhdBE3e5QL4n
BysTL2hu4LgOLfgIgCuDrG7yPmUAoJsveBWHPfofxLBXhiAPAD90RPq6XxGGpt1R
FQTdOGIRK/iSoG9FPFxhc3oByJAMnBinqrROBfMoGlZ5jHtj4a7/u+f+0UqDddOv
rB3bUnwQo1/bDaAG43skhPM3HfMA9wvgM2HQwPbWjee2q3KzxXFp+G3hjN7YmJMz
HwZyr0fRH+NKaMwYS5TDXco0V6aSuEprA/q4Yj1IKEQTd2ImyL27pjSWMs7NOaSu
/kjmR7QqkC0iU2wlmP2nYRnRwx3CWwvECy76eGCg2Qtel1QTslXfTENpPcA1j/2Y
SeMpSsb330P8Q9mJjCVYvzLzbLRJnmbgWkesVpGeA0viIC33DWZFWNQIcLLW8bSS
nMtLnhyndGHGZ9Wa93YFl28vPgI0Af0GkwrrzVlratFFj4URYjE2QgE7qoCNv4Ud
dTbcZaJZ6Gyh4mGdnR02et1O+yGIBc7VX8a7Vihy1fdb9oCbuaFCSy6dnBzH5cT9
/8aPbg0QKHPYgaPTji0pdmgOBh+pR5UrJkigqxhhkTTnOJ4t6Nu1onAab1OTQSOn
lsqf4kNkhizPl0QA5mHUExDdnjD9ihegaFLTGuXU4gwJO+AZt7qRj5Ru2aHkrqLg
cmMYkUKK1SQTTv8oS3NPCDDHPMEpw2wHpYN6gvWLYUREpKOg2DC3MYCzIxR4PXyS
BGP6qr+m0YrH9tWhA43IKpwstvSM79mWS7AdQ7cOx/Tj3iFAgRs05h47gR45cjty
wxZ2j2/R8plHBCcQX7+eqekJMuXlYiBHSF0sIkD9Q3mehUoSsOT4wQnZ8r/hnERN
RGXn1c9qdpFOE/uZJ1vvuGIKmNnfwYuezd8mriPCtRz497ugkslANIQ6juLiuP2g
ZcUnnF8RmBn2oumu3kRgfiqTgvN13532GK7H7N8XmxSlW7Tt6OMWNQU7pKzfM0Ye
09ZPu2jZfAV0AJZsHzl1C2saa4RTO6d+alN/c1UPLcFuJrMOcHTsY2uzhvEtj1h3
/9INF60u3mbtMb4cxJdZ7x4PdjpiJEJw18Ynj50f2YrA+niPSyPUyeZ/KC4A82AO
9TZRL1WfMD+3q2YbXHvMVXPa6WJgUCXb4wDC/aScKfk5FHaJTw0YtPw4cCsLMhIP
CzYIX52N+mVUb6W/DaF2+XfpWhbHnig3/KmhXCIvchkMa+j+5MALk7pZIIYIPahc
JzpB5WnOy8cOdCoyNon7Q+qwuaUcV1w4Y9OCVtWYp4NJEOQWO4Jag6OwZNhMkF4R
IOLEcbZ10dSzr4GImuJQRNofy0n6K65AOZ8vrm4kCBaoM/ot8l33vaUEeQasZYXx
Xgu4yuhj060mpvQinK8MxkDhWPLKoROtOfUYs/kX9mCT14Ow+MtqPfcTnD6qg30p
Av4t5cdkTNZFVrJylIrNtuEbQfEcZc9VdAQ7MzEZs1+xXotT6rH8AU7J9+JqirLl
+G6Ep+U0KiJie5xy68vcMhWeHaTNKnESdoWAvtLxWUv9UTn/bJUveuakk0IsSy3M
3D4z6Ur3s7LMeNimqh+VoQpiO3e9BIk7UPXl6GZMILDlImtl957hqXIBD1GEQtiy
esvoJNGIVKEU9qBO2kPhEcX3sTqejyXvsdVlAIqDC7ENHLcu0r/3PQXbEPgQBrwJ
iWxBbh5R+BvrB1xcb2PQPVfqzjW/HOM4muAgQJgjcNseyeOMurutUWx1voVvogpd
d9RzPZUyhyFRWuhYoSAmNZ6047b2h6CCo33GsREdXSpYjio004LX058nwpIW+OMK
xumDrIn0Lz046EmbyuTXozOaYhGaxcaiFpRaFeGNEwdc6/xzzFrI/Rb4iutkNLg/
s6B7FmjMocxLi/03JBZwJPF8aNbfrAYJ7/tDUGRyMIY/eBaTjAgrq9XEti6Ct6iS
VglA0MjquyrQpLht583U//vi7ySIFsIs2rGiiDfOg5PMP67garkmrBIh78BzMoWn
r56UP9TmLtrr+U9NB7+w4iK0CYMC0QBjzITdoNaBboXx21XQKtRhlYPlaRB9Uxzk
S4frWTH+fxmW3B0cq3b1HBejn7+pEnLfOkFaceUDA1pM0mqdsiluAyXrhKbQ094g
fXH/7a8uK/Lf380WuX8Mj/lj4OucI+LpiNxcWdU2LPVuKFV7vfiHdqzkp95mT7Mn
z2lTTVzbKMEupGpfNbgeQ2HEpz6BS6gnr5dIHrBirEO2A/vXkNrqhTJPTAz94F+g
tr5iMVCY7M45xoCL+7/cxRyUWnn7JJ89yu+I7DnAwvSsZjivGbMyuN7O/5iOAHgC
bX3JYHmRynBorFi/THk7Idmg+cSfjfxaLa5MViKgL21YpxavP9qPsfX6CY1LQ0kk
tUyBpSw4nzZCC+zEe7iFLCwhXOxC96ABA2Q74QPZEkfmELURdOMCA9zCa5gXYxAs
0a+whe99DSw5x44ZljmmZbyLxl6YByqnaCZ5CFwrL3KoUTNtJ+SoGsM8pN4E3rXH
7e+8igp8gw0hjUkBD6CGwwKuGmyKm8C6DA6/ZKCnSM8P1KlAylDyClpMkKvddvxz
oaseP1Fq2Hh/RgxT77F+gjPr9hBVFmVJ0ne12covvza5Rz1NbN1eQRtGirnG/6GD
idv6w6o1upg7Z+5fPnK3PBsSMsJ+Zyk7UonbfI5E4D1oERE8QnqeCSPqUSbP+/4v
HpexQ5mTsAGe1iPouxY99vS5sOUF/mBVbf9NhBf53j+fyXf+ffyoYK/YWmJMfTL4
8oEQ5VGo+HvPpcdhOcy1JPmPPqojBwnYsa1m6l9jsuLfcVEfm03X7lgiERIxcdJ3
riX5b682TyUWkLP5NkFXjKWDaly+bHVxuC8MbLB0KXg3J/GhUzLxa8HpzfjsaOli
ePylKa57Bn/+8OzRSVPdowe5/woJlDIT5EqXFvWG6mel9350KAk2wBxxdxv7O1fx
0rYjuMdZO+kzfDyGWW8SMim1lhwMeBFLnPx75CaQKAHe2xwwHh/jQzb9bng+3vpf
/SjIB5aoWu/ru1d0bKakxSvX08WCC726S6WUohddE2H4Z2IwXHifG2E0WCJj9IB4
/sxEDgz4VcnUrXYOo6DKDT7GFI6DRJ3CkLyfa5D37YLHtsUUi5t7ZlJc7wqYtpzj
3RjbfXFtz8GiDnqgF3UjJIcyr7MDXOg/UmlH+lsygSDmDCJI27lrSBJZcKrakK51
rcrQzEU/jV1L76fmD5K0PWNoM9Npd8loZfztycUQyeWGJmYGcLt6Kxm2sSGuWp2N
4WsVvY06AvdQjye1eEOHjz70rj3DfPbm7I00qL57YFG8wl2/JDFfFryyi+k9ilgB
3/7a97XZGjEC2L0aULP9kH6QXQo1gJX3aIKmFhgctTUFd/v5UQ0uDS0GzvWRWVQA
5C5MCeYXjXfD4N6iNO4IJert4izf00GrMaWIX2K/sijQa/g0TuM6dozYghJU+zoQ
93Kv/mC7rsH5pEq0vkBdFuynC7PBi2xjZQhI9aT6zsD6mNFrMVqNqq6nfxquVZtk
lW6mcJ56Pxxw2OliIr+lT+j4HFNSJHaKgSEna1KkUtXhL2eq28wvrri322JyTBzx
F7TUhji3e7qvBQd1KqPkzIzyW98/xmctcInrePY0I9GuXR7J8YFLusfAtoMX8hjJ
gRAI+oKxUVZFOerXjODjATNo32D9/k8OLRVNZHrAN+4uI5N+Q9VLn1iRvlf3O99z
TnugHHUi8jUZVMMn4aKt/vssSNEaz+R9chhjk3qlp7k6bGlbnjL8IQ6/CzUmI1h5
OQokmaT3cwVU2e4rr5p7oQxUqOxNH7qIWeKl19N+s7AVkfdA8MIrsqk7X6jcpQli
AaUmwDlAsPglnIKhgPR1v/5Lzz6fkuFWEI68CsazjmSgz2PLvlZJ/D0CUTbwwb7k
cB0zYn3lS9n2Kr126P98Zb6nJn4DH8tWRXyLDWiYSRnbAlid5B1oTnEaxmV7qnf6
7erIlBgZybODIbtw3hF3n6oCKU4i0dux7DHP/V4AveIv9o76h+nXQUccAOasvyH4
g6KIpQYZDPl1Mrd1N8HZLMgOB2fEEedbmeTuk5pfKwx/5DUDlOHUDhjyIKoTOe/g
HvKNFjh1RMQDsr8mQwRQQlcOyjkthDBXTcFYitZDdC/ZEPnQRTlqDx2nY7ME5gek
2LNZRHlkkq0SuDORO413fA==
`protect END_PROTECTED
