`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VaFKJDEoVHsfnMYLZrUO3Haz59zfphC1jD31P+5I0dCw+388wIjS7nm2Px8cdLAB
KfjHBQeSQJh+1WsN094ZkCuX7OZYArIOelDrTT7giWtDy1moylM5t3BGL9GzTN5S
vMcViv3cW3uFgY6lfiORzaz/ATL/veR9aHE9O3GDIQx4JF4Jx91E35KO+Vulj85z
+s5GfubfKyx6CTew4D0ONNgtpItBwjqwTAaiQ8LlKrWdpn2QOy5oaN1/68kedzf+
txnEexZfv2iqssK80nofJVPrAE7CUPFtXOP9Bv4r51YcdYGVAFC02xqFVK3LhTOY
YS6cMlFlhKSUF4O1THs2ySLX2SE+vgSKoTgtgNyAxAbIqsGqgeE3RbDD5OB/6mZI
221l6Cxssii1o5Yxqz+4PMdY7GEz+UGxvIbqcdJptFdDcLFcl60VN7OUrDxsc2J7
u0OZOAfCoBs+iNaXVmEGvfVuTnkeqm/Y2/5SyEA+YcfYaqKHFLJ++uAeBxDXPEVB
9LDQaxdiBHr661U5PWS9zZIyHm3UsSyk58Cti+QibvQgWVOf413bFZXUc4tLATGs
AE9HIRc5jB1+rMO2xPVmpaLRRF6u4BBwD9js2SpnlCFQxBLsfGimHZAolE0RYTQ9
tzVG5M9GHxFpCHqqwz9kLW3slShRvcN+usqLYnm6rUAIRvzXq6KLskAsRGSkd617
n9NaTjOBvEkr9gRqdgvwE0uqmelrPcpORAWz5xMvwdePmzKvtWvJZNlxDJpmD71r
1gFK0oFf1KS2JSn8DW4E4+4Xu0p+BvDZey4vwgRRZTv/rJoryBbmQQ5dD05EMi2t
M8G56OQLwyp4zWguykjxOz985BIYqeIAq91cj9JSBN7Zp/p4nw751q6bkZ2tTf3M
npQjwPEJywnGESHoyOL51We4OPqsd+MpShTP7rY1J4iI3bYG7W4FB+0k803ED2YE
0jk8TRwAcKaMrgSmONuncV5gYUi4Tggmb9GcJfjofmB2TjYVQjUqDzHAgCWvqQ+H
A9ykvnuC48nouiANLan1IhlfDxr5KgKbfPswBnnDSvRT41zUrUxp6bn2u6vXVYZE
+Qefb35z1Z9uM/oCMc+a96rSRu8jJy8v36aC1Z2rJ2Ps7M+z19r2MEIHIgFI2nJ4
RGe2ORFij5NWYT5LGWsJFXCNggWjH2mZ7ZfSKljiEM0wNXyCAnDb3M19soK4hlIV
HvyQ/hqt9HdvwC8d3OBXE5/TjjTqC/kjopY4oJTIX/G0MJmtyIGGaMtNnwEkQRB4
+HEwD43gbV/q6V8DjK8sTuOXQK8HVjVtz93YZeVDPCXzrqv7IZ2557iZT11tMSbv
hbaWnyQxMvZ8FyrCei4NaxCtLvQe5pc3pte3PlUxEvoAAm1vo8tj9fK75q/pyo9k
qbsh93fu7MIOXAwDFf0+RPEFRYtWmKceLJj4Y7uM3jC7BA8un1Frq0nuEawFxbff
Vgos0TDFtofGkbl8TLK7mJZU1pY4wXZQ5i6fcPFqKhcOZiVKEfNeNeqOocUrTn1e
MRlXLE5FdUjesXJ4mMWQTSr9eqSkG0zcvVOfkllYHZHiPNmXLoRuxA0AXwNRpmCa
Z9Gb+WTWVBQhkdJGmlMYkLjbxGshilnAZNo8IooJmlxK1Dt8sCn1BXMb5J1QP+is
hRA5a6rdqCMi/oQGLJB2CTHOCYTv/xwAwD/WAHS7B54emrRtN0r3dEadJh3C+osE
bVRO7OJil1cmQgIJ0XuiXtevAdGNtoHTviblkEHBPdy89nqQGNZ/BfTV7Jwf0BRe
AB9+n4fPnZX6V9gAOO4ia00RRqJEsoErnY3QViwSEHuovZSnVw9XOW04kymgboTL
NqbPtxiI0MjXxe20l7nLXD+AmGVaWTayZ6fk5kmfn/0QIYpzIOU/EO99GOScbHv7
PIpGqNfq/fJYqoxd4nGCAJRkxySlgKRz+iXBK2TGIjB/TLTF5wabMtYFjbFP2aDR
62pUvPaFfOUpzL/C3noEFTQA9osG2nYeK7dk9HxHou8xDtJ6AwtCqb9Utfe9eaUx
7R3PLc2O/AOG3OxvAsKR1jq/iGtTs6ciy9YRjCB4kftpxTGDkCccLNqEzZTtTuce
M0Ahoj6LzQAqJJn401bwGseJBrXky0oeXsQNjpZ8bsCulS6f6qtq8xWLCOgp1TR3
05Q/72yEixG09oC+IXwlP+zecSWu4/Cp1QyKeJBgeIiW54iZ76DAIwVr/o19iIOV
C6vbxqaBEec6HALXizcpTkgflnsfGSrmbi6BhfvuYDIbsWqkCIj7xGfoYsESkvt5
hwBAXJbCnxNINe6StspfBqtyYHRbYLihTFUZe4OcO+CHwCpXXUuhxew6dkizERHw
HowGr2s7kth6YmhQLameALLX0U5UHrrMFTLSs2Z+B4gRUmWRJXZvtE0b90Qld3D8
1uf5v1jU7stQfFP9hnuv7mUsTgQVcuU1OspwzdgwyL7Du5uKAF4K1VQ+1rtaKit4
XsAsrr5ReaB08rCpNCQSHH5VUw//sgw8I2GNNDAG9FfRaFASBC83HbLEd3iyWIfq
wo10c77QKmDw7pu1GNqHTLqXGsh5OpuLfPLTBTMV3920pg6f1r0OZKAtb1u62QO4
UVvZ3Ky7HdXfEicQ2BOIMq5XkGK/LKUzZSt7j3fiFDOIMdHvCuc7ICOYSia+CQ2u
Sm3xg4XLoVUcb/pmm79hbh0hXb2zb6koF+FDYAT1LkC8sZ2LGiNs/7sev2Rk5Rgv
MEpC5/c7qolsJtJddZGEx5cEUm/x26uAXLZZa59373LZYTKn4r2gm1QzjHVUbLlq
jBoMBNFzOdsSSAlj7/+KVUQTGp9oQ+8eQ1cUz0fJrg8JICAuPpJ49jK4rgNPa5Hq
WZMn+Cjx8zH+8TYiH66Yk3TsddEcaYdhVmBFCSwWjBifrQdkXFKS6tbDMRqqX0ge
+lpJ8/UdrQ8OZaESjLhtnn4l+uayfDy6yfqObnD8nT9iLY/UjUJQvDNwpq/nrhnr
8KaDr/vbD73wdFSTjPdmww2FkDfhXT4rjFzQWxajNCVdlfmNeJZEzQGaNvNPlgza
+9tbSEgqduSMcowifHan3pN5bIfo8MQ6+1ssBbdRBctSmY7NxLSpQu7tL109zSS9
tXcjD6lWEqZGZ4NaNGpPTrgJOqKG/OBqKzMzSe82TINfEBJZcCB6Wn04YWRoafUA
CgbVVI71FOBbeWseLsbx11QAHyr5bbpkgLuN1E8ciPileoKx4gZhryifnSe301qQ
xqaHOPNTSJOYKjuGZeVyTGYTAnycVIp5tNrDAmcjdWsUwOuWiNngrwJkok9CfM31
C1gRbEPwWWjDnXEMtEEWV8QrgCK32QXISizfqBLOaGtgLTKs2/YNNgDFSlt5HP0z
GtfdU2u1cjx42CwuVGaX1ify70jNmbiS7hWo42eAFKnVkeY17P/VsOvH0OmoV5uO
TIiOqpmJ4CXZgKX571TykZkN96Z5R5VO73SQDYkAwe+tsdh9pBFRVOPSMNhze29Q
QusdZVah5SjDkzL8171JOig7PG91t0e12Y3di2/F66UBq3vMa/e3KZiy1DFHU192
KoA5+OlqJymb4zjLYbZaX3dM3tLLlG0SRH5O6gV4MfldI0zsJofwOV3Pc+WVGycX
N/KJlNe3hhXU0B2M4tRUUUMKxabXLk8SzbPlCMq6ddNCBMAQdWlKqf5/wH5sm22k
EOVz3E+90IPSPS+VktnDISOfvQbN4Q4XL1P/cqG/gKkPpPhyBB6xk2+a7BSSDnIU
HF8c04kFllvAXa4zvBqVjcqOoUyD65+LrrdWjs0G8OvjZZB9pdaoQ6ld+i79UW4P
6+6oDbGsroEmfjWCztp4JJ/1V41Wh8u5V+Nmr1914usEnLdQRneJDT1eC/zh/bG8
BY4RFUjKmSdsMOHB0oNgJIW/WBc1UJlakae+f/k9GKR+wpeBB3oLAce4UU0q3lXq
RO52EjcOMCTjHvNs9RmnWWJ48NqE+XRGXMFJMH6p4lVYeEliRoaMv0KHaTXY7ym0
AlSA0pXoi78wBV02FU7H+5jTPq3N4gQEB2yDXZH0xUprL8j/XUKmkRHaUgMvjAwr
YKuOi+0lcXTwupIPQI9/ojAtEsRewgH18rmPUca+bjhpF256Y6tEtfwbg0hqViwW
vpCdgEnQmF6LSONwQS7KWeAhkxVoSdJP3FH/RbKdSW0M39aWf6UMMZUwXOmZZxi2
3m9ga3gZnHMdrH7KETOGAt/P9A5LOd5yNvxT8BgdECz5TTjl1hpM3sQA0e2nQ5wm
UG1InQgqN4bfVPAHzdIBgsiY4TnbHiEtWuQjNZPEtu/ckVsaQj136k0kpJSuWefx
HeXpsqUtd92my1WeYdwbp+FbsAsuSrn9YOtq+p8pD98h+Cxm0wGRMn2QfUYhcS90
QPhH55HZSdSo6btJEdR3oeirGtn8CHUi9oXCYhcI1dvW4QjCCbvtaU6kKLuLvDSP
8a2eI0vY7NPj7l2/jhyf5zWIkqY8rmDseNqdpqook4y0UAJtEaeNHyedb29wqqcQ
J9hV13ZfhRfHgTAdekkCsgmqGEzmsGYkoDi0ZfzGsf1q0y385DruBUHQ78p32wO7
3pc/NL3hznYXWMPbibBjjXeUFXDCIb5F4q/Kpk2og4xTMZIFuocacOS8r72bimD/
MhrBZyEqNcKvbLel0dMvzcirIwj9LvDmAd+l3XaD871UMXn2YV1WeakJqF5D6OhD
mnWvUizzNEv8p6ZZVyQzerVos1Mat9+PUky3Qw9LaN02TD0mnLDyaHroOyjY5nAK
tV74/JbardCcPNd/KVItjpl5QYXU9PLD1s54SiyzqCAfDaZkcnqYHap4c3I6zh4F
pYwBgLyMjGRrkId1EwGPYz3ZmtIEoIndeha/Kc6mJ9nQhd5CQFiihTeMJCjXmWm0
+m/OrbtRv04GXFwAYEyUJJLlAS67n/nnE6P9AZub1Orp6/hyfh0iMmv9CRGx6FGe
5KUxX7kbv+X7zgtdl4XH9UvCXDeLizkvFA6IetP62JQuOgbDAasDwlqPiK+hgzxF
HO335AChJODtj67vENDwvGwhUuC/z7Qx31Gk/vMivbsu78TsmIWMIFC+P4Sub3KW
LHz6pa/aA3uvvoqIIGkAFCg3GFslIiS9AVV+d5/AsR4phHm6dsSSTds8CYLQYVPs
9ciflD4Hb6U/OtVBrrA9BWu01Fv+6kwJR7tvbRy4DYcIwOfHt08MhbPMyjiVe8RY
OLg8vIhTIR8yGiJeVDbVt2VKdLqZjueQugmgNDlBE50c7e3Mj4+MDqmuNaGTfWQ4
43M78f7Icgean1RGDSTcQjpdyslNCfZxpSNKN22/ry+PXvmRre0NzbX7KI32VLtX
oV0acv0E5/sdjiTOyZz3ZK4vfop9VT+EFZT42VV0Zcgaz/o1aaZjSbF2D1xXG9CX
Ao56UoO59LWJeKCXlcyBed3hPwOMJRraCm/MWJNEv5CC6BEHkXuQsep8okPRyseM
hBJ6KjU7XZK8FdGW+85oipZ6kGk7FK/dz4d9/7O+1AEXt7ndVhBAILHsQXmLAxqJ
GoGU2R3pd1LcXhpoenScQw+U0LkC6RYvRNzICHCrRayK07xCiYfgEgsOnAW/yWW3
8FF/wKQDC85tq6Gh8oWQMafRNEoHVaReQxiaJSt5Op0guRDwaqY9ZzfCRiZgYyUJ
CX3c1oMGJmXTqFa53+/33bXf3dhBWAOReGZKJW44i9GjsYSaVw5Nk3G8Gqzh921u
nhJRIIEIHYwMgNsJomNAzxLvmJRN94JlfILkF2WJjY2/gCiMHx6zcHrZPaEMNkdg
V7CmQCOuKVMnFAQ0WP1n0YBCDUgq7oPmunD1riPsqMo65SN6ZhaAsd/rlQ0zlaJc
E42o3g5/FS/0RD1LuRcYGJYrDRhV9ozpIlI4FGpyuGv6vWMyde54Fezl2z5wx6Wl
sDbtOezTDG57kLIiFvNE7P8ObTL6xas60jS6LvMs4TA4/49/qVQHWYz99wXQddzN
W4QodV2NHp3QNEEZZ7/7mn7k/ZgiKQ0IWploL5X+brl6nd7ksRdSsPwT9NA2nP0A
BYkOXbipgZ2T+vtz16o95AUFy/9Ak3e5464Xm6SIGWvxESoOwg6OuSKNpHZg7Ba5
kr8pLOOa/cYjcwUgmwcAfaMyxwWD6wykpmbIHaQdGouEpZyE7JdHVFkxRrgJTAdg
dQsbUqzlMhpkzhVGaK01ZzBu7JwKLQriePmWrNoiqXv2SlzpWdVFSfDBLfss7WCA
exLWwh5BbDd9jXK6E6Tb5Xf89BcFUdShLBn6bzGe2EZAu/uREngcKWVf6IItD4Qd
8eogMICBLTt6ACrFoDr2hNJOVDMfm359xspqzzCJPGQSKsej8I4fwIzLQHsX8mvp
wR+EqQWzlyEwS7xH9FEGLOxcHEXF9epf+BvWHGhDGVfjkqd/Ct2N/4IXYYSanLrL
NDkPyoYB9gtYNge7KqqciJLZwTHxfbWBRMFN66wzDygxkIEeKXnKeJZzIbAqdYtf
78iN4OzV956H3AdSQ3OkVCw7rZzglj7t2W0uKHrXL1g34/3oFBfxm6aeKmE4VhC3
64+Pke8WZZKWL8vJ4J/Ob8GpiDXsTvGviOflzd7qy4Fj9+e+zKGfOhDkxwtlE6eV
OXd74284PKAG02RBdXOaDYB+r/b+V47dviLbwIB0dp8B3gBeUGOhRlJKvu6bST5v
+PZjXhxmkEp43rl9PC4AmCAazcMV8hO2i7UaTZEJz10RT7D1mCNuGM+teD8n83ql
gK/DS7Fn9XPhJi2HTlPBA8hKtls0ACM2zfVZKIES5+nTZ1aFM2IAcXpNHR0Z58Ku
8DHViYQ7qQJLEvJxs80vhz6DaNfi0UzYyLsv77TaMslyTb/iJ0gkqpmRWIBY1iXe
xaeWV8rtNme8K3Z6WSMx5ZjjzwfTtdzoeLv1d8V4YJ9qaojnES3vmFl3rGCTqsLH
32iSukDG6Qayp1Gjox3w+8S0i0UxlTdTSiBV5QlBU7ED7bxoNgwTWqTSoiXoho8u
BiTLH/wFPF4K1LGgZe5bgx+tgdgDhaOEt90SNUXBLBhkb5za1tvWFq5qoaN8I32M
OxBTnp6jRL84EX61+Ygpi7MGlumD6IlXbZllYcvPl23lY7nIkFKBveZGuPcVjI3l
tshQKEDGvUzF54NJQ9ECrsfU2Bl/QQHeEUMmm5apKMMgDCloG7FI+MvkG2d9Wk5j
Ps1HjagdpXEO/CrWgST7vfGSPhPkZvhokXMvggRfRCrX7dADN00xZwNK0HjNSFcQ
Ov9806pxYAVB9CxSp6B0ZD2BQLJrzwssMDtgYl5K7iRl6NhyGIKd2RiYosmVYayo
Xa3Ksp1Q9Sh785C11k+ufYN9LBJ2yk/5GvAmMDmRIJbDTrbdsMhs2oBeasFHgVhs
FNfh2NLCjkhTsKf/psgYh1iQsK9lX+Ac699DlHQXUlrRd+qqF3RHUgVndhNPSMqc
56Z1ZXwXJIZc8/pX/8pLktpj0gzXmH0iVgOCr41WgjmJLI3fSmfpxcxP174oMBlN
j69XBJuo9InnMhxH4V9dKUxUqsyk5xFqUUAymd0V5EvUQZdRRc7W0dw5XzTngDkc
N8/2BxlivjBwgknDNdYS4E6ksFuvbsLtDIIodjNZcJeMxxH1PBGagyk6nG7xtswB
5upGoRWyV3JMpTGUoBUvf1ajKK1Sv4jS4USKnOEzxP/WQfmiW9+n04ba10CYNDo/
CpRQ+9rWyUuwZzrz9SmmmWifEEmLLhoCF3P192v9Y6hxgyHRS4QCoMPxr8ivjR1w
6G3xmFxXpu75DLNdihfyafwcs70d9DVUydYcI9a60QsbOQ4xKaeMeGMz99x1Hl4k
XLCIPAmD83ERMvQUzhnSibLVRBWiNJbk0yuvOEfyjtaP8doX+D2b1lp4h3mmLG+z
uKXFKtCa9fuXMn3iFa1Vg4wZ/P8p4uvxuy2VgyclUNTVG6K6XT7E12TopHNoSjbq
JIvmk7rGOkCFvjEe3t+gBW3ltHwcKFy8y/vIGuEU4QrhpY+f38FvaKS0uGh7TiH6
a/D2J3Yygy/FQcNI3KDMavF+/9A5bOawqZKo5EAfKfqwrN/mzYXiXNBft1vX/cj0
b4sJ2NsPLw6YzEENmDPRjtwM4W7Mbb4ccfWV3JM+PHqmmSJbSIpjWeYEluIk0eca
Jw5rdAkws+0J6367kkYpUOzl4DzPdH2JPmwUy0RN+M975hgP5VAt33mBZQkDr4B4
qJzUuMlwqIG+pspLuSIgziV94QEYD4vLorMMQjeu/JAasg6EIgR1RWgxCxE9vkyP
0SdcEleh0W1mTzAuqYpOvgi+i+fL7M1fMG5giNYJCBy6DHG9byvEtmtFWHNl8K11
A/2FQJ2ckzsUopa3YFR2Rk7rvz82Fqy71txo/WxhyAD/eTnx6pJuLZ+sGg601xv5
WIhla31lYQyAp8u6YlqJ0O0jsQuC4j89bYioVQPSdP1VsRF5e4nV+SrRx3H9ULvT
6P4MiHWFAJscEfM+1o6+MfkSDtUhgh+A/3NZIckgU6YV4oa2MYpQpVJrJH5m10BR
eTVBOgiT0CDh9HUelf8sCIrqeJ7eEtkarufc+tbNDKYq+i2t1qoUif16S+3kltOO
9kTBAT53z3Jk/ULJdePFYfSdFuikutWaqniJ38L/K8YEaPn4sMXVQwUXW+Ah5B1J
ZXZc2hmD9b0augTKF77yFP4NnUiuvPBY0e0jTHEKFXwGIq8+Ep0QLSLneKUvG8B0
B36yh7+l1yp1IPLqpWx63tS3B6FipXs1MJsSyARu3ASoOSeKTqWh+rqn10aubF8d
rQf7Fk131r9+nHfeS6BscLUi8IF3e5auxoDTNzVsypLEBHu7Dd70MTGI3Irt1PSI
mFu08TsS24+RZSXcCyTrI+WrlLyEFOnEV5cBsev3/wIxIwl3jRdAfe5tVdmKednw
k/AwAeOtwypR6qEuw9C15/p2PUHd6fQm74qOiVK9Q89FgZjH3JBeGVBy9cARqpED
x3TYwWH7JvOWld7tgNWB2pjt2f6c1MbnTSvkE+bO/v5OoM1gBV/wZnEqOv9jydyG
l1P4vmj0cZPiESuBmL49FGwHmaq3N9JKMA7eOfa75VHJICM6W78nOIMna4bcx8gq
hm/LPXap9q0zo9kQ6h/daImjX1tZ8UOQizcOEKN5arOMmW3Xk8gSIDgjCxg/4Zk8
x9GlE1tHc8PDmg0a0ZM4TplfNT/GwJ1dA2PuiL81CS1Rthd8NqAmE3Jo8L+HXySt
FhLHAPAgDhrcMQoZh7dE4Ehc9JeDEzS0GOKaZJH63hRg5IzpvgqVvBqewDQuuqpr
4uxFvFX4vTQT064B1hPJ+nuJrWZLKZMD2DhTIl7CpM7OfXVLcp4/D/pOqNbMJFvU
RWN2pYfVQM2YxXJu/qrYnEm2xZ9h0bhIjgXZoyyrLnRm7qG+qA+MMl78W2ZEm+jJ
gH7lN3sfcr0k55YkdfKlfHMsScwfasfC6caGEwlSbGTpF10xkEO4U5a8CFjeKqWY
kV0QpStXHiIPUXUMZ3qv03AnRvkBGUVmD9sTQ4a0pXZd2AMwoBOSTV9+TiOf1czt
b+5CMiaD9oOlzOIwzPivlzq/Xx9FnHXWLOcVdZmuU3ixNAV62bO7iFBAZGY1nKcO
Lz3KKnGh16afqSX599iJd6GLfVsMHoloWj1XWj5re//k57xbm3sTto/Dx8TDMzuB
74wHqyDbd8ArAsrD0w8jBvozIzYFsXjuN/h2EOMZ68NsXZ3we+TnQgZLiTfgbcCC
d+Fz/AxUreLzY4wZZYJ9upLZ2OCvZJ4FDPtYJirZJMhBiLH71bUXOMW7hp5juI+9
K1AMt0RooaXpg7Eexx+vfcqGhmoDaCdcq+oXaZamI3UO7L59RUiFvoyQSUUjJ605
7vHfvpAeposrl6ThmQASgbCnhrfg0Q0tYJAYnaTyg9RMEeZR7/FHkbh5S2ke+feL
quQe6S/vwwX1bHY9AatAAMgK5kOkdV5vDXSyHaBd27f+FPldb8B72viH7ISFVdvi
dgw/KrULBiBR5DeKACYso/BAkXCzmkgNkiH2uM7mk0xDUZ9zMoe56RDDJFuLc9yd
bwcmJWBiWU30PhHvwVHUmpmgH8xF4kmLqk8wmzPQtFtCxEtlLMhQ8pgPLC27V1KR
Os/Aq8PFiruZADSW2XtpRq5gS3c4c4gauqzbSZFwheQGrDLUdG9jFrVfeRsLqbMD
igh8DVLcUUJXiBMwxyXhAoV7e+j7t07To96PQjQ5n3kSQ0sX2OSm5TSerbkzVcgR
taHRDKSdgEF7dMuu1tzT+Ar5+OnM399X9KLrCWmMLoV7hZ8odrquzbrhlF6YTwOw
5XPVgFEp9ifR2YAIO8lWPRXznyXe6lZwTjyFhy3Xa5o3HAOsXyQS4GUAGnZTlExZ
wCTNtSiQ+WdRC6t0FRziYETUdoVoh21zBU2Bumcg6H3nMstPEsP4VJwKgJOMb/fz
EAqOKlBGxMDig8esHhPWofpDZUeljuzdN+0ULFgkWxKTXP14ZRZfjGJIgN5II2De
4FFEBGUsjkyZv/ZtaqpYBe3EaZJdD6S2u/36/amGiRSrH6bXNMwCi3pK8xX0Eg9H
PfhuN80wI55Vbp+XPa0RaUwKgaI219XllZUm/xDjVRoTNalkzoWi5hHcsEhCBIhm
zOFw5URhX9V49+ZJ6x/+frmptNONsuDOoxvmF7W1ewUMkF9U3dWkpuxYpGKEKDuK
F7NsTmtSuJOvOLuNIYx7bA2eZoJmMT3H7nm0gnY3mdCQJBdM1qs66XBoHDlj+x/b
+zwM1kWzYOn0pfxgaL5YdLG//pPTxYv1pSBpteuVWX7RqqNuLZnbp/MQSrNTASP1
5CPDKLIqa7fyVAG008lmtnuTQf+L9Vhu0810EBFsVDy6rwDpLuaMm1X9GjYVBnXJ
deUypXqY1rzWnv0YbGDlefeytx5JKZn4uEJLOhzBGd34uN39SBZpBhZHRjJUmhof
Tr4qPX5D1dGH4xVGQI2YtFPLSZ3SxnaSENzS/8JKvMFp4SXiwjGzKCwPubuu6ts5
GSvi3OXRAPd6QQDXhPP6baCiRptcaaGFyyglqigILpTa+nzGDJnOY29stIkvBq6c
wZoA3aSnrEZmyc8k3lZiBVvPV30s0jK2L/3T2L6zXaig7e6R7ghksasv8aRVNWai
l9b4APhcwu3soyab/baWbfkz5dCE64f/WC5TQeG7fj7Z1u5cbwUW0zlGLPkzp6dI
oyUR2n0StN2vWttT9wlP5COOLEqQbB/TcCcBl5IdvO7kpQxiZohVVzOc//wslad7
ptesFKUfgSDlyW2Ej42JpPHlnBUWyOiXG2bVuf5/8ZAhe+r+0AoW/6llvvp2Q4Zg
jk2G8RFJGPTyJVKgPZEu02/UoxllnCNJPiyvBJxvBQ67QjlTeFyxig2pJ47cSqVf
+1YjGE+dXUxNGliZ3kftrXAWhE53QpW9HfeQPBJqLWpotFBnJo5K7PMo2HGJ7Ptq
RbH0Ky4EnaHolwmtMYxkk4vRepU7CvaV83RTkEXuwMzrrWUCyUdZA64TL+RNv4xV
d3c3m42aqxadhCkbF41wwfoQLnfxDTLulJdGYnmDKZjslojAzTJreyMBfvDudCNz
hTFYVtRH8ka8YDO77x6pFXPR5btwwa2CV+eAbC145voKd1EbgqqtpMZbDKM582gO
Sw9Pf+XGfVGIZtophzd0kdhrblGtlambL1O7GPHKGBhdLiTa6uSEzuPDXzb5yQsl
1LC89D+IRRPSvoLwAw/jK3Eha+ZaKWCyRdIJBeBIX0B/qw/DMTKlhHwmKt8WhrpS
5tcAAWQnc3Lo5QGuvJZoKqbwA8KxnRy1tfwI+tANEWQ+kH8t7UDXMRn7i2Wn+GqE
zANxBNk0CAoMHKjoCvSgGDnRvpzxzkuO41aL7Tt29cMVSoYYwR6FrYvmog64atbI
y2bjrOi6r9hracQascc5zjaeVm5TNZCtADgch1d6xa9bVD+lUEFBboyKsbmHmEz+
E5JHN6H4640hIEvXPdkLkdGypFvkMM71CAV/qAzmuIoSkIApUgHgEhDLnxxWsfbg
jzIbhqDUDmce9gr/bKGzVY+TC9OeIUTFW6CFExu8hSADeq8POqQKt9aWHK0mfgXi
YysmiNmxZbvvUT/zefodfS64B3OH1+VmDBuudyPXTBU1J5XwEZWFh5KzIn3pxxlb
7lOi/q6Z8qFttEtxloixYQumT+ze5DoGWwrbvj6D5o4+YN9DSmFCdeeDey3vtZ7z
nhwjKTk1R6VEI34qIssLQxrcGe9P41MhrqbmxX7aurMGH0fFXlBH9Tzn+qyvumli
6SH4uiEctRmEGclOvAeX2y6b3aQ24CANKk4fQgZHs3/1dAjLzUk+CXuU045G11ki
7gMoXu8p8hteltuH7xqXyKou1fuWFm2E8y2jShZHAAYLFb1V+LeJpTqu8oLsETN1
IN2OBM9FM5yB+R2hJkvQZftja4p71WS6dfsldxCbPGTajiS+1Lo3zqg6eIrGVAHj
DR+DtdlpVfVOw5jw8e6S5cUnTREO8whOMDItozgqFwgMHvIegITd86mFUuA6vZtZ
JThu9ZMoMTV2urRrS6uPUBijoOIoYh2Mja1ExRFgJblw3CJABQuTFpG38PGU5Nu0
erzkqiM7+4Ut34eSBdkBuAOUIn9ow7jBSLGwQ3yljUufjCcbgqq87Ew+5DiAv43B
gksCqOezNWtCIPzhvcPN36d6HiaSIqSeG6knOF90BtjzDdjAlTfeHLHomx+yI1i6
0SPho8XNnURkpOE/5kNFNpT1HYaIAEG5FXatlV8/BlEfpihshBjF8Oony4A0Ww0y
1b5NXX6zS2nvnpJ16InopqxeCBhDp8y+gpltLhlY7ktozXZ86+3dynZTreljQrmz
2C00MnRnIwXPyKz1fqMfc9QTI4ZmYfj4EwrzSHH7P9ghO6K9rJ/nfXabsm7syQTM
cutKQpGSAYtLsc8CJbz4H3p6xw/Z+W8Gkcz0Ks2C7BIMnv4bk0O3tg0gC3/56NhX
+gKMaA0i/o16rvUcPycEXdom96KAzRRg+kec3B3GLihbfcbmD3VUtw/HUkCgE+yb
CCrrky6VkNJs+OknFtf/D5l7+ng69p3ZMST23qmRayRTx09DQR/3znpw5aucGjo5
GJzeZp7DEYMAJWrnQBNVrUk8Ol9gXF2d7EfhJQGrcNeNFmdYGPLPdFAT0fSo9PNx
E+7dNedPWNARWl7eya9LKJSKS5WL8lQKw3BnKJS8RtUKWtqQ156b0FaXspSPwXo0
5/dP9wveFGTl3AKYPWLID/j3ohe4KtbiDQ9IONdFBU9OznQmxC3ObyMxrGRRpKLs
D7Ivdk/qUKdCbS44deMRkQCJGWc3xCwxc6L1GLm+P6HAzBBh72uTXPk4exqgpxXO
Aki3iGXZelpCylN4GdKhrwwrOcyf1Fqgx6JocxzQ9zCVRsD847bzgpsQHJrC63aV
RRoX4CR0h/ewtTvgNeBpSEQyonJIuiuXc1n1EhOgSl4VPMLxe2Wi8zM8JoCl2F/f
Ro3yQ/BXqJWsPyf2N4MRlY/eWJbauPdsMHfM0/3az4vG6jJ0RXdAzrUjy1GBqG0r
KPJO1AQTBWEnACDkYdrCZ54ussDQy1GN0em30pE95On+d1kCoIrTe0IqqSR0iRqS
HxCn1uYBJkpYX2U8c6AC7OcGtX8/xdY1bJf8YCliMP+Z07aQWyxIG3fHeyQ2dhuc
TyblvrUMdVLcF5ZLA3XdIWN7FMrcswpda6eN2NxS87HaMmJ6xWaj+4qMovW6GnP7
mj3TrcOUJzLIftcJe+rFSmhi9njyc1sLuqRhiAwgTeZ/pm53xV/W08dIW+Pi/eIW
3VJym0gKG9lYukDVxNnfP46EZd+FLRo2pS8bXIYFJehXVMgBNDcnnUqYqDQQ2RNO
hU0mJmKUhdUD0DQWkaolEx6vRB8+osY29naX9DYK7+N+CcQXeZ3spLvRDy6coJrc
J3jsCZ7UbmVXhCQRiqKo1ikfmWo2bN2IyvAmDk904FkGDnA3nfrqOzybjI3RVbEk
1pOsyB10voeW29UWO2/kkIixwHLu3aVPDMeeKCB/5Tf5qhPJv7KOo0KOZxe9Xdam
QFlvIwDkViX+I31Sql8/zFI7jhd/pNXW6tvSA8LJHK2+yZ1jf7Kxx3vQGC1GQ+vq
MO7BE6hz1SEgQtbDrumeBChYa5Hie/F7AeCl5tQtSz5q7jjxir9RL89w0JovOoBW
xbTJn+r/GYmUwotzCb2A99f1nWnvfh25pkufL18JS0nYBUMKqCdC7WBSuqSTnf8q
O3mQmk36NhYUCoj791bitS0k63R2LfajGfumyMAR4HwQJBqsdZlIZ83+pTnPdbML
70ZsFIXrWCtpe43Q5e3WyFIMZOgjphEsqdaz+J9Ilg4E2stPVQFH4g/9gbBBKZNv
q7eSY8ZZ+Hc7GjitQSA8r6nZiFQtwIfpif1tWQDzYyoETo9A0hvT9KB4Xp/y76q3
jMNs8eKKiup4iQRsgtydoDZQegTwAhWy9zmqx00ObGovOkkby+oKPWKEHwccmxCX
iAdRUxpu43wKQyM9nhcw/0+qs3LMSxEM2nvutGpqcoXYvSbU45XrIq8yRm4jMA5E
weOIqDuwYkxip9uyCTHpvwhleTP4zFJ4at1UUhtAfkasSLtvR0Bd0Pch6eZm2D+7
mJEQhR2eUmaPYkQwTqkIVZMcwXx3zX+OB4BC3Mu+HJSrZwNlxaNQMDniJreH5OhH
ICZcx5QYggDXeQyIX36fmq44GqQRZrEyhjQHEhOdFfPrXbtetFHde9PFU1rjKUnm
5IJVbqMhz2ZizGnaD/GgCilCbqu1z++hVU8LDfJW/3xmaVY9tXOdLeaD0JoHNR3p
QCiGCIkgKssfjy0/P3REmpa5t8Yu3qY4xe8vyJ7Q92IpRsf7m3HWslSNnknNYDos
Enxe1FR/qF5n9v8SdxPNCm63ndzaa/+hbqfWUWEnXJyJSRs1WaX7ihkocOy6W5gE
HXsDXwJ87wGzedeHF1GRBX5xXndRYm3ZY3eNFYPDUGijDONMRpQ/zU+QhmrHg8At
10AQCLGIkGXg4sXsKWguYB0r6QkGKr8l7iVxBGqqAWltPO8NeFTPJ+48Kxz9HAU0
/+Lo7fSb4jGJ+SP98DE6HcFPD/uekJ0bfajI8zBabGlEAE0br6tb9QOPZWrSstPf
ND9abTPZ64JwOpSupPhvDyixnkp6sHpXoiyKCew3fid91wljPfQWw3dod9hjI1cz
iDLdSld8n0fK8UJDWGvkh+xFdQIrceIFkMH8jnmB3o8ZWSMSxBChqMWaTCgI8Qn9
CLUA77mHBHlKDYDP7cZyFx+ziUSO/ICvIJgw1Kd9icJDFXiCk0rp0PxOczTCsI5A
Y2z2bZqPX45nHs8zq/8op+oHzBL+kEhz9wZvlWTcOG9lv+OjN1rhnykfWZ6/D9j/
vlW0p/836kTv3cEd9x4ULPN/AMaIgzjRZYcw6jYCxZSdbGNWGgrlIU3XEA/dNeVb
t8/Mhgz7x9t8eY/7DU9szwbbOt+hSzl+4Qkb7YzwEZdLL4zyp6FnAIWgYHoihH+B
NgRC/IZc7lJdQTWK/m4iUXU3y2wpVN7eEELsDeidd6Ae0b+1P2fM1g4JBTJjGmhd
hKLn53xKUVKPijhfNvd0NTSChuvVgymuaaHJU+YPVgEeCw93KH01DfmG570CTWF8
Uk/68KAC+f8N8hPOUJAu7U1vJKmR0Ge8SC730+DiXRvxXMAhCp5ttuGVSsh7ts8o
/NnUN6P/hB+8NDreuLGFUo13p91TjMslDR+ZeDZOJVpIltuCBw+afseFL2ECbZkr
QhDod5pTGBT79t5hoFs56bIkcXy7UVgjvXdt8k4v5ALI6c+x/HtkX94B6cbV3qHe
3WMCfzTjcHGMYmOF8eYOrzz7o6koQ/MAg+zywirSGHDUoXW7srhJv0pIsJmv1Ow6
9Zhu0hWSSywq43xqsxyv2wUkO4wuEwphqqXXWdcJ6lQO2Z4x8AnYGhgRK0ZtcqfQ
oenQlBp004WAuAn0B4CW+EWB6udgjZgjzkg6vBwX9dJ91WxhlMqdXQabruftcL0a
i6ad3kXj7cArv6eC7gkVerDooxjzYzzCpbFc0Ijl9AuQyWjbxZufkYlUT5VTRsp+
AcLzWq30ORSr3atkh639eQcFiLerJmxq7dx2tWUV9iI+OiQAd9UZiDow7aBrEmsf
v0p8q8DJPRfCBrdQ3ikac1m6ql5kR73RFMjhP5ZjVOZpEAiCscsJ/UTS8FjoqxqW
mB61Ac3UdaHXjI7RysOv8kvVdZObANVh0e+ncsXb1emStEz+I0VGmAnH7yTfGyYZ
kfr2J6nHSexABklKf5Yeb2l0vOcICac3J9KvddFEAetqUueHF4aJe3iTG6HVMGMu
sz+pDDZ0fPc+HlWpkhUvnxqetUmOO4R6gZ1UXKRQtlkPyiFfro2hDVGarKR+n1ZR
bvZddz/r3LUIJTak+kbdp/fBzF8FyGB9Y/Lh1xL9KDDXsJe4vCeXdHV2WBvGPFqN
Eoliqyjo4AJFqBiUmx99kojr3IzjJP1EUONZo2LYNX0yE2x0+qAX3G+F/gL12A7b
tRoj03MAgIUFJsESvdmNPp+UfEtsY9DETAf4au+Mc/4bUHZuI+EGvDkx3ZLu23aQ
ex5MFFsjoHRMtjTJsvNYKsRW9msR0wnTt95xZ076pii3gFTBFHKawaWPNhkGRCfU
epA2DxR0fQgDUpP2/gBLPDRBAwLhKJu9kHZ1DmW3KD5TTiTnJZd3WfyeSBt0Oyqn
IwspFbcpUXgY032MqLVnk2mFdsnKQT0K2fxo1q1IryTTP5jV9slD4//0AJgyd2Ko
ajMmyPV+riV96JTltcK5MtnuZtnGA6WsneXpnIjvd0B6aSQx5gkMlh8Y0BcbTOcB
UZPzIYvzExdjzIN4I1RSm+lR/lb2lDq+EdROGTwqTaWDppmUdBxUxDXvFBMjMR1+
XcLUpG9DYTtmkozspP1WQ533UsJqAd5FvXb07fPDKHlK+tjNzh52lcSA6EgO2sLG
48Ecs56qM1RPAcvF1Gl+0/NTbG0LlN5e6APUXywcMyLV8pFVhCp9ZskF75rgVYZ7
1W6P9mwdDJDwa1FepRm2UEisnz3iVSfamBDNrfUWl1md+06+OdzleIb0+U+jBKht
Xqkj2RPZ9aPHfWNd3ov+pne2vIkIK5qskmklGpNqNy6q0BjoSBj8cUGawYa3yKyC
ilfsnh96sZlJYZey7nczTtHLed+lw4mF78bgOyOsFY+hrC5IwQtgjUHRnSWF8EE/
/po3wpEELn5kI1YMZD/QmUxQFPmE4LD5YA3OdaP9z9k7syyBIupuB4cEJn7fO5xr
ex6tRfUVVwe0qbTtzx9iG9b56loCS+Pgy8r/Dy09yJ9I9N1J/2tfKuJQlx+a9/VG
ExjXE5yND9KyyHBi85CosF3gJZVggnXEpZVWEQqCSmga3ri1oyyBWCLA5c7s/MU7
rxxg/mThceBf6+ioR6wFNKraYC3rxX7/yxpxXzA/nvBBg85x5bpXQVlOMjCA7Hjc
01YAYWrLhS3Thk/EBclB6aXCVWRd2sXtr3YTzBQPsR4vjQ4pTmpy3dLth6DIphfg
kEo6lHFM+FN+Ox7Qthqzdt/MvXwvhOXG12mcQ8YdpG+/A28IyefPW9eFMgKwapJk
HZJZ6Su+hTy6tbKKq2A6D6NUgb8qVhcjci2DX6Zv6bGPzzCJYhHSoIi4nR2plDys
fNF7Y5TJFiuG8irpp8uNt8ZGYQi7jM5I9XVPkdC6fgzauvUo/PiHMu1zbDagWX9M
JYMW49uEkOEXwLIPjKsDNht2ChTaaPb7ZALwfxr8VfMMe4L+8FqGyH6+dxNZZWDl
8V62A1t/yFkY9IRJvBZtqG3+u/mNRX1nC6LvkQP2MykwMRCfg/SnIIO9BT0x1Fki
dEY99e+DQOha2glDeV6bpzCwnUQrQEDrdNhvvX7uSAw+ml6v6zPOxAEg4Pwyhvi8
GX/2iJtrxJyFcQvIwu2UGSmPQftbqjtcPT/81AmE4P2UwTM8nb/ntOeJDqN3u98n
D4mFBI8msWXMeeAy4frjaqoZqEAxT0o47kqPnzuBVNq1yjvWX/4mH4Jv/iKBJ8UG
iWIyJaXzLXZGE4KPGHU+zLn15teuPm0jlq0wt9omcYx7b2rOWIogYHX2JyuwBZbH
k0NHk94akO3H7dSy7MeXBJvJDRbyZa6ia5usmO0RDWGhFhP6FW1+IoJw+pPmeonU
+Tnh2NqrE7xhFRSCqiMh5YU8bN8GgoeqDaMJbfw2K+muLxNDQpV0d8/1FYzB9n4U
gGui0/zPFsJNffJJasUVJ9s5hT4fhHb062bvejf4df3UUHc3YwqsF9h738sOvnqc
D/j0//4xlKaNUSIgjKdxEhmebOksxI2CNpYx4ebP4OPmPTxnCGYS0MeSYVQLjaKd
FLAZNu+8qIo0FB7h6kP0OdLsDtMDOmMafC1rphGf5B+dhaWjv5F/fGOQjGZAFmh6
Yu+bVGJZ2xZvJfQ1nWfJm934b9Jyj8MQ7up8LJJE/k+7LDlf+dcdl7+PVd9TzoEh
gthlcIG6SVDtSr1VoOi+l0pVb2C/Ga+aa4qv05yPv6bGuHf5djG9g4U3m5/YW++g
ueg7ypuSDsiCLqBLVGvEhPjuTcnDOsdvuHjRM246eo+rkbCLVEagITgMNOPtj8lQ
KzKJvZNo7x5JnjOibORfhFHkzOoz1Pi6toMxgyy61+pbZ1GY12M4EJ35lJx3njco
rYVK3nmr68nmJNCRcJvUkzbF0CugxYx+QimYhFj6SvYF+SnoSs1qpxP0p3PgFOoU
l3bC0XLu1OzIbVBuzOUtVcbfhEHYW6u9OXoeJI1D84Qw5Bs7oQK7aGoYdDaw17m7
kGU7/5W+upEjT0XwfpvDTjgkzlYxYhTU5EfEM7a8VymuJmRPvFCmuNvTWpVLEW4g
M9/QdyUeGhS8QQ2KmIur78R3mmZgi5XkriMRK9BrXUWyMVNJCZhYrtn+P6i6KuOO
IEpZuSK6VZrq3gNtJtX/NhdSkv+Dk+upH0GephNnuV9SOT+gOgscxcXyojnezNao
WMhOPsoWXMXAY1GrchGwjP0KuAp9KdjXD6dHt6QQaH2v6UG8DxREqgZqVbofxNKg
Ri/y7IKkzMYCFuZNhoEU/S0we2cy5OGIjBA204Ds7J5k7bV86xibrlOfN/jpgbC7
Mh8gvKt91P0esLj/WxMpIB/vyek1C/9SEAJ+2Kj+NjLUa0xlGynhoCCgH9/0U3sw
DafPlmiwWlajMuQcComZsYhmQhLWEc/9NaGGiqa5DvOOnUXu8AAgbz/NqFWAcwHQ
NNEYDgxvjLBZT3NvpZrQIrXDbiXwGWggjBmmADxoZ89KCbDpcYoCou3F44jTmY1s
+xo1OmhIs3wgANQDuvC1P3Ex4pwyGTNcxdSXlh44OBS4WyRbstli5MG5rzB2IwAD
fPD/vc+C9LQxWfH50Had7RpLhOQUHu9D74xNrW4157edl4w0PUp8VGbRi3CEdj2V
d4gkBFmxXZpj9hApAlFqu8+aNaTlBUVGqJGKncmXyA0883Ap7Uqzs4gIBuDB4EzP
ugwsQ5JuWYKjTJ2h0WUjDMbIiqub++NNY7efPdJEvCzGakhgxhBNs3UvpxkiVy1+
5uDWBtY7eGJbxa0IPMJaAtQB6wEqIxieH4qKQEkNT3pTps2GWrYUOr8n4wJ9XHYF
WfDqGHFqtWx4WR4zEZCcJokehrb5HUWTl3bRhx2k6KImKDehJB7kTuatvGr7vJW8
MhNdRcKDEYTcsdgTCmm+exezdNr3Q0eLL08Vl3lkQMoOsLgQasT2xLH+GBPYRLe0
ajNTpu4QMIVaqNX2+GwVHzCwcryDNIpSwaCLsliFWPPy/rfZ58yIS9WtLvJ6C9+7
KyDicp63I+tf6dIDs5/V6+YlzuQVHhzgDQuxnAdJH9H/HTvjZLIpPV8u6TMmuxiw
TvOtdcKTKdiQADKPUpyTAaHw3buVIUjj43MoVe26cw8oya7ECfr4pnfQ010QW8u3
V5v+0SJUhh88axtNdmUZZb9/PVPivlzV2eTiBl8OWuG/uhbA8Ewx/jWI6iIyC+UQ
9SWiSSQh43piVN3x4PeT9/skgKvQV4yVk6x95Tr4oYbgZo0CfuAdshVibjjYrnB1
SSF111uyezzkHMlwcHPfl1M1Nd4gLNsm9VyUA/MCd9vKjYp3zgBxL7DL0X4ErP68
JKndkv7Zg9qqiWMgbITc5vwhCXRgQ1KneM0tB1dnaA+RYjgAvulZFFKD61Slu3FI
8nLN/kqqHNwzply/PG2q5FRE0diO0WfQgtHxyt8BqsLW7MiRgDYTYHx9mugP4vFn
XMIixfdlsZ+bHCJGxOP7mep3h1GeGUdXGTiIbWJwaLul5REO0kpXXGPrn0Ztk3EG
4+np88rUZ1QNlYQ9IKYd5q6vifGwGyFR4R1poTM8dXi6gdwF7ViuFGgDJle3fdr1
1nObW/oyuyqkH5GGiYfSPDwtBttlZs1D7ObpwX/71fipj+Te2h1lrffjN6NvWsBY
MzebBRxJCKUbBvJRCSn8L+LgP28htQivpKxL1DT4d41TOJOy0u5S9+8Q8EifBsiS
qyYYby1XCW4UQskHGVRvQyD4tWu8WSPNK886hHoH57oyq92T4ADKfGHWPy5+e4Hh
PFo3pwQFemJxr7G+yeFAJM1ugG7wCP4laijB+WqrssIh0T/N3R9nA0bINyTdvbCG
8DWNyM04aHXG3bRuk0MVOzD+tBzq2nk8bm7HsVCF9vImMCecb2jRmgeWzIPLObcC
l/5U+5Sj1KB9JjqxVNNYEB5dRv33kcI/tENwqmTb6QXyFWpaOgdjepomjGrkadMY
TrARp3wV7ZM4geWN11JfovLyA4h8wvq3OC2WWqd0Ge4Dnz8u7PBjkkG75gwlTzVj
vSID/wcvcllm9yq5D8LPy7i+OvtHGKFmroc7zjAaG4WN0GXSLfdeQb9opFIgXs1G
WqumkHMayzIfKCP65oktdf416iDy1Hww6usQjw/P2De5kKXEm8Hyv3pEwlX6q3xp
2oMNJesXr0LrBuE/jlOay/Ql2j9BIkG9Z3asxaQOwwp6ZiB6H3a49LejeVR7+dkH
mVoP4HZh3n7vYKpjxbVgob6XOpqkZLQ1uypcgzAK69z5a4mH6uyd6OiySZBuHiQZ
KmGBdtsb0Sv6XZNRLecXN3glJr5/OmSTBcbA3V4pWxacVlZf/D7TicX6EzBZnOtI
KWl4ZAempYKTkxTRxO+fLclHgJ2QS/fFTEYwzD7i1s9CWadot/L3fnBhjmSP+B/c
zBtiQFOsfB8sgf9S9v/lBRgBtPXKtDrNFbnL0HsH5oO3Z7PduS9RjfX7Z1BNOYCN
wbSTPDSdaWeSD0++bZKTuQy21p5+ZloixHnFhH9VAHbQ7BbzhHmLBd1vnilpa7oG
M7STabFBbCTbkWOZDmWgDO60Bu6v5pWrob7dnLwtkn3sr50PL3BW7AkC8gsUc+dG
UDh3WBmUM4EpRVc8S39EbFSvi/da6UWI22WisgNtEpiKXWKCBSaSQvqluTRUVkOm
gtsR3BN1FRsHI3eR/Vew093KWYebF00GEXGpwzGjUT2aspib4WaPbeRee5sldhda
K2NXtHHtMJ5igU/Xv7WKvyPHuNiPt0fF6M28f+4ww9O4svZPrPAQYvfwhZC4GEeR
V8rJjht+k60dydOWl931lVq36rWhgnjkv/wSTL833P2zIKaYuY+AfJJx2USxktIz
2ubTkzc1pCC1Su8Y9DU5tsf4idoGwJzVkRIgBRY9mE8Ylsjw33RGy4y0qroorLuD
TpITbglME2LHem5hlG2+yCiD9JJ1IdXRwzy+v28Ff1wNTjL7MsebAimslY7Qqllt
OUBvK+vftfZ8ss4Ev0D/700XRSsP0cRC7cObxRdQkVXMrl7u1QZjIcHfgCWv0rMq
IzWtutyQMpE8xRgm6LNp2RcsZtaVbzLG/FruRq1VgEsSG3+J3XIZxGTXWYYYPGYf
jJN5R19dKGvJhRVgksxACQ5JDMlcY4LK68QtEb1tpRz7DEcjjAEa0I2TGh4bRZHr
Zfn92jvH/RJLEE13zw8ZcQMDVg02eRg0RSKELdAZzZ39VrGKhM6+LE50V77hSxbF
2VHO1l82HgA7WwMV/PCtmBZqR+ulDlp6eHi8pZJ7QkOXW4IQ7wjZhw8XIpeclHQ0
Y49tevTuDmw8Ka97BpdQMnwJjoDT7XGxscI9eXkZ6VeTsQezs0uEzLgzduXf+VdX
nbDDdoxFGuWkp7eogfMu7QxWvlYYLMMKKZHfIYErGuoERdKa1SIZLfANQSEBPl69
FkbCm+elXcuqOXIA41c1zLkoToCxI6L1F+Qc2i2H1xSruFKdar+FZHHNC+KGHCQ5
iE9mpwRXcfJDqeyBR0QVQlcztBJ84L/hI/J9fULoePGrzdb+Q/mFMejpC7cnOC93
Wq11v5oawiWypio1aKGxhMRQHs76BOc2Bunb2QxIuzALoBh1GI/vQ7xdUveeDKLo
qWzNl7uPsgdLI58vftYVHin4Vl8gNmd+xrt7IFjp4LEKZsG+F/8/T+iDHKHlNOte
RJmn1p8rHb32s3I4KTzHCAQAJYyV2SFDCR2eNpPW/vysiVtdHxQjdeqJ3+5pXYZT
nHpaVNLyw5kc7TpUJFV7eP4+BRgZC6EDOmpKiuktn/pL9qIhjWBhQHT1kFSAmKHh
+EYT3kdMdzDxKN1yBQVd8l3EGC8gh0aJ3yEWjXk+VOnM6LHdypIcJoJ1nCoxvM3k
Hd7jUZoMKp826+2BX2HEFzW0N4tOVXcXfF4LH1nkTrJQNS7/HI0035uAeLzJNgyn
sTAuEVhVceHEDp+FulAJhp6wAtC2ojtEazJgztPIkWUZDdCAKp6cYyY2NMT3jJB9
L8Sdk/mR/MddXwZSqY650f6A73rgHA4QECNfnq+r2RUIotj+Ei+TDrHZdvEu+4gr
SvwC9Vlfu56sg/13JGR1UGngm8OkDIb0X1Hg0hGoANfZBsBx2CIWwCqzUle2RuSz
Wp6iGM2P+M4rGq8meqNsLgrtFhtkx3QYpIew99eYQzQOaXQS/4gjQhftggmU2Vcz
BK4vdh2Gy5WVcRr8b1zj4xqmqr5Mg9u0Ahz6ESbApFoTjnvrKAUpBpFVDEGLIjI5
+qfWKd7IBDbFFC9H3GkuGitmc+o3YasLkc9Xkd/R/WZZc0wkTeGGyx6h/I4x7sdS
r0dqCj+RExR6SLQW+8x3oRz/KOB1SiSM05P1sA0hPO9Lmi1scjahRCMUM4uJjs32
hpIYdZjIAFxXDxNXw8TFcDbx4iVQ+EQwsnOw4x53mywD0PTqo9e+u6ELtQk9WCoY
/pDk2bSeMGEb02e+cjEpVBd3gJO4UXz85v6cpvwIOrF9KJkh2T7Vp/rsT0Mtyh27
7dukX04R4dRV0m+uP+oju5+mD3AQlDzrqmnkmQJVUSE9EiTrlUNiLY5mwZQ3LdT6
wD+IRMTwiPQz9AGYWONEldp6smkZNnNUKucsgkKl8qs4zrdwb5OW2rQ2fD2oUoxb
H1GDu8ogcsY3ToBF++r/t+QqFoRoxWi6aG+zsAGOAGa5pc3SSWG+ALkiGNRIVAHf
pmQrg0jDshMyIiC793YSC0/88WrKM2bKjzdmLrXhTBChBI5wMltFuQZ3ugVGOz9o
XSqQTgwNpEwqXoLWNuoFRt36N7XSJBg1zcjEDl++8tfgHWN5cx/Mh9r+9HRz+0th
RxOE/NXm3AfMa5BS6BAYK0BTqoviK1q9dpufQmWriJ62ZipwNORugD0yTVuCIfK0
DFZBxfwkDUwbvw26WCfVW7SFqts20oFSoHxutqL/psLYkkvHy/YfUQJ9slzS46VO
u2PX1qkAB5bnRWZTz2ArNxW6YufKttKuIGo9rC756LT4Z90ZtsXEtglp7AevYfhc
bDRJJz+7v+/hMhR2poLjpSIkMy7OnWKjtv8jvV6LedhDbd0oDYHfQxeg3jxxIiuu
2ejcI/QLbIDNcpOc6nAhegRvhdwi0sFPb1Ydo+XPrvUS+YTwd2HC4IEtOqLZdU+K
QpCgD7hAKqt7/rZgoY1FcoDiPDGEmTS57dBzYt6pClFUy0O6nXSouydXpkviW2jy
iRIpq/1fiX3cDOn1TTyhHcJxv41iPJO/Q3m3eveb7SocAFjXyGzYcAMSmTSlBFfU
yeWmuRfAUFCXJWoZi37fWlPWwrTUf/hgVXxKBDiFr2Q19Cd8KERCWaydWe9Rr/dZ
SFwBPL4sWMDIuCeJ+0Wm0ybaDuLmO+XGp/mJN7xrgMbmAvqNzwGp5Kjw7yNo3/JG
PnuaKaQya96Sj90K+UPcEjiirMlk0EvJQRW3zV1MXAYzImOBYxY/7w+br4aI5e1q
wBOiGhYSPQv8Vq7H+nJ3Uq2mgoxutSuyI53q0MOT/yX+/xdmmF4tYefDO5uP7b5f
PCQ/ohCKOOFzG7MkBcWmr+L4n8npok0bV2Rj9Y57sFLdIcHxu1qDoMJC5ce9Ybkq
bYMECfLf/uay1GLKLe7jFStZwKUOM56QgkK7L0USWpOVzfEE8+JnuHyV/O29sMy+
Tsrs5z1XeCXTOXvgUpkPO61W52Qg56GAnRLeyXVJ4PtfeflxrH2Dvg3/byA2nJ7w
K/9S0GTyksB5ahVsDGtlZzgJ4t2aI74ai6pSmpwEBirXCDXw4YJCxAJXOzDAJTvr
Ki7RxOHX1x4X6qCyvDh7+h7g0xtRfc1mJaldEUQkYLfjqrSS0Hc0/r+bKwrW9b6H
fW7vww46MSB7T5sLng+4q2z77KAzwhnX6LuwrFZJHP2ItekbUvewx2LBfob0cOLd
l8TH2T16N7ifZp5j6t/R5CEZtBOHmUti+YK3u9gvPOCIRd8XY9/Y5qIB+SnoRyOX
ndqUpc/4XSmo7fDTN9VrmRwvgszLaG6Ad73N/xEARabFmbqRGDvvgaKA5XxtTfyC
h+h1r57OYw0o2Ao03R4VlmtkfQ5T35wqyh+EHWEEfi33Ezx21MHyJ8G573tdECG3
F7H9qdPPbhscB/G0RI2Ckjyj7OWVaMkyWE6JskLPNpM/R3R83sv8CKGRRRUnYWYk
1v8KxlLLqO26BCWSWDoVZYOmjVkoaoKUSlyxRyujGRe1jXwruA67In5dbXe+PyCB
nNVT8hnjh1qdMnw/hVK1rW5Mvc3zFOb/ZpHwGcdsimaci5ww3uppstPc13QMgRGn
Mqvnmc4uX2Ul4JtMN4uU5bKA14ZVDjvUKuAyKkK5Y1+OPMhfJfV5fdWif15ONgGD
zqRlsMaBO2gH6zhCDcZk5DfdRusQB0UU1EwS9Is9wBmUiUoyEkQOnN23p10Br4gD
vQ2gFxmu4yroH1tbUnjtCkqgN7isBZ3QYPoYaAxs22+S04sBmL0lEguw4hvTGr1n
EEpD/461c9us94n5b1kxp2H8g0OaR/8mv8X3NJG1f/EbL3m2asu/lmZv5YKGNH7d
7plGYnCfgMUKg+ihFn/Fx1Clf/+E93I4i0G1JSqBUUeD3mS7s7CwcFK8DHW6/Gjw
/Mm6hmy5KoTF0458NkQfNcliE4FFHyAEMVW9HtJUWkeJGsKZwnaxOIoc5mjmkz/p
jKrAk+xEdtQh5T+nsMBz0zxzYV2Lp18MVx2GL0bTwmRfGPFl9LJNqkDAsxjpa7WC
ff4xrWGUd1ZeUYaKY/VfJ5KMDp0L49tNA4D97aswl4la9Uy5XTbekyQgzevLN85q
+y0AR2f4MXjhhHUWk4kTHxX1w9TZo7Rpu54numnkXvla0z2EzRBwD5n2YNVvrqUV
6ArF36TIct1bF3lsJ1qVk9O9xmwz96pKYtGB/RSvXkhH5TBIoY5W7KpFSjq2qmwU
3QGyf1Xegmrcdmdn61cfqHjeZVq/lJE+KK2dB7Jv3qs4cWrnCzI+ti/H1G4l7NTW
Ml/H3DZNzWL1D8XsoX1Y8U1X0DmCZS8lilKCsBcDWJ0kmDDdhkumZ7cs+9PjLmFi
kL6YgUOYs4dq+gZBv3VlCtMYfnBiR3z8e2FvkOTz88/AcVJfsqpZWPOEV2RKY0By
o6sLo8DnA7aaamG895RfMTD+Bee1+DPOnI/dOyA1Ibeg7JKmQGb0RPT+WFwEg9cQ
xUvUlIPRBylPaucSM/gaeS3MkV6VxjOMX0xJc8agdT6F2K9geTDMs+Y5125tQ1in
GQxQI6S/3vjvP3jB/dW4/lF/p70GGk9/ea07q6r44dOJVl2DnWJKnnXMJS8wOZ9L
ZiY8eUdvmVEJA7KfNWhBwSUxitG9C0c0wHo8Mzjq7mYHDQXk9JmZxExOb8LJ571q
xyQqxmSbTblFi+Vzmzcok4J1fx9KZ7IBXIziFGOX5zYzlZQUVtDpOcN9e99ShMeN
pXqf7fIBlbXnEHQL1QHQdfblzN+aqCQun1RwDpYcoo/Lo13v+S+cwFWEyY95K+NX
Uqj2ZROQF78VZ7L+OjivyFhOI66ekOm4aEG9iv6BBfJ/6TAswJ9bgRfHlWHuMYXF
yNE9FJQhFBdB5YdyLC8ep0VIQKABVS1hMFNOYTouCgW2fSGvfIKXKm5XLoA/7lXC
0faZBsIk6SR4x5s9nwvZIOna/oQUTxtU52xAmMfPkrjG05jrmh1nia8elVu4gLhv
R7yGMCeoYi66KPcUpG3ATv5bNB/gpcFhDsxvorCIsqHSIArKe44ot1UysqqXd7nz
wl4Nx5P+B2V9j+Pm1S7bKcrNvxHWAOoGzKEBZmFdjTwwJoV+FZFrfXul0iJGCZkB
eONPmGpj31TSZeTgkTsxdgv8QmQ020ZjaKEB6yMwDsYOYpzD6sCI4PV54eI4VmsU
zCxm/ZIuWYNg7NScrRKJO9smo/vS3nx/B+VjBUaiY2GnDzQ7QnOx0D5iVmKsouLv
VBiVnC9EwUoDgwQPBrj6YCYhBH57+JzG2R1ypCiFnh1QB6R438TaMR588p5ojY6f
vZarhXNgpH0+AgNY809fE/fEwGbiEtHqSVFgm9e/+2629fQTRWs5oNstEegzIgIg
1bAou/BveuGu63iafzmhhMRpiYpEAgbUJRf0diZohmJdZYNeoVgqYRP0HHx26W+0
MvnUuuui7k3WuWTE2K+8EIrYVg4GpFKSK+h48iUXJo0fyyl8ztOI9LgypJCT7bTv
H9CZCmPCNossENBCge3Fa5ZV9TvCNOGOqCJDTLj7fcbV4lvwnI5wYG8/kVB5FroC
MwrOo7USlA59h/SjRSOy6GYCImnQ6R7a+lyJNuo9s22pUPeqSUSLc0hGbGbrHugx
CGyXNcWSZW6qgbhPipm4y5vBaTCxP1MXhTkJUJvbCC+ilU2z53YgBDebz9we372G
q7JcR8ufbf8pml1Tj9t0KMU0E6XTdCU3nOtVYVqo6ZNcUQvGHbOWpRss8jd4FEAh
cNkS6LBzB/263wivuVBnFB+sClXBhzj0FSR2SEDNlQ1Hs3QSlfJOwkKoJlvP+Ifz
duI8jNLr0D5gPF/TiSNOmAT7uJUp3Ns0mYlVWYQFedT98x5dv1MEe7morFB1PXfA
1R49ivQSd3njnWTTh9X8I7jUUkJLSwqgfSJFMgwD5M0i6LkMggFdNECU7B75dzIf
GR772GxGy/LIpB7vu5yvqrAy8+3QYayAZooKFrXV8l/Syld0ggMExLFfnxBytQhP
j+Sj+twpfpNvLMPbiKLG/eHJR/0cljCv0VDzGl91c8c/tCwvebwKCDf63hEBA4yq
l1BvSlc8eXDbA/KBj0pl9IIV6IfI9NzAO+NEjwN9HaXVeX+NJZYXls5UM+dMW80H
bx8rSnop/Mbkw4/dHu6AUSsfYLA5CwQakvTPpNf4hRWIw2LySxIgLEiQo25yF/o0
iIgWhpypLujuRSv9qUPGGdjPajBG4rcXW1k98GD1Zm0Ws7HSKZqlSSLgsDFe7rRI
ZOSn59QYADmd2Qn4YprR05r8TGp+mpm266hTND2BpZCDJ3KJJEN+ztLDRHILooh5
BdkNL2vUddK+sMhIRvV6OY7Sqbx2L1VHOMVSUiLTvv1zOmYwcDWp7wSoOjdLFbWt
XBbt/ByjzOIlH8IiWqCgv8ujRsse8Xjhm435Y/tibz7Ss2evS5vpGEmb1qSzv1tt
nSJczMVt5eieXkqNd5o4pWff9qOaOdQyprJ7ZWoJK6kpToyZv6PWSm7sLUJjk8Ek
rYpbkILM2uGd3DLOc8gruuayNb/q0V/gu1be/eyXWS1MT//dz2cNRqB7jHRrUn2a
/XGNbWCilw+yq6yUFvuSr1kx7ytTOLoUa+MzOqHrjIoXSnjw4mVW8Mm1ebCpBPCe
9URhjeFUin4Qe8iv9Ot/ifJMvG67IEZ/lF0M1n76kQNiDoEXOeujFbyyHsMBu93Z
gEAqpRMr34hzNUKfa0wigBSAs6s6dqGwapjIdwvq3FZgBAQTU+15oUxgxO1wJvHv
8ch7KRILsccZii6TZ1NqQ+jUY7Zvau9iJnunDpyDRLNHjkbI87YMpByhNOH/tti/
y+w/veuf2sYnNKwyHpCDlzPfkSYeUK/1w0/hvjZZvpyiADQxwTx0AHoK4e7jJKAE
KT5XS4MUbti1Pk2KYJdrceKG/sDvLZd7ZMuL/utSwFRMXgNr9dAZBh7tM++jd8Ej
j0SI7U8tHfA6K/sPYA/N89IT0keMvw9x7z36ssYElHYo76P9BVg8dXQ76Jq9UunE
hluJI9XKcdD61f7Fu6Cr3tO7LTDQzMZyw5407zt8x3CrFmd/lcGNMieIUibR8eD3
6O9dj9FXITgzCl6oShh82RE4cj9IclGAsM/tqMmJolqsgQOhopA7yUshCVvSGUNv
6UDvwcWbywqytDpAuoLm3N7oQjeGCXWTwBJ47weK+Uy9UbLfBjOJ4fTD9QlhsD3C
lQ6ZZBpYQWuDzD+KLfRo47hPJD3zB5rj/KQlSGZFT4n/C5kvhSm9vaOTLC1hqzXc
IglldpHI2VASOi+aH0Xo+GVZ/2tGq7K5CH4Uu1TlmFXEsFNJkZvWfeLrcVwKqIQ1
/kVCif0rtsijv4LKUzQrTMq4Gn6xHDskzYRqbKJtPT28c9Iqlon5vsbz16gRGip0
NAnsyJns7J4HjHqx/GKqWbnAUdT0Iz8sJdvmPVOrnabFHYu6onCAXJZqtutAFKFU
Aidc2lyWdYKIMBUCDVhH/WgWHcihadLx4EVG6h++qhIvPFL36lP/TmT2IZ+DxhHa
udCo3dObDJ5Gkh0p2oOzKJTJVUm8Y28ZQ5LfCCi1RAy3TrAmdQaihz8zbeE2pnYk
RDe7noQglj2eZrSNSjckRu4szeGAH4EBW3Y2h6XQD3kf+Kxbl9lhp7EN2CWLLaKD
mkOb8z/nOv7RJYc+/b+MxNtV0nvMkLJWkFcoBzRD1BXovOKrwZMuAQ4m66h3c7vD
3V3rJC8FJ4G4WxBKiU/XLLVMZAx4uFhOpn7pgLgxuS1wd6H6vh61tu+qBDzagAin
iRzq9OIEffv0vqGZeiiyCYyKYi8cLVp37vOCUWnx4ikMy2wHaFKF0/SbN66V/i+R
QP2bI0GPUBVJRdB0Umevo8pe7ue0T5t7hl14EBrOEJdNpkdwp58/oVak+fbbmeFp
V/re7mOyODPJakNmFdnogwDT2Ep898PwlQ4e07Rznue+K5qEk59RXuhIa/j81CfI
Srsd4O5urVySu5523O8KAXAapSPr89GO+4v7CYXM0onIvHJCloWFeLvoBZMzq5A+
/x+QSL4YBGU6aaz29lcnqWtSKVSmeoqn3S29dy8cWaBrko+PPCvwMv8bBH+8UuE5
c52BNe5wbWpE21khdKTUd5DqMmJe8NtVFgR3Kf73YCai7UlAFDR98CxvKwrlpIWb
32TUzZy41aMT39wd9GoKsbDoG61/V0ZhaCnAr+veFMmYcqNbFaee5AHRwT7L1pcr
G+U2iY1Z+JnPpJzSUkwseSIlz++zjwbRiSvKgFGrije0D3e+OASA7QyHQDKifXos
Rb0lOz8W1ml0pOQpIWJRWFV6dEpgUZ+4fjWEvwba18ut/7TuP9nZrhybhgtBSZtt
2YYDz+lf2NLRWeb5qxzERf3U1INISFt8Fkz2fQBRSKCdLSbL5I4plklMY3fBZlph
qcCTDlg2AiRnYWmqggMY71GPaErT9dC9dfL5d6RGe1to8Epe0wbLlwUDEMM2dniF
ril6kbo+Ecn/i0CXZWapc0XzoMMmjEYQa6keHVN+KLIOsmlV884b/QdgHeBwA1MB
WLiV9O0NnvEX8RhfhckQxDNx4rO8xmxvNeQGdPqMNzJKW6Gy58oXDlOLDn6qO2yV
1vYln7+77ehk4GviOn+SmZF/bhfTHtm77tyb1n3AlPwi0E9FWYOreMRvbwHvgl+N
luUI6VFnJ9znpzn4Dwd7bMUZ7dG+3Hgmyx7HkI2gznDlCreKYA3wr8YqeHCtvoEt
ya3PLR+24ZxWvBTI+nTu1ku4+cl3tXQu9d9GQQr4/Nm74RBH4Ws0atXmtzxJaJwz
Nix/6dqw0i8qxoazI/YFpfvS/ZtKJQXCiOcQcyHru/knKHQ51pB/Qwg6YrC3AMP5
f5guWZjAiNix3Ek2dvEVq9NNLWZ48iSXt/O9obO4NGLV4xNhPLcnelqXC6rjZUMu
n8DY6cpZf7gqtw+LGlwp+jaXj81K5JpIhQvRdeClqxivuhZq/TAZiEAIwjSRd2Ur
q32dxMFHKj5x1hgaX0fYQBpycY994CQwST5tRv04ftovYPCkqrLUm8R3Myj60/fH
6ilD5GEChf/tAQaoNoHKWaweb8xvgbAVSfiu9XnN4DSza8Gt00yObziWlP14vJJx
tZ/vFGWwiE4GnczKpqbrKH2usOK98L5cO3y7YaOrTuzbih6nfXBhorvYZSgrsZPz
m0CIjfLd+eVc6MZR08l66vLEUH7SLvoqGjSeNPwAbJcSIdt59GbG+iEw11uxRVN2
ZNLKF578EtInBPl61EeLkrEix8R4WCzL/svEH3cl2QB+1lgIa1SfCIygyA2BV3Mx
hvEkCSVs6xMBr5/e4bkuxQH5QnD6ugUiXtkQGFCThtX3FsiDUxnJqBTOS8Gnt6H+
sE9ie9KcBM8KwRCN/xZa7RnS263zpX0yMYWcXSl6fxm5u2Y/o0wTMnV13u6emC/h
lnCPKkqiEeMR1/To+hEWVv38GF8EjdZIFaIMNM5YdxRK7Hu6RkeSwM7uYUdkNpBH
kMmDzgIqFRKip5aEQAoDGVEKyr4Wvrnirqg7eu5gPfBoOF70/9f6RXmGN8wjteEt
Ip1a9ruxHIZn1fow0zxosgLXWmof7KfNNNUhJs1SD6Lq43s1so0a5hh1SdF78H1y
8qfn7Z2ZQ1cSYwc551HVPm/6T0vr+3fsm/25S107hFIoOt+7vRfyvZiqDArfvUEH
/k5R6zpq52Jt5ItAasnY8/bnDFfGlbxLAsZ4yzWk8IoiQdeJ9x2tM0Pl60zSljha
i47x51mzI9LmqCh+Ko7xA9soP5wdM70cnbLN9BSs0T++H0jMLWglfvDtNA7DMNxd
HwfCOrC8jc5/aubxkzy0VLCH+NRe5VeWkleGt37LvrXSf0pSUmlv4q/9U/Qs3dI4
vq0GKfoYE4ENrkJ+ygiUqcZpXyB5qlJqnVCu7WXsMF7Xc3MZNJyUInJUH1VFRHmq
xROs/s+cqEEnYa7cOcKhjk8Nh19mnykfAUAsGErDixUrLJtHRZ+gmuqPgLaRlap1
K8vvKvUzH2cB/kmZ3KzwbNtbwTG/0QR4WTIMINhODVs3VZGKC95Kdlb95j4ImFD7
wHLNLDj/BrUDVdzEjDZ7NEhkSvzFM8k43y2GksVKHDqfNDxiDXI6Xi3Zr64SwuWU
a2YPZu99onIziF0vfD+2XE3NzdyinRrxlRIGeWryvLTXmpWPoTUX95bpbcN7uEY9
XsN98Y4zwNjWdYa1GKmQzCl19pW69ZQbQQxjRxcr/iBZjvzB1KqF2FIBb7wErLfY
2Jh34H4USPqkp/n/mX/ptSDAKdPkHXg8kBSfqMs8+dvrXEqidA/b6pcoxnLONxV2
7De1X01zY6szkYA+d0YMPxN1tJjaselbLRpJlRbjT8YYVUCtpaiu2y1cCU1UbabO
4x0LnVvMhdpf6id35/z7ozlE30Tdaqbu4m+vSIbNPTXadhlGOqwoICoyA5hnKsWv
YlkqFQRPd5uXqexYQKJiZp68760eN+ttKKxfNlQdfBbdL867tD2HGRtNQC8YVI9d
RL5mieRUJGS+Lh69FXNHzcUsF/kSPa+cdO6HQqOifPru3fmcsKbJzaoLDllojLcd
4CBmQgnISr58CZegcrxWwtCEhE8dvxFCHMZieNiI6FDpdFytLysmfMigcvjR2bMB
oApPdO5QKQzyiLj0yFhhCys35ORV8GHBP9bE25YAjbm/yM07kfTCYGadXc+pZ4BT
FmX3VzM1RUbHMDpkc7sgoyTWc+qDDhLStDmPh/UnCS3rdh5ApiBhEkVuxrioDg1C
ZTIZd0EGwDZVXQksLrObQCIv0GKH9j8a+W23W3geIfOSolHoXJAOmxOn8iMoXvWe
bMk0II1yc8GxTwuzsg7Qk48a328JRPiOyDBgPuU9Ecpy0pXvJOU5ohpasi+PtEPL
3wOjsVXlIFXLO6LByf5CWYkAN08n5W5qhNYfrYLBr/UnIUaJ7/ychnI2LoGZ+Q8H
SgZr/b9Fp84+2iBeanG6HfCVQ9W2UaMtg58CLxN3RzgsoWjZvhoINDhcJzjyaxNM
mR0efU5S1eQvr923eao3kPCf8P0SHlhLOxAIjVC6EbQtPKQLhHPSbDHe2mGZLfmI
UWJIy5mGz0+Fl70y9zmwnut20iJBh2xMFWy4zUge/cdi9SilZcrBWeyJ5p24+QAl
66PUdUOo5Wy5RaRV61STSIB2CIt2OYehT0GdLlAIXmyG4OjNIjjYMDubdp2P7fuy
FlSU7KDfhYhzlDXbk23Md6Iyv/WBJyCUvbm1KXmmTKnwIn5SY3vDxnVOToghb2/9
hB19yIOZ1krcSYsWYMo5koJGM8r37BKUjpQWFmqIJsp8htDubFF+2Mq1eOdTXQg3
6jmWPbtFvFDvIYG4KlAKm4e8IKxe/SgauwCijmFPR4vWu0OSgJdaQ4yqjKFYk9cA
5vU4RU+8Tv+UYhpisfsrk0Nvk3zKkBVyYMQrttGq7vtg8owZvwG2UVEgwnTYG4zm
7JJLLWoqfp1MEz9NGA+S4Zf0oYf4xWS3/lc1bnOkC360fbCCfgvHRg5cJQzTgUhO
mmAF6dPd44gpoCi8mugn8CNqEZVW1/4WMT96wb6KJLZuk6qQyu/QtL00O2HgIsU3
HUNYjtV/+VvDrDgmwT6Nx+OUBW9GAnMZ6MwX3qt31Rm2uu3zuHp03JlbYv1QqgDo
V291r1MK0hIaQrqdTB5xA+kAfYTHUaskjy/6kK3dzPkwp4S0eSBawHfYfNe8JI5h
oMcIkh5hW//+l400yoh2dCZEpD2lkZZZwB576Z1uj2AbosgD+b6mwPP9Dpm4PwtU
0uBnfZk1R0r15ltF3pU5Ofe/fbMeoIXxKM96yBu+72sqs5BMvh0koHUgzYEhkS2c
ekz3lA19fFRDSEjCpZiS3MBGFRKSOpcmrOrvQ9HNDMSdUYNhO0lMYK2aAZxN4lbU
34vttXaTZkghg0R7NdVHip1b+8SoS8I33l+qDK1h35mRf0qai1w24tCbVVIlHX1D
lP4mR3H0B/bNmMNz1SyLdo6IVcCSKur1/2u2z2g3bqZMbVupNLSMqpGMXPGlbzlU
R+5W5Nc946smB0bulqIgTeuvWhEOGX1oZ6hIh/K34GgVwf3x4r8vzRY6j2Skrqn5
6U6KxnheYL3Rum62lWYNq6BQVaeftwJ5RKPuRqZvNE7EjharWz2B54pReojkvfHy
ByWA1YLr7fLVwBdcbpz4kt499tUQJD1a2dyuZNyDBGsNrM+/CBiY6r+DF58W1Dhy
Rl1AHTC8mhEKUAXExJicu9o4zvoW8fA6euuw1MTbkDroe3jfX1DTgSbnIvfY7jBR
ikNh6XjFJQhxdevMuaDQdhj4wA6DerHP4S0NDtfxM8SAvWvR2ZpLl2xHV3Q6yrj6
984jzI7p40b10xWiVEeiZ01YEEgbIgCM3SwkpxCNy85LaJdC8MplqUWRPGhZtU0P
V/LFJu1U9YA7LB1jbjqPxmf1KnXEdTHUHiz4EV3GCgD2zlcHyEXnsQSLdG4Ragkr
kGyMlEeEPkHuQrheETQi4HmHr+yWR9+nfEd7lxaWAqfFylQxpmnL0MomtU9tmWWX
E8AnrL43ziIROE7Ew7dDNVgKhAW4mNIeNmBaD9QAxOy3nT3e7lVyGQB+8Od7RGWl
I3wdxYfVB+NYumxeUQB5KzEg8L3ju5kmLqL0R+9p0Cml8ZBhE+/613mFZsGMTPHE
Ks8jmO22iuxUcsUVZ3agqX0CVLHkmjN1BvRJICo60u4FvSPak8pKG1xQkVF72240
28iLN3DkiTTvVaS3Mxg3IB0nnQEgD42Oywqmi4IdOnvBkIsjYWSuxWR3EnwmHF9q
gBzGZ+589g0r1FVC/LxOhnXlFrpLxnpUghasxk+e/kpWebcfDHTFtZUnUhNi78ti
eXKeMcHRXdt1PWUK6GySTg/r+PsbBBN4auMejOvj094F3S6hQZwsvXouznoaf11j
SsysGwByXXKNVy4j4ejbJ6ATnUBiWRew4PitfIZH/1Wx2rk/bF4V7R6HEGyLMBta
8orYMWTXcuupXqJ/+ozOrNBTPCpe/UyRDBnABgkWDIut0bdpkf9fT3LmrrRBjYKF
ScRKmGQSOHM0hWYeEnDPnPO04Ni/HWviH434gjFREwz3gx5ayKSJJ2o5xVSyJ1BR
l7m4WYiYKAkyPXVw+b6kMmTodkDuDXxlgw2+nJqq7zvHU5xEbKMD7NiBir5JTYV5
EJ3xHXwdy34MMXRLMgRGftR+imDKHdh3mc+5iFE2405HLFcGTzF5P7fi9JfIrLHv
197UGgiOwwXjtChFdDWHfLwe+7rAglEIz21lZRyF0A7jQ4TR6OvX8/eH4Jai3LzT
tmGbPNfeWlBkI00eW9m5u0wCcSsGxCefN2Pf/FY53WdLA9PVRnSma1SX2o1ggawM
LOwyVIyFng9xruYg8Pn1X7wqMxNDi0PgY523L6ag4RQ6sY2ZI+bojOrjm1p7TBHh
vXk1psFd5DMT2zLzecgMpdHDpYB5ztmWkiKjGOn2AjAzzi5ZlMAQa0n7wBvYzu0H
lU2g5QcOHP0Fz3MjPPtRDcE+WajdvYV/0fqJIy2aNbj+MRuyXj228g6ATIGXSeRz
yzAmGkV+w4M6jWfaDpIkSTWNcxF1GRKNzcEN3FdyvWAf5Iu4/u2gCmzNkikXKqGA
JdYtZnWGk2rKzG+P+1M0iDBG9ZeoCqGC+bMzo0hglJ6W3xW4Q0Q8zYX+IZ1HFOgP
LacQglwvYhViTjR57FjkdvWk0fcvFOqwdRjBLZH772SvSt7tV6m+tsKhgwuOsbT4
k/q6O+OPlYQsSB8ZMKXsMBOPOVHCgDkXpKQEgGWwUkis69W1opc4hQYO5GWMWyy8
sbDUwhZafml16BMGV9loSEIQeJcj+2GFPuT6vr3XRAiINj6H5NZ5h5cPp/1w11vV
Lr0j2fB0zt9XSheiuGnXaJ6hU39MNnAmkiXUo5Cp7jjU3J2TNzLjwImV5gaVjISo
LjiXMFM76iateEm+LbK4uPX4N0XjA+puCtoiB0A6E8XUdRSWD0S37+6kqJrR78t7
vNpnT5umpET1Oh8MW3EjN5Snzwlw50rvtKUzuNxCU0Jn/oSbKCUlCNuRaQX7RZ5m
3FkwWllaaT2+sFy/PzZeqp8oankZVKvBHow6qkl9xOp0EXiVBCKDHZtZdvlr1oxD
NPSZykvthCfohF4mbeeqG2JKqNz8hrgPdbu1cGaQBOtx/hrMvdGxe4/rx4CZO0yE
IKhlybMm4KsO6fCMcBP2yyFfQftvRFH0c2Bj3ZxXogmhBkUn2P1dK7NNqpt9xKeu
TXwJbKctf+exG+V6GwPTkqunIsVAjMND5NYFzB/69t2iixCvdfM/r/AEXzwo25Vp
zhr9/L7eZJpdpr+DxhhvUJd1mRNhUFiwN4GF3jEarBPk7x3GLFaFIzAY4Zchqmb7
32EBiEajkgl7Gt25rGxb4HZSF8lw4buI0i/wn6jwWa7pTI2topBx/ZjgiN8+Wik4
NOltEytFfHg5XxaqI+NygJa5hiYFHVTDxE6z8sLzlf1PSOxpLMnhb2RH/O4Lobfk
X4WVmixCQKZ0NqOuvuxhAAgybtz8rK5auiH7rrJJUG8B2Leq7TIBsmxFQCp3cgJg
01otsu5Z5T/1usOmEK8adJAxNv+DMdZf0JcJcJvz0mHt4a2G/muCaAduNUiCQROU
h8xahL+QaKC8s8KP56UVpnekiSI/MJ+Tf4Z6scmGjwKdGsACWloyAA1JOHf+pxcA
juAMB670N5mldNM3P3AfszRwKN8fQ9VA98MT38NL+EwQcrvwS72MnmUBa3/lzhaJ
3EeczO4NLHba1sZxoMbe46/lFSdhN0NmrkdWSgqXd1ype5G/P1yaAn9cgmtbdN2R
hdqlwWZOhI7KRx0fVlLAmF3pY1oXHddTVtn93jHO/VKfTUxG1lysZdJafJPLsQch
bifJiwETqO+ms6YHIMLLj5znpfqdX2AbSI471qRE5KcK50QU3+0W4BxaR5ZvIm3Z
gCsJqbxZcCI+BwyRKxgr6T1GvtK1ryuWIfGwDFniEEixA7+pVBWnyOsIWSCEMAFX
JRTxx6Y07fXXISq/vGOxaxW7TiC2jfbb8u2j51LJh/bphZ6kXWQa0Dy6/cXRE3PH
kGRuVerWObsPjoETRYaJobpbYdnOaaiu7pqc/ys7yVuDEz9kNpRGEF6ilYU3GzFG
69XTPcIro7546nQm0R7WShBUohEyBCI+iTvJS0c+YCPnv+6tgFdCDgHLp0lvVyKy
qHGa2i3l/qn3BDHESFm5Gc2z9Z6glUjJ47CzjnKrvYV9RWa2lpK70/QPp3cyllXS
D3TerdgEC9pXpBfTw+wiYwZWhVXdaihOSeUL8UYx0egwrkKoh+Q0qm8/Yk2qWSq5
oCZi+Y4vjJFGAu4kRTHaOH7QC+ebdGV7wuaxi5/pNLpudYQaL3/sZ5oTmKR1sf6r
XDAczJph8g7v3nOnKUDV6d6oziVDZvO2u/euEFImFB+SH4NYuRYe8D0PRiEg2ffA
UivgxfSghtXv6RpWk2GRYIdU7hJsstyYv5TxFb9bO3hoCSbhThpQ+Tvpifrbwyj9
wszv07KCVu9r+8fr7aMp6n+j86mVIVGj5KdZTEk2NpL/Rw6OTewWi3Es4ryMi+WN
+VdV+hN4sVCFBBjLUXJl7MCceb6b/i5siGFsBN3cglLeE8ugQ+RJQ2lxKX6aUX7n
iztr6VaBm2vSmbPb+U29R6qBH8ceDf/gO+B4iF+fqyab80JqBaSVW1wHk4FKqAqT
oP9OuTTNY3V46ot1sFnfuUZLskm7BelkdHgFMWTTLnIhSS01Wqb7NhbEqfIEb1Qh
Ziagc7vRQpo3AfS0N9Fvc29T6NDqkps6eZrpRHlDMp6pY1DQUkzi2iJ/iYv4Ty+5
zbUZl5w2eervYe+hksWXvKgsSCTcayiSpY8RdNj6ogILNlrqdIPGbipMOTt0TIpI
qVZxCuPg3lvv7lNrVSTmDpGHrntUZTomuDogrFdgirTtfLFxfkqc/mAw36weexNt
DARLrpka+DexnbD7umZ4bVtm9GNeSFIn66Q23HOSEkV6kzn0HdyAboewBxyGzjB0
//6+TaCtOsSniQgRVbtJb4bpB9oyqd9cYgvD0JZ05TcSe3vXdDM+dD49hDk5izhq
NlBV9pG3aMuDGyz4rWXtOwf/LZyWJEYxLocTG8PZOj0Rx9Dqy9y68DDLVwt7RqsC
U3UxX78kHVU6aXzk6MMVlyaZcvZ/82jeAipf1iSn5htyo2dAGJ9ODNxGsIhRDTFB
FmqKMTu46L1DfArxr1KMwT6B7DjB4/YpQCIZyoK0IL0ZDyw+dwZ7mT2XnJgxCVpC
QDjI2TnzFbQ3IFPaAfbA23ISlqXBeF7soSC6HzvBbrxTy1BjZDZfTqLYX5AyREar
OLsAYa5h3yT/LRdiPrUfCNvao4PUquufmcql+EREh+K926scOZrMQExfrvgZDhSP
aYGsxWU/vpJq6UbbA3xQvmAucEjZVA50pQKgPRpvmn4luUiPC/ckOtH1O3kXBl4G
GvVj0G3Sq1SKKKdBGipn9F6uwpkNgCEeRJmN+ub2K/Wy5IcB8hIRmJwJ6UYG2qft
AukzJrQTws2O4PLo7W0qGZhMJXdNRQXM53OG0a/hOtNV1wPELmWffXA+vsWNLNF7
XgjK4dQr3/eBvh5FHUClNaYwjjJo2qRnQxKD4oRXM7tXmN+3TLntfeI8iG8X0pJm
BcLd1ndQO/mb6k6s71cHG7eFq+uEvCiyWhIjylUTdMggmBekf99MsZPMOEqJfiT3
O8KfS/qWZUWV+p36zJTHkox+LRJMT2M/2iHIqcGuYkeLyTTBdvYckjbKx8RnxTwa
om/aWDBQVcW9z2KrtjcuiPaMf6IYDAbriGErf/D1lSQ8GVhGR1kwf76UouNEHXs1
jJXoQwM8UNkqVDuJqS73qes12rmOjdYQllznbL2bc4FOSCaYcBqauXgKTQB9KNVl
NAoARE9OhyVEX6EQ4I4swu+z6RjBHyxcpY8r1AG92eEJ4YmxX6/XgRvs0mu5XdwI
8DMQSkn/MKIIaRHHMqt3jPlUuCHtYg5WDsHM1jcv5yS07E38b7LCubZrLffuZ91d
6g5p1KTdIweHAv2nPTh1Iz+JG3SCxQr4axvFqc7Dtf0roJVG9hA9eFOOaySzxAC+
LBUULmgJ2wnIy3ivgNKXf/QvkHjGco3/bFfUOEWfw/eJ5U2WnfWs+vzLhrlODCjJ
Aj99hZLUXuDk7LfTmstuEyC77R0qWTTlzgih4RZ52OWYJzlPUzWBTPfVeJm4mQvN
iwyfSBErbdluclUxnnttiz0ro7V0jEpGrApnA1ZwoeJd///OOaOpzx0fTlfGGP/A
9tP1CQJPOAHNYhAskkWh+uiXc1tIdrHbkjW41PyCmI3IuEgt7XKCOR0VWTsJRUTQ
gUdhBL6UmSoAw3ZHscWo3JzGcOlsXtFhw6KWSM4EtkQU8cLXLvFT5h3nnldcagRm
qjif2b+6odo7GEubPuAOTUTyLxRj8StZPvj805IXl8xm5AbIgqP3KYEBCnPwcZyp
YQs2mPQ11AQY9hMHkCmPjEKMbWywWwsqGBK7TQLR0KoOTYPaL+7yNnUcOEdZ99fK
f6Wjm6Qg+/o4j2n2A+gJyGgK1qTzw93JY4W1WHxImHWR/yn4nZtYDrmro5b0UQoB
pYqKKW54VDFYZQDzji7+KKXZNy0kUqaTCwD74t9u9lg6RIBThlLc5fPcrzsH/D7s
JSlyLGZvx7kOrZIAyWlzl3Ir9Mnn0Z/te7LEeDPGKMP2pRsPj5/hvYqKI/sYVpca
9s15A6PGHE6Deyeq8zLRn5x1p1vNa7ZipJbhyzWb2Fx0cMeb3CBFog+XzB0tvOHJ
YucSPl1H1VnY0BuXnEm7jLbXBhdfrqcRC5tazuAdr6uQ9fiwlt1vo2eWpMjtHxiU
0I96FbviMapi+vdr+BBOCl4u6J+qCLffHMnFC2HZMgUpyGRYmELBqQz4OQ9diX4B
rFfdFIRqEAqkEDXadSw9AYQaKaA1ciX92a6C4Kh2re2GPsd2/K9eSnd2CRTMmjky
vo+UvQNhH0C/+vsC5aMVG5zuFjyeNonYahuloVow0cWeCuFArepR0NrWbCqaF14v
oX2j7cvQm/kkFopR9z2w6uina7lRolH+urameZjDG2eyGCtHcrh2ghiJ7usS92b+
/UGuxIOXx4hpTPll1pVr+LsO0kWQpgeKolgdf182dDEXS1BSsE6SWOp86pPX6wcR
YDt8iV2EKtxVYnHgwVpJrj7MWYQYuAfW6pqPgj96vOQx7Gw03e62o0ZlR833t3H9
Z4TitSd7xoj0dTphk1q0+mw+fMZAveCYCWFKduL3+BuU0sBIbqwrjCQbGLwEmrWm
fEmYil3DT2SBRTz3Mtz1Cp3tWq/EvPToVcjxp4rPW3jstBimWUoSGYtmYWA/PgwE
AeZQ5oaINKyqwPkJjZ7Ww1y9kEvOACL8cfAwwodHGRG4/D53IdW7Acxey7LheTwZ
LRnCY95CuAcfM7SKnMRC/Tz9ADMjDXbedCaZoU9aB6xkDpOjUrErVN8Z25CCRhvp
2dKxU6F7EgoP38cHBQZh/oQ7KkVkmN6xCNT5sXzI3YYnmCB87eslouqX2Tu3qOJR
U8IvVUN6uWriMb51/SXCOhw6Dhecrc1WV6DkupQFvLyhyNpiWXJ0lb76UJs8lxVX
CfGUt5TmOpPsEQbT9F6so1FS1vo95qnfmk7M1hqpYRH36EHF7Xb7zvxpCJxN/XlK
Pv1Ym24q3wwd+x/hMVBfgGBlemGHsPznRX2CT7adm/D2Dz8ndLuQzKT37HwYDQpV
ZMuDYxj+C2wiWdrSm5c9vt6va+2R5SuEezjaYlxOaCKOJqvIE82mnvZvIxGt86EY
0no40SgxXdP6PJ/Cnu0gakYGUIFmST9KX/6wqRds81xALlorlGS59t7qu8Q5+GPN
QD7DwNrKqs1Js/JDcMztImhTXS5wmV6bOeVd956Qu4ekYxfA8C/H94+sRJucJede
3TuhSg+g0UJfAJr45J46CRh4ZvOy8gILhA/Rc+SwWP1bOyP3XEuu28rEqDuSiERI
cbWhlbSExr1H1ty1PzqB9IiP7I1Ip0hnn7rEPT2TbA83r0VkhPOesOvdIlcK+eh0
/60oNkzEKkjXRLQR7Uq8ptKqLeJAsAUcCCUVERJSP/uazLjUxvh5rs2dg2vlaN4R
PDg+ajVjR5eOlk/A0YbEc0UshrUIOKwY//jqkGIQy3f6VNOq0+Xpth0OyFCz21KA
XhngbWTlDDiBs2MeI5K+cE1lV5NfyRHiQFOq//AxURaUSgYiPMUhuw776TSBB5eT
aPIXXf3Den0azS0PPQ0x1w6HEjN70oJ6E3n/yGhd47i9WhCqCcEzh7MP/Bc0D73y
TDBQguR86ZvY2AcEfJ6yVp7MT5lTHemVPuIWGGodQ8wDuv7FxZ2+mxkjOFB3320U
RAFjavq+WWNqdH1JKIqC9M7OZFszTwpNxy1J6ETFFGm6Dp4+BnfLVG3Zgafj4bTI
10jmYJ3zj6wOCjonlLOalQky1tXqaPGz+oSLjxKF1GiWp926/ZoaW3EoN6epm9er
iqiWopctM87K39/f0SkrcoSyvHNWtaxwdbZvoJ3hlR8RaPYkHpBhtUBGLPfCR0B/
QnQYit9LIo6FLLOeSTTOjTpZFj7GohVV15ceSBYaQCZ6eiIwwD1Sz6zvJUKCvuSq
ex56hX+kwYq8hXQiOopUnF/1aEmnMTovWf8420LGd57fw9+YJVl6wSmP1//OHUJw
eTiCTsxrizaQnuxVOqdS1eb96z8v435tdENZckq6OEaIhXJKtHHpKuCJHIz4P1mm
HjZgks0AxeD7htPOPBo1rvB3dSb3GcxlqYVekVw0/eyeWEZ+kzR9icCMXW2hYBHv
kZkmOuCKq+Q7wlhdT92+t4W6sr1tfGziiFC7wvGZAR/q2yn7TTC8CspeERb0m/fh
36ERY6FPHZ1CCJZjy2nKKziqfvU+wdTrm4MRD+kFCWiczVmsDHXMohBFb0H4hXJn
Y/pV57qFFex/qxEtJQfVHdMn0PQEYNmwQHrSk6RGt4nTCd3J+cwmRIpSRwUBtxDF
Y/H2mrp+bZm2MwZh3u20DO8mJEiGNnED01NixveuoV3IwAmqcHNZHVKDp+ALjVgY
xT6AklkWdGtizUblXWTR2xS8faJCD2Rrk999y+QIDKjjnenZ9oL+dTP7Dvp7I1az
tR9AK/nNFVsYG+JS5yHoWkGniaD2PtMqcWH18GfsMaWWEggzQBi87TgwVSBWItOt
2whHo+E8kFDdFqYkhpCtDEbrzPP8h2ID5F8XjbrfReSvKXcpaXdcUw3pLamsrikO
tuy0WPz4vl7q355cWaroHgdLmk51Z5sbVVOHJWLnD+R55zTZJy/MaMKkdfJ1Klb3
RbAKuIacRSvH1lVzXlO/qPPZLBJ7wSK0/rOOBd+uAfOlyh0V8WBKhHuJMqSVceyg
yxQtwwNCq2FX3/duYHabyaUmkI9dgCx/PPoaxtm7VOjodWYmUKwDzivTOGSxFrsg
84/l+S8nh6WHVBXzdSQvQ1y8QMsIo94ZGr4G/GnNy90tXnIkIp1PtHOAm7GEGzfI
uUzPXWmXH1PaI5Ex/KXsFyQbfWo74zqdt+tvXoqzJnj2TVZENmHNUEctcI/E+gnu
eIvNFw+E5UN21xMQvk+M7XnZpPm0A5BSubLo0AOJK4GvX+9YkVgWeYOuczpRboka
7cFEaI8I9Mut/zsH3cZfA2ROmbufEDCSamQZEKHZMc9zkwsSvXtm9MFCBxhEejf+
wt983mQJPUedjGMHXOUzQrQVgIUHQKEhJkhOT2ruQQAFPI1O4dLlwqVkjmOxivUE
2If8FiLPPnwNnH+7kUaFw6j6t5KQGGiYlt6f0DouG1a3aDSWsGnQKnedJKjTmQLd
/8hG3K+bAD8m1rMMB1q8xCZZsoQCgzY1SBuhbw0wqLdaGSfADwB0bBCsv17ZHc2H
T74DBtj+TJgK+ty8z6m92lPnSOe8OW5K+NuqAj5Cg9jWvKANb8aoJKz3PXSLHOFW
VlzINy0IZtsBCpsFwI4VWLt8M+cuwHrZ+AKqa/PNVE2kvlYQV0LZOsK4L4gfJUfQ
+b8NAZmev6VsyMaRjIH7C4V7+SWdkvcscRJM9uUfSYBMuit8SdoelzziM0hDiO0J
vEoz8o5NxDmR/nk7GpA8+rOV9Ms+NL+HPTK3lWG4TmFtb4m3hVznEiz0Z/UrncYU
eIRqbjdbf4qhYtUg7Bg5FoEt7rCOlRpSjfeb/thnRjpLsvYekiowkeXTkOtYEmUi
4ydRWGQFJHCKWJBJ4FyOXTzVIvU79BRaTS4rW/5lofLBzbriHNpby+pwjReDKqt0
91tBMI1N7BsQKL7qMOqT+k+4i3fMHzxR0ZmqSebrwL5adXEhKJFCMUQUOb5E7Nvk
3QGcV5mUJYX/VNPo8N0qqYq+MSPpzi0sPGr95Sq8l5zcq9OjZpFWui5n1iCtE2WC
Vh0sdJTF1uBi0lckujDwx20KBhAqfarCt1tPnVUvFLFVG4TvpouA0knXsuhxWNXs
uy/CltYWRHYGCJbnYWLl0qIr8yl+6G/hHhhzDJBFheDn6urbsqA2FfHy0P6R/Q4J
hWQsiRISpq7KXS/Lf8Vdf/eJlRGVYhvHM5cDtct18lOQow3CjLDt6Pk7fuccd/dt
Fpo8dFdKLKpCOsBRLvb4BwlCcfvBelDYF9JzedUDcESBfYVDRMXV7QNSZZtZHyPv
S3rfoUBH7PO+Z87Abv5HbkJHpGHyzdSTi1wBIIq001eazQyzeDmntNZZIciFxK7U
N9O5LMN6FSvkeWvmAW2WWZUTf3M8XDefRP1rg75/7cvA1qP9Jokoocx9n4h2S278
8De4u8v2CWZWZiW9t8vneEJkN0DZIkiTHfL2Iqey57El0gqUuLbqWUnWHHkSm17c
dcreC0p5o/9jOyw9Y+WilEZ//MGttKgyIr7Cr+YM6eW9F7BE4Vk7yTrGTOZ+SsPQ
0TmxRA0Bn5LGdh39O9eEp+MxxOSnVxxrh8DbHgTZXQSOBZZGl+8ixv6NwGY1qTgM
YsR5dfYi+37HmmOuq5Oasmc3bqwBMM8VGiAYb3lLvTMnwxuWM5mSTP+Kc3+T2dbq
57pHLM/YyOffa3YdScovWsyFRjA1/idGzFmH0zvtTTo7xTQWMxEc/BFKMIeiJgDc
+Wu3C4lt2t1dn2wkVq+g+0l4Jh8zTPOUcoSjuqXfl1Vb7ficY0ia4sCffCS+ZHHK
tlwoM2cv59tDLRLyUjqfhrL2WmG6DomAOtDYnMpaci68Gf9GCS0QRTYUOcvUk9K7
7nkgAPB+RpGd8/Bkt/rViP6NbCH0MYlYd45pVfbd6/b/wbHeybE5/HSeoOi7wkc+
VF/7IxlfRjnkSx+Cxjfu8/z8BVmL8E50NlzjQM4s5hDi4eGQ/0Vlx8dsUGtcXmsA
EQBJaFCv08XUdDdwKYPFTlEHht8+p7jllGmAi63KMjDL6H1CVt2lm093eB6ft6Oa
O3zU7XXXBCRlWuKyup03rnxRhEM+//GWvUZM/3hKfiUgLnu3ZNvJgRijHDE/DLXc
ePOJAZ6ew0xPPb5EiW520DFEEaEU9LYs/bmRziijuaQ5Cvjyv/0s+O/HZWboj1E2
jcYrVcjvikRnZttPk1lzxAwLEYQeMQDfNAJsNjmbJTtM1TC+Jq6YljenXHFWJUAm
o+oFkRVo3uAsPVg7Ojibzu1BbU2IeOqjScm6lZgrac7nT5l9Ly8b1YyB5klY5YEI
dQPomKRrODBPeo9EUkcsbRHyjRhsQXqu7tz74eGTBpxpRp9xlZuug+EV//jgLob1
mD5uP/ZEpjyp9i99iqHU586riI/An4NAhNCIXqpUgQoNhMvGwmcfMW7l+tahFS3U
/8Q+to/eH/27vQxQObO4RV0QNZcxHyO+4GsLQ0ABLXNZiRovdf6BIw8LioQsyqJ7
apBm9tbEL1aqoLM4poSD0wkGx1GXqbUeOxqdsgRRXceCZMbe6hghOh78o3RUbnc2
HfHsum4LKl7p2XENMdmOTVo8NgWT1kCF7OfDw8fa9cymW2sutpoxltm3t487tAoQ
F4ly/LniKTDLd/pBX2nV8QHO9WlvTKjC5KWERhYQR5pTy0wlyOGfTRRJ3uVgJuw9
l3Ic9AEayxZkdjXQYpsAt/3ew91vMvHqrLssSoaxilAU4FoIZptXkPKgw9fq+Ywn
tNk25JUObHgtTJREqXYRpFDPteEE6j4NEzyU/MtsBKA7GftDiMR0XBBuXnM0DUpu
Y6Pdec3BhoN0SdVrZlgkMqjYG957KN4PGpfCq+bH3ELkKEososdz6IzIeyb5Vdwp
4ZeFxhKErttQCV1zYNaUJ6itOL9vFssddr/qBVrinYnZeik/ND9gMg82os1P+iwd
xIflW0jYd0InytdThiGtaceixagwuawpv1I25Nt2EZvohFZ2ajfHHYwbPBx1k22N
kYFPZzwoUVA29N6Vy1YytQEt1CQejQv1IkF4NCd368VcAqDpD7VG7N7ZIsHpECRO
SykCg8MnZmXUgEY85avNvfxP0p5aQSOpG4sb0RulsrWX4XCJOuV5GRahlCcIicXa
+oI9YOnJF3ldF1qtI6FjKhhmNdJfGVT6gHia9dS1nSnwnhU+bDefAVYUf6lKZAv+
F+RH3ggmNbtVMDe76PE8PBGPwiYgaWanTGqvYBXsUSFcgIbTbMtit7eIzuNlH6x2
ODVcNqVHDCKvevlaYPoeHB0I/+yf6RNqzmEH+inON4Apbf6+s3etP3YDfCRh5dRr
/Hh0GVva7LXoYWIPokYBtvxYcEXcgAGRqcMFFSOEUlz3rsjmrQKg3HYP0yOBNNIS
HGd003B58naxI6kvjfCR93FOXSUeC4Yl6rGacPf1DmrjJIgJ4NJQ4tWpjTCZXsNp
Fr0QSLZ/uYQdx9H1x8sSX/7HzbdPTJMsMz+duwjtJdEwEaXRWo5ABBCIFdLRYm7J
yo0KaNbkJNyIpecbZgLv7Jh+f46hDqrPsf/0HxnFoKKFqGjWv1nJFw0AwDCrgSg1
y8C2QtGYRjNYUsx6bWHwj96QBPTN5WHA2m0JjMJ0KBnnlB/YQSwpqFgrqUl7rE/V
QB6xRoFeKvvKGDeEM6IvrWQybw4n8KxSldiC/8t46uABIJ1MW6Wf/QI+VQqJq5MN
aimQKhp9MZjFPl5etofYaP/uioxrrRNqfb5/pm/kb/UTKPGr99l+SBoUmUScf0Zw
+en9kZflpl1bQB7FodHUY17oORU2rZAFsxVp/Kse0WwYt2m3pEleXFtjaWH4BOq3
7OM3GveJ3iR/haNM7YbRSxUByQ1pAaXPI36jCaWiTlrCV+b3YrXp0NRLtAijj4st
uh4OvY6s09e4sZdUd0XhMJ3XtZpIClbudwXiUEHtisuAxql0UI/PeRR7JIaaYKgn
IvLtU0kfvQbNEE00+TB6GgnVvZ4TDTuMzclv5pa4MKnihX8p7UToKBXaLXpC5dbp
XBjpIQtgsFlpjaeCCcHw47e1gOZ0iyF6gRARdjx7dowtVaQXR42Oa+ZElEXwoskY
XrPEEfXYDgWA36l1j9dof6vJdsGjHVsUQ1gIQQATYuj5/zzt5DHGtEW0mtbhNu+1
Hm/Df9/RHt+N3IPXTqU4xrX6oXsEfW2ynd2YUHITKkjeepgYKoYFnXZk2+pyBmMH
vn26cq1+fu9fI+8D2I4lsICapd4l7bsSbhOv1DnwE4rupXSrw/YG++WWXJ8xhXZm
DzhgCbnqdlIkzuvPeUqbApIlWhEGONtH9r4rGj0+V/nWRUx8uy0Id0JHMFusCv65
dfb93ftB84bJ4MQY7YJqwRSKYLu0Rts7GZakvg9/1GRknfWn778SGSvLkuPGsSd3
pwdN8XDOJNICbhTOgDLs0vlouZ6Fplq4DkuuMtlhpGiMf6NGStzruwpsZTMXS2y7
BKl50egqw/pYAQoCjozgzkDAHn9TNI4mItsD0D1iXYqCH6mQ3qxk6NTtkwyIW2hG
Fk/0+lwvstbhpk9uRIlGjKu/yzXgrVk1qVkL5l8UwVRpVyScvHJdNY5SnYIDEOqf
wvzbaMgcMrHnWEB6QIHsEYHh+COS6TdJCgycEpvVfJn/nHAUyMUicGhWnVi/O6/h
RsoF26sBznoUvsqHB4wOnGRMBLCEiyi7Fxazuo5fWUQhcDSzR1PhCif71mQOgPB/
AQ/bzFS/SPthvDA/mRAQdMOIslKyaUQaL+17GXf7PDF+GZ0+Qa47rIMeXMQ9xWaV
oP0hxw9QysssIbq/R2p2arTvSnQJqvNhETjzHiplURsUo7DPWw6OpFM4anQRSba5
Qcjm0EiOQGFlgJeoZ44JDteW0Ndns/FMZJ6cL4J20a3dvyypMQpB7HJCXWj1kPPD
oIf7lZNgsVzmHLuGEcYJfbesoXBrOJmofp2+xbyRZB3V8XsaP5OdRvA4lCXiAgT5
TubCGujn0pIPqKnDRBJYDye3utblGrz92/mfBFV1WfLFzZRkgkxs0V2OxDEn+/U0
/xsRAgi8SOacOagn17EZRvtUTKGZfDN03Dp/x7+Su0CxzdvMNQ7PM7hbOczEYDR5
agKGI2HIQveW8TWuD24hq5A1Ep7FIu1ZZO7RGCrJJy/XxYp27fWqfQiYx3nBBNGd
iH4ORd6QorLNtybgRzNYI+iX30eRtWjyzuMp6FNf6TDVhwachnzZqCJrsweZ50Yt
3Cp8QbDCyMD/Pv1AINS6qpdtV9xvmNLFud9VHhYrFWKo3qjq+smGtZ3X/vPxNKEx
CbHELuGzCuUbPuza5x8GgoILLeuRVthAEuI52GTJ3yCtoNt7UQPpgGDbJOZ6akDg
leH7HbZKg+M5SSXWzdfSTJOx2/CUs4AGHkwuOOBQaxwOYeohDgUNmtv9E0VWpFVS
X+U1aMHjLCilgh4154mNPUXG28JztV6osqVrFy84Mg20wjbldw/82BaJE57gw+ME
E0N8wVfpmQZkHYU/P/p1HYMo5v8zxcL+zfgNNKC9MB5wA5mXgJk18dnmPyI2V0YF
xwIXaj2kIge+xqEJecff3xX4EDmWTSS75Z0UckOGS3CKPjAlccl9ubZGcdh+Kumu
YzsdKpobIlKXlNLi4tMekGBMLGxn/UNIUu1jT1T18FM3D0Btzej90GMGkADNM0K/
gF2mhtoHunzdA1QQwoNlOx2beXzvUbZfMyq9A1NVvsb62mzco6mnrYcSBhJvkrFt
Dy+G7wx3TUVn8k4O0JMJ2r4BFcjaz32J71xyXWWZNqxkfudpkGjgw156K+lED31s
EGbaikhC3/qaQf6GGU/AD0nWep7IilJVNASdtz37iSWyHvvwaIayIVBl1iFVPTUW
xVr3phArRf9/T0RzpvSKaXWkbmQdnbdt3xaNJjA17yWuOU5YX7gXbfksbxSo3xV9
UMvNt+NuZSi6WByHNtSycwapEiyi9WQHAo/UwDOE1hHbuBesRmGNTPBipTNm1VLn
mBZsSp6K1PGeX9e69uSIYTU1b92FwTXLSJJGACb+MYmn/a4Eolf8+vkfw7xwKudM
FaX/anyGGEYvC+S88XjWpZ271NBc5ri7Uwzck5DWoF0KL9PvZOMy3zNDOmm1uiUP
mIOkDGus/mxfSPG+R0kcaBaHh7GLTTsUUlhZN3PwPLggdWmV3rFlREa8eIGPxMNN
WWgTzSAl6zvK81xX603MVJ4lglMcU1Dnagu7hSi7DeJOkebWuSTxvMKu6WQf8bgk
C02kBMcK22u198j1pDfoF/dBt/IFPQRs1li11SAJgcCOSmjdzl+T+7WTl3R98szr
xmI5lqyC6gLikJf/SVzOS+2WZWWfSwXZ1NvhP2pdsBRQO3TaaI6BA1xXmNJJJLJU
idqucTDgAMrsoRo8xehRk/z3obTorjMGnLwXhO6lolwLF5SEkzLdRF1cBjCQ5qB6
tH3FmDZVqNTYZUHSzZ8N/o8xX3RdV6Nw1UsdYY3OcmbSDa/qlNqNnn44smzCP6e1
vtErla1hHBVqYbXhojXPvxgtuYjwEoVYOvRA/dMFaic4wmbeYhCbWTjpEpK/Yk27
TimZIJqNU8SRx/+TqXk0XIqaxUFsZu6yRK3oBTpwZnN+0BJahrfUEhd20kNnHTiS
9iUn3gdOIIIwpK96PaUXGuSoUNyNoNvky7nPgb1CAaFELNRUP2XgmOzKeWRoz9+K
/vjeI7bVLIPrLEXHQJkg0MOsdplBGKkDLDdwZmniI2azZ9AfQ1nyVtsXYhzPnOQ9
GtF62gha8SJofyS7wkrs7d3RbHUuJ3RTlmLE2PNTol1Dwv/LydN480cpxSYqhjnl
M2st47zxCXD8NnxrvKjvQpSBN6l7yEN3LpMnlPb0xy0GgZsjyO+xE5RRMF29fw5s
h8QfaOuN10NT6WKlgaIWOZXCGrRE8/Yy0sqNYB3SYowxNB+etyKGJMEDD7gJaV15
/pgggtjBwXoAAD0wDxHTlTd/qKyDtW8bfnsHjm/qaoaZZxfp96o0uj+mczNsSU6Z
odDqdj8n6p6VmZynXv2rH0mzlp3yHv6pKcjudwDsQHuoBPJDhZEpD3AwDunIUrix
c1a0B/nG88lbd2kbrcb3B9UKGYU/hTGyDV++Di1D2VPa+7YNsaUccGO4v5KUQIpa
lrA9KeYpmXdOhVPF3y5Xw2vr2q7kBRQvMC4PEEs9cebbJYcbdub6/zWhTGfmSIIr
0nFADniHuyS7+Hm3BSgIybKoUhGKXIo4D79TrlNGMnZA/Kdbw45DK8YSqx3o4GSd
954v/ndxYPqWYMYxv1n/KX2mhb7xKE9ifx+y7mtusqOKHpNDQHVJUMr9qqDQk9d+
mdzE5IdC+v0GGLrbbLWvrGei9/tM3y2sJV5fRQe9iMnbEl8SpVDzYf5+/G3arYdr
QbdFl8bTZ9l50w6SxCaOBTCKMKI5B2j/Yl28viFXLg7dIJBeGsBkBnL4PI/k8xdO
BftQq/0iTkCjlGBTa8Mb3IioiecaNL3CFXCDxUIen/SqfI83lNz5UPOljahLSAH8
VMx7qGz+zHAsafsTAtsCGXhnyublElDeFjfZA07kD6QrCDwMGXDwQwXs5+i8nYWQ
dTYfwpGqVfK+vHeT4hGxWyoDJC+WqJQXhq4BvzP9YtM+Vo3hq8wtEeqeKUQZKDTY
pxx5W0fxjl3mMnNT/8H0bXjY+wtgowmIAyGt1VQ0/68OcvRMAegJco996iRi1DzZ
llirUMpaZ6ApjX7WnTAKwFXBbDKPL7BeSrRv2zeDAojW3X6VWQbW6eB5WLpuqxcL
cu/lvLsNd/o9pvaaL45HksVMevghursqqqeEorAPWXSWhZ32mVzi58f5GN1oX9Em
KcCZx3jytcU4bhxFRg1v84ePhxbUPcHd/lK7VlT158H61ymPttaxqr+aW/T20Qqy
ZXA08F8Ect9ktr9ADcaLzEMw4H9Dd+nt8Zl3SqnCdWX+fy262dCURAFJ0WhEBULf
pmks9mS6ak+Z+iF4V7qaNAq7RLsNWkuKRdt3j6J2vnLJWeHud33fqp0avaZwksbS
f53NRIlsgPyi6De/yZU6BZclA866WUkdbBVJ+MWpzO53eo+rGeOuNLxm0F9S87bc
LHQMKDkOxLB9htxZpYZ4sgfTh9gtl0Pejl2e5TFPOJPeR9dSuL1QMkJ8towRUOd5
V28BU6RiKE2D64XySeziiUNGFvxtNC5WCEbbZZ/EmOmFJiYUbSvYizjpY4fJNodO
cqrzooAz6abizZpySJEV5DxjdnkzythbCzxdWeD5k6rnKSHB9ggbvcQbALHINKkQ
j0yx8oz0Yy0X3mPLpQdKXqDM8nx6xt6lIn2a6pho54+lGnPnmKQLggRI8HCzeslo
i/60bAayYGDtx1h/dz13x5yTVo42miIPyODue/9+iI9qC564XaX92Pj1upIBhdv3
zxHvUBsj0FDwAYkShXo2GDTw4zOtG+VKR9nO0YLXsq4J/PmxZ5Zp6X7m6oYQJ8XI
o6k7nH0lmcRKg+lkWRCl/IV870vpUqokGfTVtsXK4cp2fHt1ws0Dg3qmDlYCXyoM
kSeqfl60Mhe+sJHaDm30lCFvmSzeOMh7cmaz3qa5zXajxYVQG9vu0bdbb1zuoA+H
vzHwGBArrtfOyBNkN/yO9mSg4SGhf6AURDLRNmXgEKFFGioD8q9tGxlQoQA4qpi5
cCnSfeQXtyWhvPzijwFYDp1PKsGQlJc1U8m5RsWxqrgFhtAXCnRJWqKiUOQsd0i5
aM8ClVeNCe6vblO0QVqEJ3Z5H7g1Nhh4CtGJWpGG0TPlrISWODAfgnYLqO7l81oc
KHeNOOQVwTA8NGSt9tcIo656lUg+O+6iMHVQCcy46NyG0O576VXVKN81A94pCkSk
PS5MG7ScpBKbNFWLrnLb7xMjTE1ZmpYtY4XHH82WzICr2vxrYz8oLSGWu/Q+w8l/
+9irBxYYX3kg4BVlk4VHe9ZbhPfo7s0fgUWlcQPuV0CHaH+Tbv6ePIelCNja5cso
LSieNEt5JYVggfiya2APUcrwRadHacYzwaKfk/KH0u6q2WjrMIT2eBwiS/vh+CUB
qBdpJdgqykK1gUoMAdIgY8KrjgcL/9qHPXSNwXXldnaYRjqNtQFzcDbQnFnnq+1m
EabI3yGpPOPni7XvtElOTG+3smwcUXQqwH/90cOC0vP66xXR5sQQbyOx+PfseVNi
UeSLThPj4b0Phmff2lQcJJUcZ7e9JxxyRpbjDgqYIAw7mj2jd+G3tPno27S1NXBL
GpCRiFa+z8G0YRprkbSKltEiGeYTQE2DGM69Xq4aWf/ncdP+J84C/Ll4up6EYXK1
LslBqywcJbDP+3FnNwxitf5y52SYLaWpjR98C5nLh71F3+FsI5Sl5wpcJ5PqzXzM
kwHNwTs+F4Q5qtDDBAeWwicWs/qZgp+45tprlDNKShNK4CsiUHmBPEhRWmnqwmC3
7hvOa95TXOZ4WtLUjE8bImgBPV6sQEUbZW6wJ4tZdO45Iqr9n3nNi/a0bW07d4NF
SL/2jouItmHYDc4Av/1Kn67UC0L4NVhO8rLm1TdW/735YoZAA2ysUALMuRIt68EL
dqweCilcFiETc9FSn6WaiFB6pjibYUQFs+S6xFYN6+XeI/Mia6QQwaqOvvaRvEyh
NbX5i+o98HGDJf3/PY0NRTso3SnWarEmcGLd5qg9JYrnpmaXJ4Ksn69LQj8UrBJ1
Qczxppa+qq/Qw6kSrT39MbfO1f1DkiFDlg6HqGH+74XzLmvkaWH7XlN+G9LoCxIO
/Mco+ft6nDbFdPakJHUM2NVESYdQ9lsfS7Y7SAYBV+Cu5SyQmAA9FwX+8qr/P3KK
R0bF428ed0xuc2b7r2pqAbsO9xq+zrsNjyGztRXQD3FIcWS1lC9iEJ/BcKilQcNF
L9LkWDHCkoksHCLt7j024aSpUp0HGRE/xN7CDOQgfZKATA3gh6sL64zyCKdmY3kP
Q0xl5JIkQ3QXP6s907+RtLYrR+4/zpAZ/1Wg3nDiZ4I75zv7byokYcDzInbVyhTF
XbzCHaDaYUa8gpsb5s3FEhY0tO09O2LVuuCz2SJ7ChlrQkRXVAj+rzqefcgwQm6D
tWRrqpsAllOD1mGIMqkA7ALZRIvpGgBe6sSyKNlO6zI8ZsOja6QlKxBh7v4/vDQ4
OgfXlJAZrbrfFzRd0brBn3nR64NaAWDgzZiI7NkevYzGObSjTsYsb+S6pCi+13wq
vwVeRCg8pEu+z97InZlBYy9ae1uJh+LupR4SUTX0bBGXkN5uzF2unv/87iY/vUXf
PIwZqae+o9OW+IbErno5EqygS5+NyWu6I3Lq8AYxx0X5XewZPZTahdyuPUf0I6q4
6ok/13bYZSpynNgG67FdN4RfMzHTnLYw1fi3TAOgp2piGcsmm5N+C+J71CYRW8Aj
Uz/E85Oefmpr65lINJd/pStXQ0B51hfWThVd397/2e05zNhJ8nJTmO8f9TuZDOZg
T1olDPfXnMUx3kJ9fLRGcFwqqP8GCy7eykVs+AN8JK2QWwhMPipF5MGGZUzheA+c
oh55VtQPrT5cp7nNoLCsuOsbmPzKuUGYpGWhR/mhqPiX6fROImud2iNOrZnKPJlk
mLPK/ldypQcPQSXzOqk1WzJN4hRYd32X2x2fj7V4+hO5S0mkke2i+ABsF0t4MACx
0zuT8BvMpFZDEj1lo51Q5DK2z8pk67IoB2H/86Ioy3H+ISaiYbVxkSMblHrlP5Ay
EzNbcIUMR14eSWyZoTAmNjTX92ZJHx17XVBjdWfBcKTG57JUoX5b7KnNdbxffXTi
YxGScyGm7J4xMaalxjBI9u+De6ldZyV8zp4O6q2ytSGJSoV1DtajBhPniTt5G9Oz
FeONyKgdZRZ6q91W0NFcpoelkUDh5Dzq4wWEo8Ram4E1BC14V3FXYBX8Df1nezfO
mmFS4LtDsvKiUBgjy6AjqtnWXtabyk3BWt9UpbB8zP1X4Z++SUsjoWmNIrzVKM/g
w+4RlgSaj+IZ76dE3JHU98eddqZgrlFRJgheA2zpg6jpiwHJT7xz+22MCHVJ4saI
SEVP7rLUb7Hrz7nHSZNTF4i5MWVABjofuYPOCCG6K0Z7mgTvJBvliJkwoH0GnQlK
msBZQjsUuEeF365bLyNQ1Ffq5juX9e1AteLFRBMG6muEpAdwAYO4K0XKamJtKF58
P9HxwRhoC0s5+icAcr299Ik3SB0OaWbWxayqw7jDgGX1J16U+w/BEeAZXZo3GkU2
uAT3tB8EbombDB5Bg1N9DUsgTdDl4pJWyyQ11ioMsJXpIhN3p0WUBXMtOod2qaTB
KHmug5capHTQLf0lcHmDe7uBSgK0+Gu1TrGjU7tdt5PnuTFsXJKs0CDyO32bJcV9
y0z3lpNppPX0Z2lTEQRWGXcaOsgdIDtn/7Dspee3UOQ9IDSb4HFUnMKGm4/ezWaf
o9kDOL91bykiniXNI0/rEeoepRfUrgxu19F15LJqF8tSFoqAPwVO5ffVhjo5MuFD
m4VkQnBBVd7ooIc6KwZ1lsTbx/DGV4sYDTPh7xfNMvE/lxMb48CE1LFBpBFYhjn1
PqXwp3NeUj7gbo3xola0v3UpRpkmD7CoJE6HkBAxGa5QDZW3/NJmcPEd0Q5tMhHm
rlBwpOPNtyD//zDfx4YdoeEolnn8IWAqXrUEhx2H9IujJ8eJb23UkTav2J3iflQw
V492l/IFa1d3czeTU6KkhWuXdjrArzzcl4yvkMCmRHajdkHZ1Uhi8u8mSCiN0Khb
+PLGmbE2XXbIEqXUxgKI0x50ca2dEf3n5agk3/oHF537QfNWC8NeCiwsgGrGwFjs
Ltti0rGh0BoltXCrqcbAcV8RKLZH8WBK0cTeQ1aTvPAjHgPtSEMYz7HYhN5d0qBA
dmB0v03damswr6kM8TGtbkLnv6kkos+pIBK3wieWeFO68nquMpEGjkXE5+D11v//
bp0wAielvEqodJ5jCI1ZKy9Q9KgRmWkXzSUYjHtMYI/kEXaB29eL9V9S7Z659HMj
FjUSCJZE3ct8pBHOfZoOYPtDJyTM+5Y1Zfzz6x7n3L3qeKgQ0NKwPCz9cQ/XAJRp
rSzYxTwhOFm/HvdqCHEzHvCeQdV9AvJ1/gpL0rLGaulhv2FeA2wmiYI8W50ANusZ
iERQRZ/DcOhx6lMdpiIgzZzAJ4r47ssfjUteFBr84y2NZpWV4vFbjjax7KP6jOxf
cMVKGehOLPUDKGLu6QEKz6p7odZlvQJ7y36ZZ1JuuL1huLJwwdkh9ZobRP7PHYw4
uJOqDkun51XAYUiYNx2HoTHrU2DAX0qGgUwenUI/eVhtcxVPiPpyi+5krXnL3F/n
mv6xMhfvz+GwvhM4wV15oAgN99rl5Uku8tuP1NZ/UOxvFKKvHYvFu3aqBQBBBUIf
df05f5nAIIGRl3foUWF50cSThGVer2/HrQGksJzNP5beacxNpwx16VD2LRy5HYtN
CqmnxfFoM/5/SlyeG9fJp8Hwx/2xAD81dV/RfxyFWg6+1T6aID10JmAkQhIj1Hg5
P3wbbtVNycNa8hjN1jNNhUKCSS9bCpgHldQBXrvpmY2Xfbx2qyV6Ype3bcKsJF2P
851wJOK+sx7Ou7kMH9R9SFHe9hnPSaTVglOsjHX9EP5ZtW9CzYuCmpLcAxl+slG/
uWh4gPeCAlWkr2LxY8MFO/GR6rRArvaTpHTSJUbIN8GZDLnsSYlD5vWJFio25qkE
eidxwLs+6IqN84SYhcupAA965iR6kSIhnQBArz0DQXv7SkRhtAtv06zAEgexXxOA
kuKYMHx+xHZSXYjJWb+4wAdeJp36n34OOhDU/WUXnmyvgbRz+gd4LMcdHUP3i0y6
DjdVX+lZHoGLnwxdHPHGomv/8l9cvxE/SzCZbfpyXiOQecEcnUPqiNy3TNO3HuGS
Shzz+g+l46Bdwk0SKfb6WO/UEII3Ba1cIqqRnh/ZYjjvLjf09X4DMyjTFEe8aFc0
MRP5DntDbxKULgHNxN0WitIIZelsOXeHrUoY5JeJg4lsAv2B8vLO+SA71ikpX0sr
gPMvarAPA1MUBVSJqFvHW9v+vGmreUHU7gQ48sPTBF3AlpGgY5ipmjV3qa08tsIU
zYGCPUXaoxC7uqg/rZDQsxrkaQZYEj/mgYcOeah9yn4GpQ2mM2sZ4ETOLDyWEBs8
AFdE/RrjDZGYfEdtgv3NgXa5sggcs25bA0zu062A9VwI9CZvP/ZaUwuYblL5kuu6
2rQlriT58AfD1I4d+FD2npxdcfU+n5gOOvWwCpivG/qi5o6jLEq2oulCeyt5RY46
m5GinZqLoxGgZLeZeuzP4YPTWqgLJS86UaaGOrg33t6bczhuhV5kWL12UZJq6cB+
LnGf+KWJ4bPCXDOi9Yg/WXkro9Zw8tAZo44aFfGpm8WJQacbXEX0UcqfcM9Y+jR4
S/t5YIdC/wkC7T5MZ+MvaNA6/9STXlACwgutquXN20x3WUT5oOr8La1HEfEk5dS8
d6KcwKJRQTDHHMUty65KlDhhCjopo34YRRlztdTtSmJbVOt0qts7YJhVVRoYXRZI
Wob16hnIYcAqJdzdvWuMwjjIAe2tdtwDxiX0rHhjlovTzBAbbbliecPCf4QbnGVj
QOx29ysDla/N7Fkud7F6dS+6roAqCMOXAXidErD1BHbeEx2zlK97J4rW40vdriyf
NcE5M6Vwz8LEKYxRUMftr0L+SyfFoCaF7GxzIBQQ3Z9qLLzqWcMLJODiTq+9gFGj
NdkgC2l67jarN1BWj+NUAMgf4g+9xzr9GwIq992dvCjvqnTPiLnJpnI4ZLoR3sC0
MEpIaFpjHmswuzzRipUmrs2CSHMnNZQ+ZMtvAuYgmWp4vbU1E9hDfoAmyXw6A0uj
X97jpKTZ/HRTvaqP08ZaghwGRFPtRLBxYV1CdnKUKb1dlT3/3EzL1Qg146yWgKWn
sys45nglLmHa0tsrA6PP0Ea2+KUaWqzOSzqzs/xZYS+fK2j2ybp7eyggV5U8Zc3M
Sj0UxileUj5vFJJ5CiBbUCyC2GCniAcWT64ainkPchlhLIumVlp5v0INAcfri4cV
WzkyrN1zG86ILfuBI4VMlFAER4a9hvCGr+3pEfvzGkOn48g+EPxF5icabE3nvJMQ
KVIH6xmPXss+q6l2NzLSFLJ85sajSozyHrUc+D07Ulm6Of0gZ1T1uxW0ByyMjri8
TIoxjbJJQD5xhcaaq5vFeGkM47ADCPgf7t4PNe5n8CfTC3/oTinEq/ClBvZ1VDva
j40DTWgGWVqT07j04CqFofBeOkMs0Zxcu8RsmLb3omQ9D4kkiiYxs7r6qdXJubn3
OMdPQfNatrnOOz0i6XmGmgldatKu4Ax4ND25BG4Tx0ffJxouB5rTjHEa/4Egy6SG
uZHhb4xGVGxMV97FifFtc5KulYeH6K9YTyqymumoxlL1Sh1MkrlWnaW7PXZ+R/ev
kHlPPNFiwDAb49LEmEqtT6VZ8R9cGex2a1BsGgTuJt3w7QQec+w+YmpbxX5Q/AcG
zDgqA8yzOEUdnD525F9DkPTmW6q4TH4rpJ3uBdIJRsftO2UAc3IOEPAJsvQ6u/Cn
XyrXCkDPNEA0pa+FyfVQW9QM2BjD2Zqx6YUK2PTcS630qq7TJqnzd8xM2u22iEKU
iiWesE84ao47D381nDLKP+eQVtdVU2c5RiGoQL1we4svx0VORwXYRAM81ZbbUMhq
BNk7O6vXImspLLQnU3bxPnd3LDRZ0RRCTilmuLQ/xS619Y+SYQ5F/ulN1co9AvDv
7VwNjQrqVWJWDTS3J3d8bbtnIdUP/Leke/bMTV2gDJ+I2BIbFVry0bdfxcqJWD1E
amjDzDdbr8B8bP0uzuU2+cbsLTn3q95f8X1JsZQt1mn6FCl9PXYc8zCp1wVUVGVy
mDQUtfE+0aNMzRykqbxvvUcglNWr75lxeIdEi/sMfjHM5WOvJZ09oU85P0TVIHEK
bN+iBcYqOK50GlwkEWYoGC5cgxF0t5F2fFQ8AFfS727wdZP5n453NcSygWGwQbR/
qOSeHYOA1qCofR4OiBpAtJXeQoA6JxBuJhDSK4GSTmL6EsUQ0p7W2te/gA/vxByr
QTp7Is4cXge+RNCzxIasMMiOiZwFluvqU9R2zGCyIhEtx/eZYo+rCs7UOjCLrPW3
UCJJM4dZDKvqn9K9eI0aUP33S6Px7/qxAdBael8UVu2TOcBEofbra+MSgWIQEvvn
W4CqPridT/nbFzIdQhPQIBvxEEKVpALmNVDNBSCnXEl0tZOu80Dhcqx6Ys9I1aLi
nSJYjJd1HftcnBYQIeBxGuJcAgHw4HAWdJeSCGOmHmecy6EotQ29gK5yYrvv9TZp
9nGMZD+jWACsQK6a9dz3dDv35hqZYUIyKRsvnlXcjzOZPtX7V2n2X7EYFfFcwEqm
EaNNMEMPo1m79zxeh7k00Wvb5n5UXpAVS03Ahd5fDt8oh6FS3Dt+S9rAGBlbFWaD
2/vhr/QgqLGsIoswGGaWLbAuD2oQHXDy6RAxuMPd1m0sD/wmTkmv2pg9gEv+lfyW
hMYIS2yIK8NAt/e6vxT1e1GBFUsIPvjWc2NtoUvquVd+cWg63S9nTRy6hAgz0GTu
JpH88VpjJUmhb5UEn2jZJX/q30esvukxJfpMrPO7nXsUze7cwTcywDj7U6b4trmS
fdFNVKt+APHZYuJ0DzVqYeksyX70rZhyZZwXstZonnekzN3CzSqvyIjvXRtJ8+hk
iYzHoB1tnEiOU1a68iDA7pdF8twZ58/M35NTY4homumNKBie/oJejocuUNv8c6jX
HUJvXyXUVI2sa8eWPQZHWKWdgHSJbGbLJREpyQDoaF2wh8qOIm+S3kzAWaBAI/Nw
Fct9jasJ2km2X1j9vDl290X4wj5pxwm9wbB+uas2G67hJmq3/ni6fyuppmasIxjA
bIATOJDvtAorRwXmtoeksTk6DiTQrlwLJ7f2yZE3380q+KAFWz0J1FAkL3VkbPtl
qlYhoE0PFboo9rYuV1ICnJL1YbhBakny9seTDAw7zoHhUeYJaRwiSZknmtJucyRm
klld422jaxoCj6naqdzgRpYYHxyvGE+LSBYTLaPzbZCovEqhmvaFECO5C+/yA7aE
COxZGPtkc6kvaZJPY8qqiFSz/sgvbJOm3nTOxbzUAierSofCe7zcz1X//kEAdG3X
jv8uerpeMdUELhBGXfBYQuNnU4Nv/ZKSkEkcfAuMcrwYdHpfBucUjRj+qeOZ9JPf
fkvO4kstk3ACCSlFzt5WmboOl1GIHyJjDwUkIJVwr7u4Ex9LsHRILFVyJb/XUoSh
AIrg30ObyjA7q2wwqg4OU7/L8EJawqZ/g9nSTnWt0U1ltAf1tTEzWArJ0+LtyIXD
AMzswmMuX/yGMOaPLB+dC8XP+yN+JuA/qw7Dt2QClqdlNJGhbtScyjuNvTnWDDHx
goLAIsd4v7ysLudZD9kvmhBCTcNUj6A/JrfhsI1iQ7j0H7XbfmZFhekoJXnB4Scv
7/5ORLUB4M/nct04lg1VnvDwH9f/248WOG8Ez52O7FKDDMunuh/mMjK6bvdRXVbR
xWaxLJdSQ4SnDKwmHbNorhK6cCz7kuWkibsNraWAo6qZF/1sniYswbD5h/7FopWs
sP94N8DqJKnZM9wJe7Q3yAHtShu6w0sqPoY0qyPuZY75/I4vF9OB+mv+TJTzQg+D
DOk3+sCeLaW7vIdMIioVx9XBrRB9HIFw+f5BD4Jpg14zv7CkNSK9sYdiHESWGS/Y
iW9To+negy3e+xJhMmzNe6mB1bmOx/04Qyw+3oaFPF2pAnUFURA35J5fRDcCFBF0
KfZtrlxoub1eRkkrBhx/rjbajBLmtBBGKZUVm/cT9BkX2PqAr90V/J+LIYggqGv+
eEDwAXUHIKxM2dQJ1opAs27P874lubTRMuFU3O+yUMUW1xiLjyT/DDE+5cnWGf1v
I0YvOJ37c7z34caAkRpHFZ2hPNJGPfUjNLtGqmMaXMgF08bo42j8EM/xgrbNaKk/
kcD9HI+tWyt/CsBV0xCg1Gf9zvNEyR4ciiahDQonGQdipP0Dmv0FL+8fMODU9XII
ky09BfGWfV8C4gQ9HC8R/ERpNOnVX4pbxsOfZWE3ETygZsKl6edkUQPBeUXXszRq
p4CHbYReScXO4vBl6os3cYGFqMxJSydvVwJxqE5ucm/c2pOMR8XqMMXxtPxy6kPQ
7+v4lKCkPxI8lDnPir2j/W69AnzW6UqMrXbGB26yM+0KBpMlUMhdTLP/bvXOHHgD
ZR8URNpEft70+pil1Af7K22lawEuOkQubHrhA8OszhNBsBfI5xVo+lMVtDGFjzHo
TXu/ry8SiSd6/79gh9nrfUEfZ0W0qkW4ijolvNccsBCfvHdDei3MrhyFUZVOaQo3
KVWBu14a4Fix1mZa8Yjq7jt9DQfS+bF6UQaE7TFWpyXe5E2gsmxuQrSQJZBPZ4gf
RZsOA2E0UYWa72GFYL3ZK03YjK6gTur+yq8lcGNMGbn1XeCj+YY0OsmZFfYExt8E
Jy1NvrU7XD2QO4emUAF9Gfit2JbQ8Tp0feWLTKURZhRnt8xrdLeWPQtau60cysfY
Ru9blOyfrP1uIILV9xYsvb4DLH5XWrLov3wXjaFHFyBOh42efTLyIRwIeemEPC0j
R5BpfEJhZFdWODGf1SQHfv5BKYFzgBWBkkLyigzhdRjkKC7PnjhcOUea1QUKlABe
D59C7XwlQCcU2pWn6SPb6dUSVqc5SQuKTw0jkGprmDbL8iL43OuDBZDeCK8ToXfG
Rw2C9H2FMX2uHZOEdZemU5QST1U3BVHYENk4/EYsXD+z6D83c2EOOvj8vWCLUedP
wvze4SzxjEhmJ28QlaMHBAminNu0N3cIPabg/boDIIoNTdWtZbV2Uks5P+9BnOst
u4da/HpjqNddRio2UVHY5Rk6o3o18T4OmLwc3mINepM5aXyDKL/M9oyGWDaIBXXO
F+EltYT3o9v/RuiO966HgblaudLpvmbYYySgXR7txtRejfLF4Droguifm1diykNj
nmfZ1wKxzttnaVMkIRpENtImXIFF3s2haeucWyEvtkWuIic16uUwnFEK3BELT0Tl
bEVo/P2DBK4Bvnlij29bSFzGMSR4UIMw+UHbLfmevcniu51o9pAV1RL5L74hoxa4
k+c+irWtoYQNV6CbI17onLm/iwHK/xfFaotHymWyAZ9MdOFNu/cqprxtfvtu1vdu
bjrhu7g/rSnxUTjQy8XbzUVpdwTi6iRKMimXH6MOZMHGMFwDyHBBJnLzgeKL71dj
e9zJsBM5+9zfbA4TBbxBbukfM75HOZjTtwxZa9mu1uGHCz6HNs7jnrVf+KBVdhwW
ADs8Y7g/pjSERzJNdiayMCqwBZuwb18H5R7lkldlpuT1y4j6buGGp8jHZ2OAspQl
eI3jOSOUV5EzFNsclI3AWUut/MLL54mvPF/WrbAB8pSZ5cRP30mbVILIqmmxAp+h
lUjaqe+azhn1wYEpjduysmea/1owsKIsPY7RIqwqWblov1TPFZcQj6zXl1E/citP
I6ynrIaztVWldPePTfkYkbzuu8oxyAw+N2t5wEvAqUZtqtKECHrBQm/izEe4BTAs
dodRs5oIIOpIEnCkpwqUP6Yst5i32zPpSuhTp21j9vIeyZESiAvkaIwxcHJVfEcm
S+HhFwchSwG5NfT12jJ3Ki8WRKY0M6pkgsLP1BF8wnmkcJRgOKSYIBMEFoy32BZz
QQfGVodHeF5J0LDchaYzBsVHJN+2wETkSQjNWiyljpt8/xNC8NHjz0ddZdAZBfYz
2NJW9h2MDav0sbddMylYr0oTippH1aHsOlF1Q9QzVtzVh2wJrJHo/37BimQHTQy3
KMgKt44eMA3HAEvCj9/H8lJQES0OjzDkZDaCZNF0/7RNM8T/veF3GZln0dkWFypq
Yl7gQqNXFXyDR4/wTkpWed5d8Agu44llO22QbVcqueuBSAP7CvUfQ5EPoaWcLl18
oCIqKnfizCQpUw1a6OWABrjgs1D8c0SuxtaTJiyZbMuguniA/K86qcDmAVDtiCh0
cB720SHbqCT+pOjfJdIAe0OH1GRhNkli2/OuGEjuWBo1ojgh4R8AffH7H/zHOtKd
hJqgxKLYRga5sXp7okCs50/HfPsLn9nRtxuoHvgHUIOHBzOWw/P12KQHK1yyAUJM
QLCyHjFyIrY9RnMGBe6NAj7NSS+Q5Se65s7orI/XVDWprHwYv6RvhFRRH35mqsDA
J37DyYEpUEmZaXq2dDCzKemjs1S/LwUoe2qP2KWOWxzHyOS3MSehuWJ5JDmL2tgC
3M4c7k0Hz3InNEpfSf6hndnwoN/FxSYlVZToFyGGstH7IXjHw4eavXvkuCO5AkXC
BCbWaXGtiZ8z7Z8esaVGztWBhNBgUikltOrh2ivWKQIvAaPnivMBtcDJEaZuEzQW
CdpuTVItrTSrb3ho/5WSZ6RFkM8nGi2xAEAoRVVzBKXbEmvEypzK4UlPjNDE9dLy
lhGIP+j33/znvYK8S6oBO+ZKv1jLQhPImrT7aWmJ1NYbvyebiTtpvNQ0IY3GZIrq
VcZirv+FEHHgQdiWjiYvApxO4MopyHpUHUjeidyiiFIV/CL8y8zY3hXYCYyO9jO5
YDoO4yyOG7r08DBHYc7io5H9/UGkMWZFgw3Bw07mpQkfx+ISp9nmptQgDr5HobLg
gI5SZp2gXib+Vr6h0cDsuXVeqpcHfY0jKfjX3BmqKbRruRAdfV71IU0mVvgQoNwv
P1mwjIFz0hIV3ZjlGLAzCcdyO7aDQftCIQUMeOUBTNghLT2nbb9+xG3zS5EA9+rW
KqPVbMaDjYffM+sp8KhDo/+hGbJtUF+l6ihUNq5wURpY9EZB8Br1YShJXm9I05G/
FsLqNSnO+5ZpCbaDIGg7onqv1FCBaKeBDr1MgNej9nlWLbtP3XB43yeWIhRgfjo9
20Tg5dlX2WLS+XZTibGt04swZCOJwCwr//Q4cWaEnK3BjfSaY90RDS76JCWUbBrK
Vr4imnnbJrwvjiyVa/5N80/d01SyeaaNft6J+iNcFTQe6FcA9bzdBpyXyc+Q3eFR
vv+PiWgg0hPXuE5EHasMRHW51F4Iq6Jt3bqYNW6FaSylsBT3pjpPanxblDyPy/vm
wG/e54cXrRDFTpzMXEhFo0SFZKgj1juEQHdxrMDB4KmyEuDglygxxVlkfjno5ciE
+NAoxBzuVfTXLckwJZvX0nAxpIuQBctAaaaynfkkEFrA9Ac8SBySGJko0g3pEUmB
Mwj82S2UT/ZR34sknpJ/mA4rNYKaDm10W6FCUE3PhDd9JqewDiZd7V5MM39bCjeD
byCviHnbmEKPGVkw5K5hsblPUO3/F3O2trlooer9h/p3vfjDUvBvw5+Xv01altWt
9L5M8fHG2I0mFb34UgJwNQ8tn8uDNdC4omDbWIDXeWhG8aMUF+NERZhLMM5A2qz7
VUf0ptayGdpr3oMlCpH5G09dlUQFkaLqHW2Zv3a6PKgxuonj8glV6JVSNf2yBnHM
whb8Skojcb1g+SFbx3l+aNsyMb8QhCUm6MIq80+N+bwUqdklOl9tDxo/lzlanLn2
j3zPQewOHJnh5K3Xqlg8087zp+/Dt18WhzP+SZXf9Bjq4ectuPdslsQXXG9kgH2r
cI3eRh/5mzS7yOl9BlksWmrnTiOrfJh0gJKbjAN8AmT0DWG6nYXXMx8OrwmI29Jr
I3iepFLHCPflPCkQYPHLWzpbY4TslH3mazU+jR7KsvH0l612+qsRj0A3KTerqnUo
KtPIjM+0T6dK1jjA6IvagtXUhcaaiZRljpkc5oynBYCUHUdOodI4/kZmdjSnsjam
abQnEH5cHqWKElzjPoVTCq3Sh6aSr6kxHyMnhjXgsH8oP/o4Lq6w/QZ8oT23duZs
MOW4XUzukbHIy7mA/iBmrsH8/2cvl18u6nzns5w1UCoViEYNxIN+YL1KeqvIWjrn
xb/CQ4kbTU9bSUw6DKhf5UGqIIqfuZ05G7P1k9m1elOcvPIfhe02BPTsYERfBg0i
+AvBIkFEMBJeRFnrp39lxoJe1XY6fD/ng/e8qFON8PQLx1sQJJ3fIbhTZ9JC7Umv
WozY2wapdaqbI0VVVIPLC0EZvZImAqHd2bjyqtBYyuB7sAZppJNqGoerAqJFl2UD
Lcqcd9pZhQnpcS9itG0E0Lc+kxibQag7QH57NHXJn/Bw4QpMwQmC6QH0WzF5VjMZ
MQYGHrtBWWl+ha1Zo0A4GV09cIqm5CNwVA6gCtjLGukkHlAfokXUeXbASvBO/iLB
LLtAuXR4KiELNWzQaO3DLuf8bUW4l0hECedSWaP5rhUiSp64LLH5c1E7xFURv0zh
mcClF3SQzyY+U/vYwQ0jRUsIKWCJUCuXKWh7vprIjZb6qUyq5Pij/0ShEFJaD7J4
VXMWTmYQSx8vG2N5yxuCBK/CKQpU98307zr1xPuyUA4zws0IcIQpXryd+b9VGCTE
xkNfZIlw0TGYr4kjVCyPsFta5lClb+FPzEsInln8vR7E3uk5AJX1Kzdd1DBKogLA
J/j/lJWmpaCfaDRs/siOdpk37GCosj2KZRIPCbQdBPP8qU8Shmh7o9TTlG07hUt9
20FdxJBBv1KWZiq7HG++Sa7xaVpyHmNPhID1oddoEAT+adkomzQoRMNI5rbANA56
Izq7gRmpZQcuMsDOfXGSfM5Q9wvf0YvIoXgCxiMIEvHMv2YdDdu2DqdeCglZCX/p
4c6zxDEfuzqVY0Tfvi+vKeXCJAvy307gvHkE31Q66p6/9VJ/PVEOezT+0C7EXZ80
Ntq51VZ5mkcoI44pU3KXumDwMdIpVLSD9lNZhfiSwj//ESyCyH7UomfNOKqq5j6b
gGHXFiilQ3wxxiWMYYajbtcE6nmkd6kJCAxsJ0QQAyeNknsYNCGX+R5GGYzRhgzW
5ms3YAxyaM6EZoQzKu74EPxURcBErToYhIQa8gqfp4mbD5Ud/p7Wb4rCKyP/rMQw
vt70/Z0pZnoH3f9PYa0dXFTRXW8oEpqYSW5tuR6qHLicIZv6jgC3NixW+UIS9aIQ
/LR4BvKuLr+PIxYKwMDKDA1JQ419/C4vUjHSzNbQ3ReZoh1hshC077reXXcsukY3
OrdAte8e/sTIqs70eJWcaCoK83c2siBTmpHFNBBvWREaRTN7QeyNTDdbb7kGFy0Q
Lxeq6/ecvZ5VDCV9vjhuzH4A28UEaxVwlxiJe5emM7RneLbYTz3vmr86K9L2GhKQ
vYrQhVjUzhqlEsc5m0pPr6CmzAB2BfqGgu6eiWKUXmtTO+tHba/OyXUlv1Qxlq5w
3DtwsE2mGU/QAT7e1rFlzTy1V9Vf6uKVk1z/BuBYxYJhv7uz0gLLLylNjvSbr3Sx
uU7qSLYybL8NrM6y4uT5SAgUTcosItXh2PqH1Zuz5EH+Vn/0dN3WHWkIjtiZ0+vD
+VaFMHYdkjVUYot8uFA8UscsckQB6RGg2eBpx3VHhs/n8Gy0VzRmGoe4B1qEXb1Y
/xPtuqPP8sDKZZmPpfH/408pMDCBT5B8NSJ8pypulHtIhZJ0tOjoGul7THeTCpnf
SWpFWI+gzC/NjoZErx8Msu2Qn91fRTTeog2V9JPRuET2Ppdx6TE1vTPoET1wzBC5
XbPrIkk/Q2iKlc5QMaTS7ITTatVx8UyI9aUg174W9xOuQD+c2Z4smTcAzEf2hh2U
CNKypWDKGDGfyKOcCkM97fSqbDZ0JxVMMnGHP43N6oUtjzJBVpn8okYr8xjGYDDg
fFfjSepfa3sLWlmY8MML+UhqO2H9+SisEUaYAOIIKPf66cY3+xFFOGJtdBjVgFQB
m6JoJ3XLsj3+4tax+qVQWs7nHnQaMIm5Oxz2k2macMIsX62G1PTanZs3z4e8uHLH
6pjKUIfiRYZ9Acm9bMLu41RRyHiWht0jaErfS4pMRIXLO0fuLMNh5e4XcrvLJQcU
yyKV//kKmvjJ0lQ87ud3gLTM0v8jkCEdskr+BC05t5P+PSK92PmVzKNDdnqxC8U9
rf3l3TLufWQQNicmeDBEMBCaZcF1GFok+POVcMtx5rk9YlEiXWADWq29nM5X7rBO
SExXsMz37REL7I9vyr3teyKQHbE9D6bxJ3q1PWKkFiu09coeimVSG379eXVkmZWk
DvcocjLSnvtyPDNmQmYOVqyn+kQG9Wpbx7kRKyqM8zuMlPJ1Q+uGQzzv8pGIVkiG
YlXfanjrXzYH8Zv/56JSmswzEGDakTLildEULR9jSRXYOyTNIi6BZLJKe7Ef6ELa
UaBqlPcDDPFgzcBtHT5QTdQ8FOii97GtsDx6SOZjFlbMYKuKoScQ57zzwbna8aWL
VFTVw0Q/M98LoJ6GLC36Mm9oDgbF+gCnr0sPAywCuMFq1Sne5X7EFCI4cPaZLZV2
V9OtAG9eeyRH0JtWEbIAEywwpdR9xSw7/dHoJWQ04dv6UsrARxjXkUuMOxn0nyno
3SkRIEOUBcTWXJ4TO+w1xS2NzZ+Bv18F6ELl35itfMfrwx6aLAoXEHxL7l/DBPwR
6/hWzo4snYt6F2/Buwl6IinchK3Fgym1RXrDDxO4cHBeNe8mqnQUVmP+izLUTShe
HPQWt/ZBcy+NZBYO+GcyJltfrr8icGmCsBDFvwqvw1U6vCCJoCedKxhDXUZLHcbk
mIiHhgHlCY8DrW7c3r/GrlakS6E6wdlgTlsmALKxquPHwJ+rYgIt0c/vVjKHP8t2
KrrWHWxnwNsPv0GioAr/2Lq3saigZJVmFPvP4I280CLkK57k2jwYF1wqtdXkzzgs
3OqQj1HxAfZJEVL+UnyUAYmCKP+vP6Z3KIC6nDgCtrqMTNi9oqZCl0dtSyofID4Y
8C+TFPg/vdaSi/uj0hBTW3pXIBBfq8xpH1NJIxusajmssW3VqK2y7IEP5xt+xHGJ
vDxTbsQ5qPcQQjYcFIlr6g9FevY/5yrtR8t91v35M8oc+RBVG7TRbdPaIfwUI5sF
tdCzUs4aXkSf5D9tYPlOXLm+KeYUYd5aPsj4+iP/1otphSa6yocGpaqOxgvJZsCq
ChdJao8gEoOStLxj7DJeLCzbPjAp57Nq/cEyQdqipCVlfWGPqeU2Gl+nRde5gy7i
CkEiAN9D1jitl9kqvR7sX3f+xmEnIbLLoZZj/+rtM/lV48Xhpb9o/8oPp1pR2Xua
0rBerkzhad1EGVdSeMnk8Rn3XX60bR+U24iZqVQeV/lfXk+xZuPe4czZmqhfi55p
pnIxDemywVMot963ws3bOsrh3kJr6lTaCFUfHdeh55bX2ZWodBNPkevw3g6v+hBy
Fc2DWFFt4Qlxejzhnn4kX3Us5LxQn9lcUVMSN2/vv64BFt+ClO2lcP45mUjBvSpF
rrPqwo+aaUh7ZbBIoOgxWrxp3osxrWWoKZq2huna5MT6ivFvs0Q1lkTOEgXwhCfv
+Fea+o8kq4Jhgi7xxPl8z5ZYfZkzKIAqDzrxyjl/IR7V2G9ZXEpMuNwePjosBGOe
Dv1LqFqkY5al/ssJOVtV3J+jtVOiCTHg16GwjeJ4DOjL2aaPUh27LXr4mNqxa0+d
UJvYb350RP/rmyUFdiOnDQv5k/+UItPIjK0SCkljieMQ8eg5BkfG9tP71ZKVzoEY
lXkGvLrvkaYytoWpBbMtoAnckYa9Cld9mX5HZtcD5C3d+/aDEeegYPkirx3MKxTQ
QP+nMDjZ5/EWhIop6cQInrQJJ/vW5IPLwF7ZKIymFtZZesgldIktj0ecQ90d7kDf
IMpTMAcSOt9/zaKWvO98V2/Xv1ZNPufytUMktEb+YO8bBjofEKVmayskvI8FGUO7
tn3n6ragBrjVeUHWbQfoIdiwct+yFSi7fvMGMFlkWVlRuAFI/vpqE96AwYMjtSQm
+11IG1NfxCxaZcGetABehgB/NoWVJalNHwk+JP08y/GMVrzzTxQ1jHT9vgxKaAnt
5WV4y2nu2Pcb3QrEByIY18VIiop0z87sGsTCTtwE8nBMIsbsgbZVC+QzfN057TAG
WSGTsU79Px5zMwiyx5wotuUGojyAExALhTUdmTWkVaU0/YCg0kJ4O1MjdzI1Yb2k
G4L3E/enH644JTyPZeym7xxAcxSBs/foV+SoRLuFGbpt4giFZQGbLO4F+Hgi4LND
XwqT+sfdxf4ev6s15QhZPWuzbcJfnNC8xvBVBdO9Z7qhaKvC1Ve+B7wMvxFSwMGD
0LWRlAtaKjazraS99cgh6o6nka7QQO5JOb2vS1ctoy2noTSd82cEhjuPzGc+ty8P
JpzQWUzRBtnrX/Oy+QBVpyHHWyF5XOeq/JtxDi1kOAI9fsN0DC6Epif41i6CsD9c
kpklcg0we9tFQf5aLnsB3aXqA0iX3T4tqNWbJvUKJ/yKx0B9pGPowU7wY5Zognnk
7dX2gK/jbxLOpQsyRZ4MjTvRRiPpSotbES+tPPO9Jdzd5dSau5F9FCar451C/suk
tQJi64F9Cco+Lj7rHLbiqM3wqAjVPsvjI59PS1yMCCCtx6fxA39RkKL9tL7PuJeX
+2xnfGU78eZrVeJzabr2tfHHnIUBGxguXc+PuXaYDZlovl6f11wMrkJHAZEgQD9c
DhgabBJWrMs5XMtSQwVOUbUEVyH4ad5hM1yPHqR35gamI3o5hz5uS7YrQ1f27Ik/
2tpLumfGG+iMS3lEYjtQQ2tH+TlbpxeEVR66C6AAjjg9hI5my23jEolnl2WbI+Uj
AJgFztYzLTPSBXPhjLEGDOpp0CFHspzxGH4jUuovNqXyEfkIEZW+8zpgYTTBgfjb
9jPKtRoCWbX0rN6GiXxx40fPTe9linc0gfzcSJNzk4e0eHprlBcw8yWQIdhHd8lu
JQTQapVUenxDykLYYH5VbdZiAvXUnVp2mOMJy7ZW2WbCeUXS4bdKdiGZwE47Igqh
7yXuGmdiAy/UmwEod5PcYwMXfP2qo3X0IkaQjVZ7/lv1E4Qs64x34RRSiOhw6Qkr
d/ihGsn4z2k+m0n9qQr3c2XAz8VXanTTXrBaDU+0V7pcQSQNAjEpPjfglgHzUvuq
27WMD109aw31goxqlgxJcwtcu64wDq8LMeJ05DeMEr+5ZphRQ9295tCJOdpZwA3+
Mz8lS3+migL/udPeq3prunNpm7fW52bUzeRSdxaOG62dvBdLrm8dfm2FQYQTk2Mp
nqWvYl7fo+fDadt0cNrw6RYPSOrri0HAKbIdb5/U9NdpuAmr/WTcRY+nsdwnr0PU
ZlvJ9aLQrvQs14S80nxaXKmABEojW597W5Rn1e592OfbI9FQgIxmjRMGqa1hQr/o
wh7DgyuoQvZEJpQEs2AD49pQDPwNQyMrJXNw0n0kIoyftoxq0pBYvGy2M1CZBL3O
9MsLJsXvnPY7KAMqYb2LHMVgOniWmmfwht3JAKtjkjVAZf65aieS8WMJwKYgIrqj
zi44Yh2RixRpU6jhVcvXDrvOhlkRcnyCr6xvWrGW8o7ezKCFVlsCi7rorP8h7w90
JW/cFqTXT5JVWsrxNy5FsNpEaTk8bkgP9b1zKnDloSJ2mTfeJ+b8sybviW7TKKMi
PDjIYRFLmGaCRt/uzXGS0h8k93DzTsQkJxYXyEIyN4h/8obUvrhfDVOhPNNNdYTu
x6iNLMPGDhhgwDdH6XQAJ7wzartys3D1tik266aNijayWhC6aBc53vYS36ZvYAII
f5/Vo9EJH1bc0WMmVXvM5xAXB6DUZbD6MbiKrS7FEQ96+9o5hYhaHlgvJ6UTPTvq
FJaJ7ONwWoyhVFk3r2hHFLTaKWe7sGjPtcyxy9gkyxpfLil8Q8ZIrfr3JhAsXPXz
Bd/OK2ZhiTHjwpC+kYQpSx7A9YXLI9C3wSI9W0A0iclNyRt4uj8/YmkaWNT9WHNt
gb74X6UNwZ+PAkkf1leQWIcFotSetPnzUXNI04rMBvrF/GOkJyZwFnLiIbT4M23n
cqrjzJ/vJawb1g79eQclPhFffI8N2QR8Rt6fefcbjTqP/pz3fykaXf8iY8/gxhz3
u/E5NW9TIUdvbyveCcT1bXFLHaFhQ6OF2D5/3dGeb2bbftSvVaaF9Z0x0xL/aqD+
blQsSh3GknNBMKyv7qmRV2pSNuX5emS4QboAwRbrU4yPfDlJQAqespoZ/2yJ5IYb
gjcju4D0vGIzyy0RqQpW6VrW1OaGjAykvZAhckDysL+mJwCESyJRcn36FOJ9zony
/5auuCsGQaHMDCXkWJDWXQ8ZTHJBqzDML32atkI3Rm0hqLdZYdP6BaW3zh06Vd97
Tjek/HVm/edPCgceGh8n+VBmurBfNxXFznSr2RcJxnG47wz/dJUU99d4hFmYdhAs
hXojdOd7LPcbqkC6SWoNSMi9QnyA+pnvZHm+960HzM+KsQaq5SIp0Q1+/jmB0FpH
FPOycJARzLDxJf9yD39DSEZ/SsCjOxUbY9i82bUmXguc0AeE0GnDG/0YOHmUGJkL
IBZWaa6zRd5IQU3CJyt4MiYXjaVoM+AMJuTiHfdnMVfizakjn5ggcOaXSE/8ocpS
GTtR3nmOU4wOwz3yiIQD6YFmZW3V0nI/gaBxHX9ZWOh9+ps/jVv96gRpl6GzwQHp
VgqM9nt6w8mtDbvoQUspauL0FjsMfUfMEmkwOaro+daV+AmFiUot/7SfMFrEXNiE
+2BLtnxCUL6NYOvxuXF/IYM1YSHOPw+B50JNCj63BNQpNW+71cZ0Q3OgGwimTrmW
wFaMhIcAMgY/w//gs0YtktQBqeElT/NdYI9IXv3JYEWWrIuBynGZ/f15WB6HAhOX
N3Fso78S0mGORPQxN13ruaVy7l1o7VQ1nSwj8kYR+tWvOSKDXJM7hvgnOBeP1NGg
pMi54z9kHJFPmt09LpeiGQ20TDN5IlXTBYREKKROG9BFbMin5g3iTkqffhIocsU8
reYJFV6lJ91Or+94GE3zcN1QOdhV3LOS0a0R8dlDLiT07WaPpyoGQlq7O2RK2XGE
Yn+5mjcgDUxC0Mic/8DCJw9BcCgx03bhgD9hlrMAD/4tCJrfIys7Bax5s8y9Qrff
Z0oPJHpxWUl9LAjxlYyz0czoAguV9WD+zaw/KqkE3pV2w2VMQ0WpJ4veYkF9sXMr
36hd+lmlVIdC8xRDtD6XX6MgGPccgxiwWcnDGbaKFdMxhbkn7rsd1H2N5D7lb3sY
vfJFDyB5BtCiXgTXnSeezAbax88hCFZR65ZPSBmemAlbehuNQrxDHFM9Vs59GxDj
XNXquO206qBe2D8iMyh7b5VmJYVL5n4VXpIhaPswJw6UJJSSXCDHRWOBhTMlJ5eJ
+SKVWhavQCpxe4d1bTXzWSAADOBEF9ShRx/+gURD+wljAYsLWIzDgR54ItKToqwP
yNi+qw5HV13veFC3dVvn5Q6CY1sBr/7Hzqic9UtZfqUuJMWrtiwPyTKqqdPZ+ZKn
BSMQGNnPZTuqyEjywS1XmxiOzmqzAqilo+NSAhpsP9+Tb+e5BO+hqjFV+0+BiaIX
xmA1mi7hOv/9GOnG2jzs/wA27a6bufcRQeeeyxX2Fu6r+BI9o3NIv2X1SP3yZmD4
Cnp7m8ifaP9ZWKF2Dnf5J386ju214vmbw1XeKmysG6Kgi5AfIGZt6MV7SNM9tRhZ
Taf6B0TM3vLr0PTZwvq4XBSCSdNvWybor1UFjZsGuzLB6WmuVxyIf0/CT9nQedt5
uUlokRRuD6l6UF9VEIB0efgHn1EhZrnt3F/dpKEvD2j1eiw3/c0xzXdcitjPpUps
ALrIjQZEbWtiZ16l/xkO+BddmaU4D2dLN9PQkXkoJR4Xy49HPr9NMoUpWkWziykG
79D8ijklKGeCd2Icgr+oCc0LKmjJb4FOL0t/llWjI2F6yC/TEQf/CVaYafpz5nZh
rhvwMFScDSh2z7qUYV+8VYUkCFhYkaop1S8RqXL1JtfGxWH6la1G1eKB7k8AjwLq
CPIGETZrq0V6SHlkfbA6of2xXwWOpvPtgXVoyxvRgMQWOm1FctqXbeXPi52I/6xW
H6wQ4vMP8/008J+TMEQ/9EqCttSMF80MQ9fVHA37A685otj07Vc6xXcMDDUiGwGq
hG+82em/JQEPOWy8tEOjtsvHT4UjNuCjZpi0YL4wevJXbkDDI9mdj2aQ6UMUCea1
yuAMuMOXqAVM/MpNHAXeulyfF8MJMgj+Zit6kHFHTvR9zK/DEg0N8oi5UbV/L2RD
q3vAuFBXCbxL9Mt/xcSN16U8PSF0Bx2a0Od3up5KFE37QGtDPsuEj7MwudShry53
NW/RxSvYYNXohCni9YPGchFeuwYx1q/hq6fKT7654Ykfd2iCQF7Ka746yRTcGL5a
VS2F17hKXgCIu6jgDxr2tH1oP5J18D1fc9LtVmyRvYFUvABJJv2DV6OTz6ZY722U
MP4AFdcGY83f12DmlMtVmt67FEornaIZkK3iQT7KOc1qkCX0TGNvVrVXugnPQMMd
LQqTvbSscDiLwjmblvDhQdWuALU1JrQV6jrbdpPKkVfRMceW9ahAloVk65DOMrP1
iNE9If/xfPMBA9L+F2D51h64DyQI+DVnlg+KzgHWp+NNRVvWtCAv8iUn7StwRGz9
HdiwpW1hmH5Gfsn7Mg/BAWG0FtbgY8jDPb51Kpr0cvnHVVIL+KYDtb2AL2FF/xbo
H3xrjMuCwDPpFWMb5sgt/dnDHmQcj4x9C4w6PHblUQeffq3/gsPT4AsGz8q9vKuM
jCLZZXxavYZGW9zd+0bDqJuP8MuW7diQu/J0+iDxDb195hJg4Fej7Z6v9SD+vxyI
hMxeQEZzU+F57z16x65O0PkbdCFEWsXVCazubIv9HX+3EHultCUeKi4YSRzFV8ch
zzxNfPrWo7gSypoPtyeeMkg0v8HLk/2WPodpO/emcbVlfI0F4Ps9qiQMpE3zEdDn
8jFGk2Dhc94KdUvhQumLSROUIXmvsXSBLMm2PqP0gSfF+34vEEEzRlpPGe64OoAW
kma8I/ZA5yTt92GSabrzSth21sDMl1QBSqaIViNUQ8KExhuBaBZmoWXLuLYqV+Eg
Unepge99emgaTUhzu2pC4OonAiZvscPkk9iifI34ACd2kt/KBaGNpRe1dcfG5tLv
S6AlZsv8ipkb3/CWiC7TQEd3a63gAybYMD3QFa48ppBphO7RwyCjfmT36cCUQFfE
KAnq2VpYKT04BuA2Blyrk5tseM98Ae1TzuDyPh6wapRIl6RyGgZX9F2ODxJAlKwD
8Sj0M0Q3MXUblesxvyL+veXaEbKFJXtaxerjJPjlvU/gY22WhnL2ieZTocE4Fpco
k0XM7/xtlRgLgQiXx6l5lVhAEQugya7YUypJxbY7GJsfL4xWnfN6nYoxwYxHeIe8
zjMJgvFuhXzKClhc3O+1H80Qw4ekvTr2CyT4YHMCFPsml8xIBDDhVz4jcv2J2cMl
gp5AkU9vf7LCPTViyv9wxVzbC/DAWsj7FhFS9jKqoXtFXeBZCrJdFA7unq7IJHwZ
17Uaga/k4WGyEMe/1kguhfuU8cl0pzlRs8jcoJRe8LaB6jrc364rJ/N109jbq+8q
K2/dJICqUFhOe2DvS2yCZxnYxYgMGIhx4icvZwa6Ulfjipks1WThcK3/B7cLswB+
QaiIuCcw0WVFTNeg/I/IVs+H3DkK63jqd932Ld3y9QhzFvL/3bTbo+VCQnkO0Z8g
kJz7jJfuqgZCMLe+ujofdhHWhFg1n37D82AOyWiqXE0ln5zL/RfIvnbojwRd8ziD
a4n3iKRgjhhHC4wkpPWXBpck2+OzAST4KIrYXVS4caO3m0ZnZaO+QNS1+3lXsS3r
o7l2gS2C4UsthO1InuLWydWhzaxgCcPmueBPhEVDm+c/iWr9vvKDYq29d7m19FWV
suBCVN0+qXAN1GE3fR6r52kTCHj9nyCqKGSzZRUAc52q8O1f/x4nZdTUkbLfrU7A
WeW3MfOO08fW731Xm/xNkkA4iiEnd1dgbSTZq9dTMryLLS0/PiDXUXKZvQqB/YTs
GcABWMFwOABTenUlcma2bQ0pnXTHSx7m/09Btf2iPFe61w52TPYNTqbNKNoWcPNH
1/13/104JlkERnsQS4wu3NELecz0nhwvLW8Co23r6CgmcD3YQGqwZq+MfihUKoCW
a5WvuzDrlc48mG88rjvO6rOq2JfVXHDffgjpBx9lr4dS7iHWq/D0Si60mHpf4ZUO
CAkPOaj/p0/1qXe1mnKgU3uRPZgR6+TaWd6fBdQG2vD9dzO6YqinEVPWAIKIoEyB
IkkS0kYIZCKUdfA5PFUK5VfhfCSIFUKNVCDJZxqbq96E1BKenp0Q9WU84cMSmMTk
fp17L7JbEBh1qTmRdmMSFjiJHLONoRy8Nmqsd3XAWw5YJUgW04jiOteBWzf6R2wL
B7A812pTtc7uQYZsFMagqpx5hyoeU3xdXG0/wZMEJIJPg9+TADW8AmUhk6JF27Jc
frunu+uJflcjl+uPNHm10MiHLXVT3S6xFuv4eR0AKGVglYyWbj4JFA47M+MR1wmj
HJeUXk5XVdS9EtVtURii73IO7o+U/95e6Or+Vd5ICSvvRxXmttmbkgvG9SYDoEEb
nuDEp7bz25fOgKdus4uTRfsN07zEk2Dncg9n8snZRi1gAJMDz/Gll5vdzB7GOmvA
L/c+hGD2Ja6H1aaCLV1r6yH03OoeXU3e1r+qGOw7N0kYQzVYiQxwttquJAIAK6nX
Sr9bsNOXJ+mtpQkkmLpisipHUiOHHRVSUInIBk58iHJEXvb1VpDENR8+VtvOobfM
C/PhSaoFfPc0QP9yXscSBZJX6mUYMgn/IzrXBmrvt5PsZD7Uvms0/BV97wl2ozek
Hln7JHSfVBIGh1y/F6+snITVpXp7G1uiWi0Id2sV8KZS1wihlR2KNAIs7+wBzQrO
fsoxjpAJadUyseV/aCM948y/ePBgA6GUVVgaXL97fTPCvVKuM/U6J3pettrgDbSW
RI0tz8uKEDI4qWdWSB8ORBcytYVe+Y15PzrtvnYkHeR+B5+Ol+lU53YaT8NE5h+x
uY/u6XdFurtCmniKuWlf3lZnGa88hOKNg82UvKD0fU9rGHXw62BuVQNAmCxjOpkz
XxL4hWfEkGreOUSOCwJLLfBBxgiiVhvjOlgID/cbYUFHfrwUKm4QuckHuleHXmSk
LLC80SKngk1Oc4KcfPVrTUhIKrjxqEjfpaq86NH4PyNgvEcGqM8/Uq4R7rVneV4S
Y32cBFPfB/qkiQtkTo1dLtblhocJ7idJl54K22tkFSS8yaQMm3xpbWmd1V5q5OiY
Oq3vBJq6OHshPFK6lPb/bMzAYG1m+bZT6a5wHz7MQ/bSUmb5zplbccUyZ01mevPy
U7/mfwU/3pU2W4TnJhwxzmL+Hgnr3c4fPkoWz+UmFjBFVXjPgui1v3fbb9nI1vYD
WG5SU1WkUSWjyhgGcWCYC0KgqnTCI20yj8FvFBQoooO2/HE6Hw2ow49vTV+CojGJ
sALZv9w0Tjz/HvnANs6dUmyqaBTPO6M7wtcJwFK2W2ZK26DP1VtZ+itOAPSoK8M0
5xfAfDmO6arF9LZ304kDfEIsmdbZ0Ye0ktyndRBf98Y4Tf58Q0QLGSsQvhz39api
2GU22w900fpoUzp6/0Hu4XR/0GHP7yET+HIdDGKm/qh4Va04oL9NhW600aCb9Smm
GMh1nyR/H/Qpb9mUwrYbIotCMOyioq1r3v89jVaJ2KPnPIpyNQIhdLmWXoiUVuyF
6fAMvnEQwh620BoXgz21hTiZREi4+JDgE8R3c4qYNiMQQ3DJPcGWQnrfta1JfJxa
jUGL7tVB/tN/8o1RQrAxWerVAwg8cmYJOOIuyVvN25yf2Po/rdjGIeShWs5zQ6oD
fg0KPwtbJqQCE0Q+tN4RZnzQ1CPwk/LX+zllxkuEPm/AH7DC7igj251sPl+a5iM9
C1jggVctu/JpYAzrQBWqfFp63WwdfxghN172P7zCmtEBmKrK7NnB0XiEDBcR+ZjG
QjQma5ukc8HSJKIp28LD+OCjsu4cELwmM6fDCF73//VHmMTMyfNmWd/Ni9jkNaJH
7iUDJ9q/ctYGs08ePnCttZCCxs5B+ogEFZP6TSMfd6E2eWKipJh7EEM/lTH0mY2x
gLUYeVHJ21TgQkYAXHNAFj9dBw099gyBU+QY/bRAe8+mbOMT41bSUAjZJyETdjp/
9vqDLxRKWEDZ/U+LEWM6/plyFMMvycRv13JJBNlPp2X0Gjwsq+XU6MJ3YGmtpunE
CXzhxDJ3hYRwr81VuNtthTTMUs62bYliruxyGOySQSUq/A9Tq2cn01nsV7siO9oJ
cueYiHdHi8GBsmqGCgmo9kqjbe0kCMeibf962CHOK655LAuoyXaWG0p/rBFiIstF
/XUzBax5D5y6p0acpnfSuVYev3NpjQtlrShVXhArjZnh0MD4558iUoEuAg2r0pX3
legX5GKU/HiLsSxzoHTwVygW/uMMN5ViQrEZB5pm3cSEyVieZEHB45D5FZnYVN4S
Xibo7muWC3maGE27EGysoTPjjFkkjc1caksOLf9nB5yQPfbsUOLqsDEbMBZg3T5W
/0DqeOUPhjxLpYEXynofWWluISgvU7upLgmWyL/r6+ST8yk8a/KFZ8JqkIAE5iG1
yDH2B8TBOcPEXSY9z3uZ33Gl1qZFyWh2BHB8PiahG1hXnX8eNMOTh06WEe+XIeWD
XPooLmRY1hhKsEY915yofGF0hWqi4UVxftCRgVgCdXEMK8/okoJ/iL2C24XO2lCS
eXaQKEWkffeOzMXvUMQpURkkvP+Zf/m9qNYf3434qpcmVPUAulfgcLOCz2cZWMC5
PetWaEDVcBrVvWCyrxquGCsgKShYsAp54b9vgAetGK9fnYZt6EYICC+W4f0KZI+h
zlrJZsvk9Z+KTYRdyrQ162XUq/L0WAqSBLPo3X4KJn7/vsUi7Kt+QeYxU2uL/MR6
jyu3Pry9+9Y7Iv1quMQw58ZKnwLJ5KA0DM3Z7uvdskZ+6rle3sJEg9ZNhtQz4JeJ
F5qCjjB4Fd7L+AjhDSWudVy9Nl+vH1+gNfYQT+nc6Sb6KHyr5PT/RWxDpCbgJ667
zDjxjfZFE/3c7Onx/MUsEiOyItPhu+ZFdzGrfkAk3XnGgxL8YwnIEwYRjUDpuJN8
XTANaaDuZb9wGWqFkL59hD15naX/GyNSiNl0B+oMrty+5yI3dULNHxbFE4nVsDu7
jj1F1G7r1520P9yhAmKYShoC7joloIBRXtteHpfekeVtXre82HlzbFQ4hdxBilFG
UKlZRHJwERkCpvBa8XSpsEJ6ufS2tA30jcgGPzSiuYLJMry2Nb7ZZPTNaeS3ueE3
0t1H6y5nY2/s1Oq0sZYiKl2gvhs2VLiL6tZ4QY4q46oAPgnxDmJrsxpsN6GOKySJ
SYp7SGE/FSzY9Ceof36lPeeIuG9JRcHkkSvkxCsbgUKFvqgHWj4CDQQSchtD5lIn
M8wdulRwmhZ3EnGr9dRwgpR7SV3gGlFZGVXjH5yJpAfDj8E1lsV30oDJdnnsVn9x
VW7OY6E9fGQZpeQh9T5QvS/Mcdv9W5NqXHAEg4BvAu+hJDmZMqTS5WMS0wSMA7VL
HDB02fDkC/7fXDt3fOu+8v/AROKh/uCpJ93ZFqsTNDVzIwj+hESGix7xpik/zizf
ZyXn/bgOE6F2T7SjAz4RolGLQ/Q5fPM5W2NuwwY/s50r4ETNcTbBc7DFSjR3ACGm
wdszNTX/NaX6mM3adWDrS5zWffSy5lnhew6QvHcaR9IxcRAljjRE22zHRITpPkJG
3yU2uawxbihiTf3pSRNXUdWJnEyk/gW0q9f08cgroV/F/iZtXc2UA6+J9k2PFwP2
+m5T3F1Wukj1vG8V2ri0M0JVYkA3B5wPrCI/m+lgSKjxetToWb1VnRt2SOym8jjx
UElwdpkb3Hk3+kynZsr71wkeCXkJuFIpenTx7Q2gjlDTPfmZZePUjqnz8b8lhQtG
U39tAk82IDtFe5dVCILlAOs/GQKCqEqNU0fC4fC5NcbfwMIsxWJVcXSbcbJ+WWOG
9xYX3i/omw3W7PRWd4USYXHp/xsQ5IuOQUewu/yj1rY8bdYb4bpXOtxfmY3onNnn
k/SLQK9WqdeixiLY9A9oU8R5k8qxyVaQgchhBFeNuojru6gl4URf1P1sVF8roJHo
w6TRiGnPMg/Cj0TxS0ds+Y2S6TV4jhATaupXwpXlRGJSifzy5dQ7skWYRJe5Zj3K
bgCCocmGZsfB10n+T/GJHqhPDwzgsOajJmHRihlbHftcOaWyhLhpbXnpULactJtV
xyTY+DxzRGvy9+wuP87cP/rxwQXZUTnd0fkMWJ4//8+tEsS6H55cS1XQ/QEwjgPl
qSCEvZ839XVtK3ySaS4tlJDFcQhF4BLFR2uVyIt6H7MZbaPVST4g9qT1AbF1NlJr
MdIqC9gb8nsJoCeTLhl6IpKhWbuaL56RLNDWjAXJf7vETLwbR8bXifxdCuh50uDn
aJ1WS3Bf/jyo4g3RtiieVvDGnnCRbrua+HQBxGjwwfhxd2Lgo5NDML3p9ZL4ZCjn
3M9SYK/N3RsWp400Wfu/b5iWD2k6u4/IV0DvJmFBKIDhrNTYFBLDQLg5DzBHkbgq
EcOPRhsZCDwYoDr2cf+Dzh818ePuop4+vNS1s2XO47vFpqNME7zQNrSKITuIYZIh
wz1/p8rshNOlcPkhZLSY6f5/aJiJQVPKJ7zMaB3YnuJfgRHxpqVAfEd/Gm00V11+
EUFtD4JMAUfzN4EVfayr2U7OPJ2n82hyt2laeGd8cZiv6Qz9OEkzyuyFG3VKPaRN
5UCYZw9gJjhhZFNLtIDjYVAreYU3UPtBp1mM2BS2I4VUHGw35fiUdRFtt4q9xGBO
BXZlRVhJvGrYfCu96AlSOMmqzPDfp3t55pyiqPLMx8OAszwbREhvmMPg2mAdkwny
SqUhIt8eigfHJD/9PFq/H0Bh26df9cYBNhMOuuCwwhnly5uX5oEjVQx8LJ6Sf1ND
osGXyfldyuTXlc6dBiOwy2CRn2mSTKfT3TW6VVaIlVyIoTVJxwjRG3vChTqFuEho
70ZGy3iJK1YXnQzBiL/b5GydNGttduslD6qOAxKN3ZwAtaJnLK/h0RylaojAbwNJ
qRS2dwl/3pFJqXQRRoMcl5Q2lgDn7ENx5lQlhcuKCb/AhTAof5tiybPERp2xQzqN
V3WPaGXovuxu5nsfyCgBjZI24tfP/yKouF6ofnXAVdlqGhy4/250zX0xIFj3LTy5
IdZEXl7dVdodHhAfo/XEWAvYBrjmzT+C7sfcuVGgcVPS1oYQ5BUafZY7+WV7lc3S
MQFktWEZzJYZwiFc0cw2cpvWFji9pAdMapNhvRyc9h2gmNiiPRnfUxa6kIJYpE3s
Wj4Rp8RSdDLzVtDG0kt0Ai4O9U6AS2sGNrfFQ/FdkzlS2b6d7/LahKqzSodjeZd8
fq/TcdO8sTOMh8DGCR9NPMNRpDtRFQUXvCgpTMWAPsVyQENvIYmPfg+MvYFi/D2T
2zb8TKu4prPucuohXAZpTGhwUpnHsZir/JzaoVgyvZ1eKgkRJzmzXNVfxYa3Lhqn
72K1CVUACjF0X+K/LQ9QqRrwuq2BxrRQeOLS7rOhVgHXQPQaSJd02A/7AJElHJFe
/xIBX84esFEwWKCiAQUl30FBFTc2sU7s9x+6oWyb6soVqyB3MSUo+0lHQnn/ZuzB
SA6n0ueClrHD/xPX2uGRucZTPnnCiQoq/dzoiKR+3DWhzL+bf4Ja09nDV1OFGibp
EWqxIxGIDmbhlTZYN4dViPjumRjCXZzAz+XJRNlPOn7EAiyDyLEEWpkZ9RzQtbSk
T715s/9EG+5pyyM0QcLjZeIQJDtQF/Ic5PQqfETuqxkqtidLdXuS362yvHMA0z+G
eVJ9emrysgUHm/WVRKBKH67K8HsEb7RSTZt0Y2tkQh1qpUc+128XNehB7j6KqoBY
QUnyqz17Zp++keCLTP12pJh8B96kSdsI0FDoEenipvIsbVKIc6ZnPyKVWacmIb+8
cP5IVHaE59+70k1hjqybbna8ihdxgkaiam2Re03jFB5i1UkrlWmvt0XFesels3Jz
XU0CgCw3VX2ld5hK0GAYpAeNP6JVpdWYLReR0P8dwikg8Huq7NgPTj3CBlF52aH3
1CdAHdmZ2scGRYKxPGA/Pkp+3zRS/UhS78ZkFgC58v0h7pK6KRqyD4hxppY/mN58
3rO4Xrvyz1HHSJo84LEC8E9ksSEqs6Tu0QvxgOo1t/ENXItXJHULm4MNx4HFdyYr
2D7Zm/iZ/5AxX0J6+wH1rFNmM3STJRg+0E7cugxT3ihujMppjFqyBsnf1GPSNmfN
+cVOoGiBxNmlnSuQXwpnSpg04i4e+rDTbo6Weu9FWHaK5Dq+itOshq3lxeKcFZ87
Gm4renTKc1IyazC7qEazsIzNBL+EWpJ207Rq7sDZHnSpj80334fZKtGe01hHjecY
PAotL6lB7AJlYBP9fnZdWnW2BHxOO7J4wI9b0c0BYTT9naKqo1V7sGd1xp5DQSvy
OKaUElNvG11r9OpsdiuylPGWoCM5iioig/Zua3DuuPykVcs3UpIj83jcO1wbBJ4z
CBwwubH6xD2thIev1UeWT1Ht/f+UnCChGpCheRE1CAv37bMhSE4KXYcid0OIQ2MD
Y4l1lYZj1YjrvhCK8LNvGOhxr21LtS/tTbpYn+6vEApIvA1CCyyMhP2FeZpmhmgX
tmPE6xfKFCF0ZDI3e8+8dBazKcmUciZFmtg9Dlsf6ai3l+JFVWFntHsd1fA5oAnQ
RuXI4ASgRExuhWxu7q6JYhENK10W//ToLwhpTaJmFNrWJMHqnUBJA8L+H79gVh8Y
x4komizYz+5htpLub9C9b79ld6pU3WqhLI91MW3i/2PlU9o/k7lQSWyo2eyLaMZ3
02yvIplTm+IuJeCFIEV0cxCCK0N9vpFvAAo+X4H5FAIfqCDpXKZ1ZpFh5Zy9uAQN
1/QosUf+CeYdWciVDwe7DDm2jL3aUgZTtdY/L5svDKvgBTcalSYqJSThb6FWWgXE
kY3XQnUmXuSE9pawuPOiKnTSCIvCZK4DfzLliBZlP05EVr4kAZmFtpdPA3LxkQeA
ejRV8gSPKCI+pfD9lbtChvGzMvEjJuNcn4WQlZLnXxAhKPTyaZ8dmgzV/qEWaLU0
Z9/8VN1P5z9sC6K/cY9LfJANHzuHd/e0iiYIz2aapkOaDKzYSWSMCnz0/q9bwrXZ
deyZN3uRG03YGc+GqPWNf6gUzzrxYNnmiYdSY+NzRTUhPQtPA94pqYbVElG4I6fq
yY0tXzcBTBJFmlz4hi4ftUG48B79QDyml9zSOZ5nWhrTKVhycwn339phbXsXJm5H
1hZrW6q9ywhoFWKpzVCFKEnHKbDIDKgvmj6yqfmL1xnVrHxvqzLFCrxEzHF22F3i
WK6Fu7YqzLMBehqGxdp2UEZloIj45m1ocVlgSHFjCmwfZcUgh8IvIRd9bne/Whoc
p0coTyTIYulhLJ2oCrgR4KqPAgeRnn+OA+lST9i5GbCww04s16Oo4d6D3redGOtM
TeeOyecOvWmgee7EUgvdZMkh+aW1awY1h0pdX9Ui9c3lyBih23ol7OGtWaFfv81w
OGi+6NspS6zZoSZHy9gaLlRBehNQpg9GLVyDGIT/mrOF/vu/B8GY75fZxQXjto1+
xiB79ExZdf6/EEBSZ32CpC34tf9wFm1KYMVHqQLZWY1NlURNom4SHcKd5SazM30F
WYxS9fAwUDoJan/UpOtyj8L4S+g49rZZ4ug2eJMzhAVlqdhRhQashG84PTMwWMsR
WX+727Zz/Ty7/7Gz9uWyPh60HPxamS4YkVlkSVlbRss5KjSJPL0rApqBj8GqKOQI
yxPfBXkbefeInLYUjJoCjpCk/eCUCh3QfWteh7Uf/PNbWXc5/Z+FAwzBJ7IPezW5
kyXeDtuhIlgX7Oquyd8RaiSpmstfRueklKJw50OIlcBkdelntXZ/ARQCJtYcp8+R
RGcClBX6ocm2QrGEsk9coaqDUO+OnLP9DoUUBVTNZLbeyjGVrwhAhQDl+cO5Tj7S
SoGIbuUbBsFOpWaD3L2LLkVsr2MttLK2IPXXZhEz0y8+ZL4QTaJtUy1baTuprvNl
jVklbo0UaM6dixpICcKmlT49lXuoAdLaH3APae1455pjpqSgCkCkbF8IWg65uWip
Qt2t9WYiEtuFSjrVrStqiORGBQE3Pp6xmwOp6lp0UvvXyD1klNk2seJez/aXEfaB
FILFe8XzbwfQ7SvmLRM3oa59BT9pa5ufg9hY1OloEz7C6jHhauhEHv3XB4U6em9O
Uods12ekhUZ+ysW9YCRAKcgqD+wF9RqGZ/7fPzfWY+cSqN8Ymiw6DGm7IBmzOzAq
j3ZgIjjhyRyxgN49jxfLp0kT49AGIC8Jy9TTjgpSil4eOXWxq5lVmlZyDrh0eDSH
txx5V083uvhpgtDNRgv6P6m+hy3aCCNLKFwhm+UTULqcYVZlFdhuB/PrhQ5lrEw2
/sPIJZw6jzva1Tyatx9GxWPsCht+BrbuGdgfkWuOiRrlW1pPI2qJirkOSuLrvApS
7GHXglWffFrxGUnHLYeGJoW7yPTERtaJqHce8s5h2QsgEKmWBVaLoPD8ozmmVfJq
qZG/aMrEqvNFcciyj/0Na9u3P1cCnNv65gg6Hr0VzUd+/jdFiJ+Dch/zsB6Kozwu
a/+psOTgn+n0fLjOrFl3Xwv1kt1ZsUGPIXueT0Tnxow3VqC5l4SH/so/6c4OGPaY
vyq7MzYVEjxM9ob6DpoIm85fEYBmfsHvLm7CUxBozZAXFHYT028WGRWvvxEpU4K8
z+lyWNzsoGYmY6krtqYA2Fd+ZLyYMI2n+WwsYgXQO3RzlSjo9vKF9FeU6NHaFX+E
PmsYlXr12PYDYk2UJ5HE7so0Z1nf/y3tQTcd8lodmtmLi82/vQNgZDbWKbC6MUg7
exLprIBprDSPOfKvI5ejhNj8vuEqhBgQQ7RiV8IF3PxwpkbQ7jAPpUpFgHzu7kh/
1jWq/DX1z7EF1dpZGYDG8dWc106BelrqXxztM8a8KtPDtKSRPdXytHcH19BlT5fR
D7ZtCwGXj9g18TkwnrsoZO4Y4uPcja5gx3xKgdohQOjs4NzW8g/wgzDc3LvjKhf0
cYLjusxyAw3PW35kjekH2swM5fCQdFz98HrKQAU7ScamOQcAllHtNUM5G+JtGlB8
UqGZsPvkkN+g0Q5k5A0vEfqnZi7gVtqe5vkIH0E5aGSSM7xJepfQs3wj/QXaAzW7
d6hZgVAPeLr3Y2FhWUtmo4INGk+Topk/BAdTL1rPNb/KujzXFw15fUHewlbIiWLe
qHhvccWYHehOnbMazHMxeCJMkeeGrqgZtZQTlmT6jvO41VCKZ/V+atwGboCN1LUU
BqkKmoVrYs+qYNRwd1GzU87TJwi2JrsmQtAr44UreOQOuCGVv++mF5AQYWz8p8Mt
gyEykV/jtoDE6c4feh8RPLb04v6/4C9MeQe3U2Hdp9GD6BbAXr9QnJjSWfmE2JUt
rqpVqBEGN9uYLWHyWjRYbml77SbW9mP8Q9ocVvKse3Fh6FNb4UVyD1v1KZ9mLzAw
vK9h3ldyPxXwv6ax3p6KMP5eX3EClUM2Y5Jv4/AOhLKngANnWdUHWAdm8ZhTK8nG
KqunVufR5F6MzRmLcl5hb4voTv4yUtr9lE5EAHXqltsVUxxJCAZJJdXfjDUcXeVY
yPJIA+nkc26yJMIjfri0W8ysVuUA8MRW+IjpCW0NDE2Qste6/bMwZw+neKjUP/sj
5cOuadRYprTW20Fh/01R4fNNU339hmUEVDS/dGkZPydJIlpqtbJwtvpbO18Svo+b
Cj8vJ+R+qwXLTheD3w5RBNCnJJ/zMnFRewetPEE/NHrQpiYG0zcWIIZblVGuDQ8s
xEbtVSXjwPuT7xj+BjpVFBW5/jLTlT5oCzUjaUKwBiMJnKHq2bt79CTvA+YyiAPY
myGjdVBfqmBFPumzDrvat5uBsBJAjA8NJujYuhRhWsgQqA8VBe7sJ3lXO8KkD5SL
rVeZvDfPDa6R0Yd/PwXR8MQhpcrs43JDIK3qD3lXgWqSeqIjIY/dnm4XDOefkQEe
vXcBELKkx2iDw9ucdD0+2B3P/D2t10HYXkWIqbV43TusNaDkTsJo7M2bUOlu5++9
LemT6m54+BCSv+cmSdHNCeZJ5ueSLCICmbuUqW8CiOGBQer0LQUjtYiIrOB1ZsZx
qE5O5bOjCEkjG0hd1Tp0jq1nJ62nhiFmelI15TLRyvDeNbYTTfDdtqtao+92AdaW
cjQ79GET08xEHKcl9rHIt5nGiYk5WcY0OYbEjOZbzwRha/jp86wPmgK/TDjHkjX5
Z3ORCcCDNlgmhE4TvKI+qZwW09H+raJUAayhk456eo+k4xo6fhM9EaM9eVkPdhfM
NuzVXjTap3tmmvLRqBe+sVMNRRxaRN5waYNLeLaKQYnuTw4M8D1ByQPcyDVGZEVX
dBODFgf+quwNsWAswNtSbUxkkpkUqP/Q4VW12P1FGPTmVcQI+jrbDSXi1IC1cHr0
WNoaKLykhds9u+MMuOqt698d8THFC7xqKAtTX5zj+5al1uSYvUVRCBz15mJukKq/
BwwaanTp7u+UVVVRyPVQI3bcULR4VRR1HpK5qBhGU3Ts20UJsoRN2c6U1SFAGcNu
Irs7GWCEnzuEDCm+19JYsr3Bvi4BiopkIt/YX00BgzMhhqDB5KhhYKcoNOPRyPwx
2cxl8vTtbt61EGgHByWytlLtv5BsroJsg7uQgR/2s3bfXZz3s/rN6fl2Gn3V0Yg8
YpG1Gk+kzwWnx//NYpEkHA6Ukxvhz+UGYyzfxLh9ANjXPsCjt+1gPqaG1tFGYNWi
rAXcO5iz3oLnFcFqw0FmeQxOiwou9bgC4iX4pkWbJenkYqOpE9HTkE2OOBG3TG4i
tCHr4GyvYTVbgwjQWJzzeqHOdSYoWlEnxaew0MLxyU7JLow6P/YUkPDAx8McRYPG
dCV6YXa2PAUBLRC+cDR6rUxGz5lWQwFvLOjxprFpDboqbfL6J9pfo2koF0+joU79
qw6otHy1k68jJiftiC2n9cw2dNm7TSji/pePLFmYFngkW484ltv/oYm83R2Vtf/f
c8hT/NcbhTHgajsqvG+YlEu6JGI+zZVMFhfe1CZqEsHCPpieGkiL/mWE4XjEAeQj
qC50xtphP+u76M4J9igowLbaNthtBrlmr2Gnd+Mn18DEqEfVRTtPSHBsIiOhlWvK
t0dNETb1kil6ny+ln0Sw7lX//8ACdeg7h9OuqnOkxCZWOAOIs7gD2a64E4hhI8lU
y9J5Yd1owmPCm1cCDNQ/fQKVqIhfnojsl/RNje50Qw56+N4PJQjXAhkXnd9gnUC6
2VDN8bhyoG2UXJJtPd19f7w5zlEx5jcd3RlmGcc78iRFfoaZkh4UAzlekcyA23jw
W8elGrpmPngk3xRN+EYXiLUUBBT6l3vhSgSl22Y5CT0VoHM11PWNY6hQQUo57C34
HMNtzBH6ZtqvXs0k07zxqfBkmxal8jFGdabZlSIoYTX+Bx/tIZWrimfsqRAt8e0j
DsxXIqRtCvUgNGv/4m7h9SWYGlfMuDYvVcPV85YNmKc3AEa0fJQlB129gFopWNBI
3dUihT2gt+yTK8kVAxWN/FCex/oqoG6QWRuhPI+18yvWLnZfSExOcUvCzaHeoIIK
C9lShd+WgYwkCMbv9P0nfBvpq1a8CgOM1KCtVkPb6Ke/wgEJGx6NrcG6CLqHCMzY
UwL8d4mMQzezOh2InfV4AsWah/UNWL71xRazDlDVfj5ItWx9SZzqX+DaSsNJQEhF
glSv3tBe8V+cItIIKeJEw6zl3m/EYCRhw+1RrI6ZFex0+Q2qh5GCPteiKbPkaP0z
eP7qf3IqwTcotkYTa40w/MdtO3jpYHGEl2/v+j1oh19ABw/rX89lfBEVHpsa1aQx
A48zxxgnV7tEuBfqgLM0LSObejkLWC2qrWiUkYkUKTltJbqMcCovVc2VDOstSaa0
20xhIOKxCp0X6eD4BA57hbxmfhhIbIejOF9BRIwOnKyCxDX7ntMkQJekIjf2tKWG
jyDQvD83iVWhr3LVQNAUtJH7UGUjVL6SDvYTP3Br/sYK1szHrDQ/WJZuFOCHi6FB
AsTV8/7IAx6TnORX13SHJwKQYIxF+qygFbfOiZ/C9FqIR5ZwEttdYXC8XopDsRxk
OgLUg/TnL9vEH4IYTe7jdAln/GrxlwjzqhJnqypSMT5DtsQodhrw5tqajaT+rz6j
k15nQ7nB8mENGWzNhaiUOq2/ehlHJihP+Wh28QBAdRms9u32nr4EeGlojmuEowwA
xVZqg11IHL0CH2QiNmX8+1uI6cpvG1qtk/I9Gkcz5MU1YXsRrHEjEP/k19CTjjYq
Y9vnbHdZ/oh8/BmnU2+1Q79qHH6SHQpDO1iFKIDmgQY2RLGXNgvTG+zLst/B2Kae
0VaO14ErxnvNAFVKp3uc9pj4HHkqQwnEc2iDCV33oPVDF/Mh7GiJyHVU9dwV8y7a
p/Cvki5EBJAJDvSFAlyhygqN3uF7Z2lqnWSg1Aqfiji8K/x4mxqvhlRCBam9tlQr
ZOKRvevpl73X+4eoUQgs3cn7kAAx61on4QJCUp/B25UWRblgrF2toSfyRiBElmd6
VlYfD+cNTY68E3K0tftU1UmkPhvjKRZsaw5dDV7D3m10suD/oTEPEzfyhbBM0qRM
cW4qw5ZPkTIpBJJoAjs4mcWezoJUWLKKJkYDSePn7KJpamtb/1Jmmr2tQZWEbfti
PCtLb887i0Nl1tSHI+6yue6eIdOgdumRovTU1+hWWgUiHB/M9YxhMLOGLInrKFln
cZ0uuT1AFDEBDGueixFwEOMTj4uuVPahIykFlYnxOrLC7BWN0cw3urDzC7/tiWDT
IbRaKuHkBffj+GT8kJlQNy59Bb5TyT04AIa7xTj5HRU7ad3quaZoE2BUCpIPUwSs
PgeUHevLId8aYwPvhGc6u7nuPzK7EuaITk3tlGJRn0pesijqUlehxP7DrZGeWv82
AsP5evMDp5Ca/uJ5PQ/SagAmG/LlQPKCsTvrjEX2zekq+EoZIW9ZiDX7TTWOMS4i
IbsG9240hxVzIQX6b0n/ZIp4WlgSuP4HzQ+9ScABD+h91dgbQd8AYjFE2MTusnfH
3xjPznbxHRNbzUv0iFoFxMtNZlhHBlGyi4bsntOzWO367mTbJJZ77DnXjtFEWrrm
V7HL5/lzgjqhRUpMgL4Vtu2bTEzvJ+jJIR5wvaFCBtUavUQqVuF1rA3mUopf4RuP
1AGrJZN8RjIKK/8QHUSldofTeBLVdRlg4wniYjTHZguyJJU6kNnmn1VCOyezVlXr
SXR9ysUkKEI5bb98M615OsBsTu8uji4HosSj5J0+/LSr5xOv54Db0E/6CwkOq7Vg
JukrDYQGo63mb1rKvF6yko56xZvUSC5/i3EyYW3ojGvL5NlYhMwG7KwJENlqdKQ0
hq2FGRmLAvSHpChaPCbTCZH95Mx8qTiLrB9i1NDZTokSjvZK97wjB6SaYk4pBX9E
6mCHf25ilo3BZyNzGy15CzsZ2eB7qZraTtlD+L2Kba4th0J4ltcrvkBMQpgau4rY
9VsN18c051FrLkgjOPcT/VER8G/3rymlFI6xaTek1ZR6RxO+Nowx/LXOyUyK41Bv
vlsQMowwf4TmYaO8om/tX+XA41McLDhHSovXw7lFmjZ+/NH3EV6z+6xNgh/EBZLx
qCaXOGBNqioUOLbVWFP+M8/HZg/S3P3+wOc6LN+w8SucDnxCJNgwjBsWOjX3+1/O
/2e2zBLoJY8dpzhPSxFw74zv6lSxtbQrx/q+hH3gFJFN23oLKp/QaqAAUeU7FYRj
dXe3QYTRQQ+eFCLiA3refjNRQvHsQ1uKgO67HQKtbmgslUE4fwAEtHdY/I7WH1cy
ZaJsQ8N16IKwGEqaVvuZv1jW+1Bi6sU9rGJDHLZnBO9vty+YQghkglFtUlBXEvOb
9YMqn12J+PKHUzjTKn9+wK/JLohKwZqPEy2KbASM4MrRv28Vsj++phBh9pe/m1Rg
6SgcDU3yeTV4xs88bRDdVW6GyhdidXIdOr6ApRLPp/PWaErgOtRopi/2mPs1cFbe
6KlhVOsWnCUhuVCF4mU2mSwWHEk49/aOtljeIxSBr2siOwa6XhIMr3dn8aZ2yyiS
l7oqcq2Fq04nTfxTzRSHC7d2CzbjWY2u9WjCKHtj1UVoot8JYKqKoso1NhOUMNKL
Y0vUgkspFVrlAJq56vhRe+YSwZYd0duDkG9+XpcV3PitZxckmioCvdfJKF6C/+Ku
EqCeog/1lEI6zNwwGE/QEJ8iRf6lvqdSUoG1ozwvaMFHx416Hol36/h7JuMxaey3
/AObfPuzWn5vcu9Ho5aXQdiP0MZ0o8J6vbbN4hsfA7Y4pNsNsNf/XPcP7u14tTYx
B+fKaRffz/LPxoDwwo1RgA4YpGTMWHXGli3ofe8oAkKA6sUWGi3oSkHARKUKtszJ
pnrCXHO7W/Jim+ayZ8eTYqwHBZcruCozPTbgnTdMWlRRu+M8X4ofEONE+V7tb3Vb
wHsy4XQ7H0cbK31ogtmQCQyuTHbKyPvzKK6C/YyuhfsnQtPcu7Bpb2TXy7z3W/41
JFtfBsDC4XEACGbZjweN0EnL9RbHsJldW1U7nURP9UxIzaIfkEb+aavIDJukUtzs
iUBLHevic9ToE6mj1Iu6dNt3zF19LPyRA40Os9F3dNEqMdGOF3DfFlKqzr4ntaZO
r7iKt2Hm6W3w+F1TZ7h2Ad/N/tqIpgQQW89VOSVQhD2t8GKoPg6jrphFzIRaP57A
xHgb6UHD0JoaDCloIzJCKQoNO30tW6FyNHAP0FsIlaTpHZngbxeRhe4q1vYYT89R
mOVH2YXF76+hqdz+O9ToQKUecsHLsa1xHGLc53k+z8175Pk75k3no5nC9nXSG3Wr
+PH/5me8MuDP85K/lx5PJtLGB4fqwRPbfYBlfgS+nblFvn2CYgHNPBNpuWKUbGmz
ZdWKbPxpwFnffPXeoHMx3oBoFryfLAGpL1hr/teWnm9L/1gC2/EfabFUhYSGa1hl
rcsBmuxjNigzvLnJZyaUq3bCwU1O4pD2MWSyVwfXl4M9MtjqYCWF1QL8ssk19ZGn
+kmWQnRzoicmE/vLU+Bfg3bf8sHS25iZmwxUcRF4qFPRwNykRHoIGugVq0KVNpfA
mmJ0KtvHiW+v7iJvJNsTTZHcC5CwKiI5N5ataw/9tzSZ/8EQwEfsDX0CRys8NNWl
+yt3gL5Kuca97OvVFoSZl6rC5zWqa/zNEvvH3iB9L/lZOx++XHWn1aRzAlWG0qTZ
us14CEjsKvZTgKVvPEUhEcqadadG6TMJv6WDp2oUDqwpOGIuOXTS8lEU0NatC0PD
OyvoLOwJSH3j7Y0V3KFqNU7ccHDP8aAEjSlcqOcIUZfbb31UDq19H773r/45LIHD
KBtUrz8eScVwgOL+39Wi+EAVOiCThxu7OSHCgrmnSSkFqE+WtSaqoWncGNS6hNfX
/YMOgl5uRnGspRrCVDMMFoE9M7yVMLUOQP+fn1xktHcmbd+MNj5Fnn0/LYiZf5Cq
r4CIawzKSw9NEOFR+GVJdbC0aIwimwWLZNNU61xSM8k8Oz1CYx5gbydiIv4E+7K/
qdeKIMkjYio7rHaL/ViAfIBgvA6o7NE/2HP0sswNe6lk17UG7Dy5SZEVBZszl+zy
RcUcC+iiew4oprakzvbv/707Kz0KCUuEhZ/sOrV5fq5c0Cxb9FS8dHGDTB7TyK44
Xf8puz7U0tiewFANYRs781RhLGZxeK4G7xVzE5UzbcYcxnYgmk0guJ1svtjYO+JI
un/zkWw/cfxwBdCO65/i2SyH20b0BKDesJ8LSsyGPfwaVWJd1JK/e3tds+PJbaGl
TpuCWfmIHVrccEC1cWl1HaoD+qWjr/4PcKq8hc3luoa99tIopYLSTbfgrPrevQmy
6JwQxlanSDv12uVnYPvKMZ5JRXJ50Oe4gPR7c9FdEXMyrU4xTcazlpwjQBy1ckyR
Kva0bCL5/FPAafrk1XoyL/of/sSaiJSzVSrUQQFHf2yIDZb7Swmy8S6nAL8DDOEr
MmAO+fiD+bb6FK3cXL7ogIVQ9m3pLI/c6XSVhEhE3anXe7E7rQWvmTGapeuOvwVr
v9eXFf1l4XKZHb7Wm/U56Xk64btpHLsIA6hln7Zdh22zTk1FFfNWAwUZmgm0LUOn
q4rzF86BCV7TXYClawhrAd6M9q+Pd8aC5AKzYCotUSTc8b6aXuJ32k/LRyXq0GPk
2fTQi8+p2jBwG6doLgVLdOPOsBKvXNDYdCpr0S/u2n5E7mhl1UQ+wuuPWNPOxXwN
vbg0DctwQSUUn4g+ZSd9DX83Vf6nVtTHFyVYpH58IprAQk2FLQH1SSmaWiRwB8DS
mzNVe5LHjvWsSj9tG/hLT2zoTcqJZpykr1ejN+1fQq+ByK4AtwTvbmAoZOoMAwxe
dJDcVv9LRnrScsEXSdl723ef4yvxK0FOBBAeI345EsiTZGFueMQhS2OHzeUqe5Lu
lLM+p09P3AksJoXFEPfFTn65dRjO5J/1oGRiFprREBJ/a5PbWRqBdmMBgmXbajbb
XwZcSt4l+SKJL0vOh1zl7z9x7yZEvB80OV2oGBYOYDDuTbdYkJ23DW6p58zr0ly5
6h7fFd+ugxEzNusJ80tgTAFwV9mxc1uqy9Hxl+UlLywWiGQh2ZRqH5B9yO8kuIG0
j5L/saLFebI1OO3aJMNsqnWWrxXKhmVLfhnuGcr566381NMrmJHUf3iQQjGPpvnU
+jfkF6DZF5dwYJebbmryKpnGhy71D+6F/twgITZ+CB5gJHD0H14ZRxKjAu+tq9qU
I1M6UuTaUn8rNMY7GTOP5L6d93Ih3Z55yMIamyMg6tptYTYlRuLRfJ4Jl1Fd78oU
ykDE7Ic5yZcR9uga2qHvzF2IToUY/ZdmUaFg0I4Muq/nIVwEsQdFnAFMcELe4fhz
RMlUltv5/XuuxcYHByI5lM+aMhkQbG24ToaI7N+zY4IMk4PKukAN5lEXOX+Kx6dk
4SIM4lq3Ohxs4VtxgLRH87izpmLJP4nRrZVlmPDFf8wHxEX966y7YPra633J5wSF
csHGmcMMxfL1/ARlHTQWN4XSVF6zZRLjVZMhd27rYTCHbCdQrnTh2n7Zi1aImKQL
qQKt1Oquy7ZkNdC+nxGXBA+gQrchTG3v8Wqc8Bjvmm5fH0rCsPNIIokqbChi31h2
Hgcv/jBeZo4orm3ggMhNU9qopofKPswE4ae3X/PFPK917XKHTLoykSZIpGSiuDZy
htm4Vc0QkDUf1MRxBcuGX9GuDZ7c8YhIRp629+MJPlEByvwETbIfty4sxW6qX7lo
2OfUhMcg+MlxDExFx9Qt8kuUcDY9Ye7N4mO3zlAxwpioTSefEbKH7v1g9IJ9KJqh
0+2hrSODjoVKA3li41EnOQetFvO1GvRY94gOXMYlcOoI4ma08PmYqWwbleyHR05S
TWcIr3D5Cw5BgfHVKv4jUT2oiwgOSI/ydaasabtpjXQHpV5MlOMPwM1L6CIGYutr
Z9ghK6icTewRKRY7xzIy8rY98oiDTh6gFXjHzNEIdW/n3sTTtBjzHsbTp+G/ch6I
i3pl2UTTIn5+OoyHmI/ouiN7PnFMM+rXiWJat1Xzvvc7xeE40GCrKu4U1YCe0seC
6Cnan2NFGVMUZFM0UjJC4YOV52xY9C1NiFgaKBraaIwjZO7TJh2eOukv2pr9XMR2
pwsef4+vqdgTFntfwmGDvaItFLE9tJJBqPVQJrgqLuFiLgZay/KrHoGI9enOqus3
CTteycBK6oIY9daaM+Ka/S9+W26+IQuSUMiysnhGgGZfyohRhExqFWF4L1WJxc2S
okDTbmD1kqpbfv0Ca2+6GWEN+2GY5Rx+++ad2E31NlpbgRSYyKgFpuuFW+85Dj5l
LBQRmV6wk5VWXcjAsMctKcM8q0w3//vKRj/qIblQiNhQEPoy3gW31o589c/HkYq5
JQr5eHfOfSrWbKAtbWZ+CGiTyr0Lpsv6ICLi3qmZgEtfZCSUsonwx5g5qsJXVpQT
kfHYtHNOS3pvuZ4bpN4AfuQBGjTHMQQu8jr5GRYcoRrTJU5Pek9z6f2IBUQdzr2D
f7U4PQpjKlgq+nIqZxGonJeUNVa1HwGubHSyKfKZ9q+4wgasES0lMbBv/SIhd9v8
vLheT/6QXHTmM446C7wdHr8ba5EbHkp4a6NAeY4ynTPwnoz/eVnuRk1nWs73YX2D
iFp2lLUsuxJbyVHRHaYUgrLRNguzqCcJKHQaILaXTlB7ocozVR1BzIxil24SM8RE
IfPDaUvbwWEZO5ZMLa9gzObe3pZuK6vEqc1ooj0mBremC3hMYaPRkchuY71IQNFj
Ep+uiPa9nLVRinri03wKLG60TlUCGAZmSbTzrbwFRxymomsrl7/io73BWcgDCWwO
VGhB1R7bXMEPjilcpEX74UTYov6Ko798rWMv2vliK77iAg3u5bLgWwmi5KninLLN
myZuOwutoFHDj1ztHtspHuJI1yQAGtAYr+yca1Prg13GP0FcMN03euKFq0iJ1NAb
5IWXmYpBDHH2PsE/lfg2YqK0BGVBggzOMiDXRoIdX/RskI1dntL3N5ck0r7XZyCg
a2QcqVMxmEeJsquwbbioYoi2vq8IJq8P8CwWqeDS2YAD+AA0Clj3d/jViSc0hL9m
DUOZyjCgBCwF1PG2yf614C+fAQve0ENbi7GpzXPAr1+jjsJQRkX3LRpj/w6iZYKS
yYBqnc+znVbx2c4u9GTjIq4ZvLzBL1bVeB9HEXzyR5IecSuqPAu2b+jbT+Yf8rCl
k1s406/dty6VfjvayjLcqqwpv85wAhYSzxO6QgssZYQ8SePxmNS4axdevQMf1rAs
OWZk+r1TyuOD8LUr9aFwZrXsIX2UQ9ZCEo9yOBDlWZIjMyDpMCuz+U+6W9XHs11l
yHkNAF++kTC7BxXE/MKmfYU30e+am22QLxQgsvD6uzL61pnZ+FnbVxhaPiPw3u7H
+lqcigQ5w/Cu4tNd3Zz0jeBBNU1c4v2hEOB29RPIokKYpBiOAwiHP4TzAMVk1kOb
LHxpjjoY6Ai2nK4aDv0H79mT1N/lkl0aO9G1/nt15KSEadWgNiThvU85Jd0AucWK
nmcM3HwiCAkSvX2AInXiuz+aNrz8JtXo6ogbwQR6OkFBbE/dqkBpdi6HSDGQH0J1
39wO8Rub78OZfP37d0yNo6Bz8qZD0JMq+GaHUTWOp1D78MzwWYVcG7JeajoZqArc
oC9QPQ/mGoLSIcWUzuVrpztCrAgU1U2KJ7bXTOQOwXEhcAcymVcc0yS/PAdG/P1H
IztrjdHglkrUvcIngdNFD5+FwWM0sf3u4tdVzztKbpEPETxQukxfRDMEHJIloq1c
XptKs50keUXOPJnGF+CSXnnDLYYP34bgrpTB4E7URolR8ucHmKKYhxUH62r020AK
cSDeUx2TjL+cGxml69ksHTwXH7Krk4piDjuwnGyMMfRwuWCbZnfUWVU4YTg/7FDg
nQPGy7zT4GPfvzJVXARTlk3H7EdLG6VqM0Sl6CuMGRfPQV2r4qgD0V3krQ/eXE2K
MO0MzEDCAoEZZ+I+surWeBKWh81SLokb5wMxjc7jp+KvqOp3xD/V0nDM7zfOTIRk
g8JvYTx1pn7zQuBsh95zk+A9lNG9eJIETnpPsXo/oNE/DGN/I+oKhvxYWQ7PfDyo
IAvqmzFrxtw5lmR0k/SOVxb+SL+BhNtH1fQrN2y89gqxWXbbJwutLKTygyxIFV+D
ZsGLo926hRQvGgjYDDUk3lr18HdxeAi2BXWS2n/dGlVBPgBGwy8IxQ3zUKGxP7ML
ciwxxelx8OL5NJJo3XU2/DMdFSxef2CNhqqM1T23uYz2G79sn9oiSDBLVSY1kM4W
RHcnEtFfs/H8NMTINUEIb5YH/eXLY9CqTeScPwmCiq00JBC9PW0pi9sbPqaBcJsv
YVinBAG077IQ9UPaXwNhNnuMfr4BPTyuCXO1BnoEoFt5IVAgu3Wq/QlOdXcwnD4+
MRFO5tQQ82FtDuCTJLRcT3iWFPV0lFIOQq+1eg0LFcknLiCYP8w7FK7BP7PF1Elc
OqNc/7ViE/ndQoBYMQh0qHbEw1KbHBuERYrhKpvwIZA++g01Cz6o2irQ2uliGUWR
M/olCgZ+o8jhmAjEJeb6x6ohXKsuqTAPMPE9jmkRpD8mkqOm2gIxD2utrpPn9dp8
8pAQFu933sIRJwmTZntXdEdZ3tUzokE9s/Xpe2ctsPVfhbh9y5f1t+F0hhEVyq2K
nD8Wi32+r2Fu5+EwfzAiP+YFOWPsux3KHuSAi9hRPRv3+CsoWo9fgwoFwJkLaT96
C9JnunqTp6/V/JDOZUSiy2RUQb3QFYPLrNysBv01X/SrTp/5/GnOwtEK7fy8xXHR
8VacMfQlfhm1EcVrXoEXtN2FUflQ5bBVMiJBGZ/0b4PTHW32DAfbMA9yMpRdW9yt
`protect END_PROTECTED
