`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
CSjU9OR3JKnQXDIKEbC45c1AA3SfuzBwhcEQt+zw7WbNuqlGQ5NyfBWYmU+HI2yZ
n5yTNmDdOBKuTYjYEU83p7MFu9mdB8fN4PX7Bh13TOEy2ZaSk1aWItwi7ScQ45QB
puSSzFMfcuX+m2tpTjF4l80XEyGFmZiiktggqCCrPAax5uzjvA2qGJmcDffwBbRc
sAbb2O9UiUcNOiVF7d6ArKiWmPvfcerPR/ECpwRB7OlKtwVTtUygvlYF3TbDnnFl
ckTAmi8bxDwc5JTn3GtzX0D7b7GotcQFMa9cGKcFgBSRuqNpUcuw0nG+YgGTmrnS
obuEgyH/Z1NK9dSOh7PP8gAFSxr0Sb4G5+ZgiLnJsX1U538fptvvxN4u5HsFs8GR
/bY7fDFuhtw5HUvVmr4adDd1c77QTq5gkflJwnx23ZiDdhELeFetocvsplL/Rsj9
Gd2HScd3LO2RQp7IgWs45ektgLqr7od2l9/sB39/l2iASWPfL+e5V/EqFFmZb+Bo
vOfnRPU8o0VkuM5wOQsxz/M3wZjVX/zYae9gPGQD8tZIWaD5Npie73su5tZ9T8a6
9SkqdZjMoe33C+GQYbbyAfSxbml7cHUH3cc5+dwkjHN87D5Zg3KGmE3MWAaL+3fu
uVasmC69AB7kKSt2gcKNp/FH/rBCKeoSj6htxzGaYOGS9Mt5/qToPbMDF2xvdzd+
gajQITjp4hJf3WoiYu8FyL/1CeIh5RlXkpmt0vrD7897Skndb2ZUZ6ee4XN9sSbp
x37CSA3sLNNEX+Wz51TQ66/tKWGD2KUOdqLJvOxTRaBViryp3AvGpnrmjYoK3E4G
0TNzQk+ePqRf6+CtMvJObX7nu9V8Y18zUGM1Rtsxdf89KReJxmuvahUsj2p3ERzF
UMEydZ+hozt4bEo4KKJggowReJN0tOpRwcKMvqr7yGjtPyRa+GOatTntoHMDUF5h
SdelQx+inIYCet2I57zaqA/4cFGjk3J0xrFE5Ic1Sd1ObdMgyUHgVVDSm7xLxPQL
aFU9KTj58GwdekbJNh6F1tKH3U8G6f76PnciYPkiVMDgTz7fmCB8c0CB322/88TQ
oLbXq0jzbX+LMYO7vQPwKFXeUzL8opI0IoPMjivIAUPyLWTsHkT+y9b29FOhVA8W
RpjAwfduLkPkRDWVQD2gcfWDwk5uTe1Bna8KOEAPhAa4s2U0QSaytBaPLnPBzdcZ
25p5rsjzC4xmHpvvtN8f/RONCoW5MnS+5qtdtPUREy9zojPsUScRWVARW2Ek5cHz
9S7tM1gT/Ona4Ze6sCBuLsOrx/hgkPXO1fQ6k6tW7en3dkL8hR+oFKzphy1QgR/Y
2tt8/00OPMigtmF+5sHIgVruljR2bbBK/ylx4MYGKig6x7Nm72hccIOvGqhHML+S
A2EbAN6tdnnOaikFh2nFwfetYU1G96y29cIu85P2THsOgutEOdnS+tWBK5gr4Ggu
/O9lXlAwjXHIfgevFhiQQtvqWKBT0Xg8N3LjpmqTgvUNgMDUT+D6ED4p+JdkXlk7
sd6vAiR+S7FIc5HbqPb0+aQMqY5IrOULO2eXfZ6L7j88UW0NucuuefmmAm6zUp+7
lpDn8cFla7ufvMOhK03lvGpyAq4I8DnAlfXPP3/9TtJlKsYNeJ+BUuAYUzX30MSG
emu3Ith1R4UNG8Mfa5vU8InsN6o95gXX7yt+7yuMtTvumUBxXN6qaNNGcuZ9ai35
ZiOdTc+kT0nJ6QPBuYR9T50zTk3FAfk8btkNlj/lSnANw11KLShSdv1Z6J6vzvIy
jVl9GYZsVKW+ZYx8i7KIu1VJnd/PUAwzgsLzl6/+P/5f496aZ7tNRqIzKnD3cOn1
X9sDPVVM6v4px4xEAK5Hp0xjv9Br4zq2Jit1KBtZ+vt8rIEX43xu9wQnrDd4R/tl
OtKA3Pa2o8/nX3d/mRr/LUeyJR/6XJdn3qU0RvFIEE27eU/NUdbxn/e0eL1x6Aay
ZNGkS1DtFTWcA4kVmlcp9XvAj8CVfDh4/2K+P99LEAloh+iehWJn56eXeT5O08kU
e2cqOcw9pW2KfDslVB4749UyOpjBBzWX26VWqv1wcL2wTZEcE2LmNLVbHJf8m4Gu
aw6LMtdPGQSv6G+CNKPT2KFlKhyIMUa5A4pCQwXhJBaF7kVuQGjY+D9YwdBOVoPT
V0XcsUKmZF22sp4uAsXi8zSOM/zmPyX6a62wHh85qSuTfuBQLZKC0m6b1BAcvmVg
9Y/ESFTVBvjthTMbsdnHiy5xmdJWYfAZbsfzYWLyvtJQy4dRy453PqgLSLCQEy90
DI2FbYbk3duMhL+yl6oia/PhrqtVJ/k7SL8yzbwalA0aAkCs/YuVeCTaD2z01Oqb
7XwVGpWeRkV9rb1XMM5c4H7nW8lCL0t/n5OWKdNqezV5fM0nC4fJd+BdPp8oaP+8
BfTlRAJPSUCZYOC6iRNnWETZLqncN3+SDgWW4H1iqTGyxW//sxOAUHWrUNdrpJ6J
wxPVgU+8G2BogEmp/HjeIIz/iRWKozLNl9ThGIHXsmfQXmS9fI3zBhNxkNfjGk0K
BSnDxNGSJHihTjkbHLpkIWpWR6EtG8qXrNYHlUI8YRp/9Z0IEhK4mFrPi+U0tKtL
ZIwSVAtz7nLuq7X3vW+HzQh3af+q04HKfj9gku0VGIL/8/v/tT+alIjFdVkJiYY0
nL3f3IF0SHv9pZQd5ZF7LrueMpePu5FJU23B12BEWwRXBywZOqCIGitoOWqjU/6q
0l6m3ERw6C4mmIdTIoB+1dd9Zr2HMtkL9UsgMF/tQUjpS/ZEIQ9j0+QBz1wx0RNV
y2vWjJUVIHtbdNRAQ5q1P6WgMSQGe5Cewn6ubdoXEihrn3dM+iS+vVPF/jMrQC6N
S1HGZn6+sNcTaMW3OLH36D2/02RMCbNm2J7myRStf36JZ49KNnFT2WoK/7EYuvsS
6f8oytHrPlX/8GvaEU0VYzizjoEbBxAOLDZezGaobeNP2qgrBvifKDnnRCBPgoA+
bKIVs389EDXyFGG6Y16rJfDbG0chwc43NnPdVewDxMtX7vINckW20YcaxQGvH9Im
oiRfd+eoWiXFdVjfUsDiGty7NBYyBu2CJxQTsJjZl+Ea8csNzJ4PPmN5VWaIvsH5
+DsCVzRlo2nIGrH5hFBO+JPbS+xXZcWEkAFuNwOnB96gWr/He6ZxTRtM2EpOqMzf
yBHt746vBdkQTDUC5HKJ4UVFlDEj+/aDRaGvu80yFFCSn0ctsfdf7ohDB7rH6TwK
JKSuPq43gg0QW404n6rSQQQWBF/ZgbiJL4ZLfgga5UkNj46EyVYjFcSvIuFtFRpc
mQUi8hnHOv6jk1Xe0IpIzXfrv1bopQ73M7VsMxC45Y7mWMcjEBcKsWkkfNUapLzR
5fBupc10IsJSe8e+UnnGuy2s/ny19zQns+yaT4irYLM/yFWYYxt/Q9bKSWFRGPgj
5krHjGf9oTE5XueNg1jg0CDUk0Ump/IYiDuwOdJ6AKL2yqXU43kBPUJ/9pGYYpGI
GAp1H+SE61/gvXjOR4XXOAGl1Sc6wwApATZheixgjTd/alNhsg8ZWdCPBYV7vtCb
DAxKuwqHLaFdQbRmfbK1DYBbNVyOZTovnwfU3gtI4ebVk+tx7eGGW+F93k8PhA/N
0Gn1GShxCHJWX+cd5qa1Hnbv2tK6/NuAPLGeMZcyVXCkYG4yfq9H9ligDT6Sq2qF
V2HkVOWqhCZHOrNPzhs4hIBYtEnZH/PowNMQqwSOHlMQhjTo4NGxHWL5sBjqnzqa
3oTTRq+z5e+0mBJkY1oUHWNyPyIB0EWyq+B5lv/bI5NujmhoKP+bmibJMnPRgXJ8
sbJIQzSsNX/NL9B0MWG2BmZD1p52pS5+tT2/iTiM9atMbzpIRsteW8jNazkR4FR/
AOrSaA89cohxxT5L2eJInBjIorLrDZ61KL0x28lbnX9GIvU95ZPiOeQ7rhwS2i0s
p+J+r4j2O3rCpmIZlCNMntNU7yLm/ik3J+pUtgJCg6sJ6spdf53HuWc5+sbZ3TsS
4bg1SI1D1zFX9ELl0+OoJ5HrmnEYp0w4PQFsddLZvd/WR3uQS5I1faq53ZksdDkc
23g3Zk9ZVG8ZxwKmPtoK9aaNpqZ5FcY2rWW9m4AbOktpcQohq7PfUefi/2QJjQYX
u/16eEtBWSnOy9yLdo/aHrZqxFPrc+Oxj1cBDtDnlVto0XedzphG9Km75QFgSe8Q
cIt7c8nL82DLWJ3R2CTC/FyRalLVORFZ6cj6XrvTt/J/Cr5frUnixJ8V5GCJrC6+
gIuxZ7cJYOhn+4JPvFEKyZJ7r4r3yssQkndH8oLoVAzhXaOmpFnAcBc4cWtpdLIg
cA/4bekGCefTtJGLK7HKANijp6VH6bUtZZPHJ/ja+o1ieZBbPSTFfrE4i6Gy9y2x
IOvuWvtJrqO62qXwCkm1tXLLySUlQwVcXFcYij4DhqcRBd4R4xfL/lei7buVJZ06
SyfFxMo7IXvlSev6PQJFrbggJZDsXFVwWQmXb0C+ytk6ZE4qo9UBkKK+Nfsz7LX1
j0LN8MxoAve9kxkv6Hd7CxswHC94xXhJB+AnXpqb55O/nz8/wlgUED+spLtmRVnc
ZVUSW6Xs30Qg+gNL6zQoaMGZHlVQ2ZpIYYOjVSF3J5OFTWNT1ENF6JINZrLixna3
VmpkcpTDWwjvHBCn9TkCnqMLkZBw+QXhZGx6mP4u29wOq+f9AyFWK7JJypI3+4aB
PNHoNmKgu1NHvdwJ1BMWNhSeoOgaZC4XnR0nHAyvZXAPTY0BVnwcniDh/xRDp++7
wXeovLzU6nfCVNXl8bnGlnilTyzLc2Dy3MGubBcBuCWp8B1DsvyNCnDQGesmKkbs
MoLfkL89PE+LCcHRtmJp7eyu1kf/u+d+3tw4DCYXhiXcTXD7feQWeItmpQKQmenu
rLE653GI/xcq5dbvzai6GCPerHfrlUxbmFzUSLRKRQwixh7kWW0oDBwjek0eTlo4
MMrzmrXf5+tZc7SLPRzBqZhjdlXg9mpyiknrrzYe7/Co+KEydwcdKRO7Nwtm9pI5
8HG6EuF93N8L41rZ/WnfGvFmqrHrMCHSW5eA/Wq1pIUGxpEgYBoU2emnyM2Fii/3
udTHEBQ1qM3OO+5OTL2/+w39A0f7gnT18i/x5uX0utUgY3T9eCTKCNCfOXot1fdd
TZlgPHN31TgljsWfzMfqMXd4jygddeKVfykMqt/0aWOxVm+t9EtgDQT4Ydwxz1v8
FilhkuqZ46Yfs9HJycuzSVg0Kfg7aAiqLr2w+BYxhRX2VSvoqw7kBMQ1lHAus/RA
94fmJxoY6bUjm3O/ogBuKrNkr8xEHIAuNOwpHOJWWN+SgSN8K4OGNyn1owAzydeT
g22YYxmkUQlrPrTbalO74K6zF69go7Pn1KUjmEPqiR39EiVFezRuZaKiV50K+NYP
qbxnDo+UzkcsdspwpEjhSUqtH4KkDUpOHWadU9dP6ZP0+7eX64Uj+Mf+E6HFCbSi
Oseg3d9uiQTPGvDBA/IIFr06mcKOPkprEKB2Uysv+UUFdrHp8Sk/DGDzgT7UsKJd
DllM6l0sI5nVFgeDOsr9GaVqsjA6o77LSVU2qStk9NTV+o/o47s65Q9pHEZbIgae
vQvJQR9I30S6HEcLXe+Tp+lqjKa3Qdjd4g1BUq+9pWy4GHqk+lpTMK3e8fPlPA3h
`protect END_PROTECTED
