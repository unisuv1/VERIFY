`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vecjb+Iw7gFtrAlyct7l/zzQ772pz9DDPGct6ZHNktl0pzJ42bGcZcq7butXwBkU
Q6S3HvtzBw/bLEXSp1Um1rTm9cp4IeP+V/r9/hfFdgBO49H6FBmvRH5f0xnkYXft
0Ru2hcTNOY37+aRuEv6UK6TzVL6XhSZ1KVyCehHl9yQYziMCLOZ1XjneGVJIq+8l
1j///pwenle5tIdJ6OVeUkojuvmT8lp/PCxSzyq2+zv3x0NOmLdC7iDbIm35eSXQ
Qet+0fMz5jbxogDwOppzhG0785OKBNtqAzYUH8YDQPFDJiOA/QBHqU+M81xJwwsu
uSaIRMDnCSyvIAMNMmO4W9un3qwV9OuRygvCXoED0v4C3xgLxHPIT6ooIhbpUJ2I
HuDkVwaBtF+rc8A8Dp0uBTlaEgYJNrqOfIToQ4+IWXOAjRfO/0GkecdGB/n517bu
+88XeRJVET6VsSVLn7cWFzW0EUJ9IozNyCJ3DzUtLP50b7olhwWrjQNU91CxirzV
AdsaTg9CsqEy5QJ1S6uUOPAzDbcU4kb7OW+RUB4ydnl0WG/0kU4J88ALJAirTYW7
mtNKyVIRajoJi5/SG8p6Ci4gbbHxd6njmY/6wyoM4Xfv2oG/WAnqJ9oLKBXKj/5r
KpECBEUCPywvnQZm8AVOPTlrgz1LQFAn/Q1/37iWFhUKjYrjb4f4YGA+lvGXfk1B
4YNvropR1laq4jAT4v/g8lAwHrQj1nq4c3yJ99lWZGpSYEg9rONn/VWyePOKaR/m
wm9LFiUJkb2EJKR34hXjpP3UT4oXeqzGcs9d54l/5K0vU48cxh/2lBW69CsGU8ft
Wly1KiYkfGCdatzH9dQGTA6s0kAAQYG4H/al+hJywPssoNn5VAkI1RExmCVjOfB/
DpCkpLupuz/kjesaVBAF8v8B51xr1O+EQWfqTZIjfYgczHJZi770FdUXaq/iCz57
qecySrNkcJBLX3Tj9oDn5uA/yJitGVXGGItGMaPBPdsK+YaSnTDrKO0slX5lSOT6
smTzC0YCOuLtjs9u+FFjITqwXhD77b79MwmzIKt4gcd/Dh1mt2dYgvgx0SDoF4/y
g9/fx6m+sOLqpfsvLl1K10ZpDVnWlgVsrclq5qn1DwkUkP+OjoVvhBmBxLKGC/Hx
OYTMT7E0izHVWkrpS45rA2ZU0roB6KJY3z08cGHBBEXtpffzry1p0kgmadL+xnwx
zq2DTWynF188sKs3C+FhYZuhp6u1bU0nPb8hRc+SoNPqIWZIUityYobb+JEO+LV2
vdqOVI+ckM66U4Qa505Ub1VSOUpiD4vwK1usjaxJF3tsg+YNbAaTg367TSI6EGu2
JlyXIrzZqDTnqtzCHhvxA/va+VQ3MVagvQHEZMNWvQb51voe0ZQRepna9cQu5lr5
nOqRjyJ86EQcnCN5224+UG1vL7LUTjrb0PTuH+EAFbP+PYTj1+ObrrMSOmNXIoxC
QbBDpBiBTqWvlMuzlZQJNyAyx6xUU0TAw+duLoNT0UhcCggY+UYd7cG/dv5QKdma
1MQGLTJoUbHvlwYBy2NKMRweSKY1henmlTDHPiDJdj1Yjwz+Zdf4HEaGUVHAWuEa
DW03KwaXoqcTby+EsFc1ytldMmhAsTRrzcyLRj5+0w1SuR2+14mrsY0yBMpTanr2
i6S6MlrW+uS2vEJjh+yEpYaJp7ojrlMmVaphgtpVywsmd3vGab7IKMHFQZlhxK7W
d+WcGLvruqYYNoI6y5zCDHz3lofeUDGcL/OeNZl3pYcbMeaJcBofIJB/2g889RjQ
XG59QOYRC9TADhtYHWKd2bomkpCvTCh1kS4sEY1Vo20ohrwpd/m6M3kuuMe/I6yw
BeDPo1jD7g4MsEuoLdxi2yrRAXJ3QVd2xeP1TZv3yimJxxV2DkaCPEdUyhNMP64z
LPp78IA5aiJpaMktOECPGmA2bfOfcGH/QqhvT++d40AwDj5tmd5jYm5+C9rB0ytZ
neRm7jWCEUin7VN9oBfbcuWHXJeEfVG+UObIFlpi/0icXpd5jrnJO05M07gEQfd7
dTqkbUi1+yJp8bFCCB9TXq9/HdEJ0QObB8Fr5+hxAtJr6b9wshmvBfP6k/eI1stV
C7WfrPRlVI5MbfHBrGgRyfwMjc8ouplEaz64k251y5TNiEuJuZwIdOhjvweb8bqv
n+gSskkKTEbd5f5V1P+O+xiCXvLd2lkCKcFnOq7l56f4wg3X1i4d765eJsef874C
Y1FWS3m1rmcQhPTfOwCzuwHBbMb2LoMCbB4J54P1lumNbRdgFfs4HgMfNdkPDs2G
OMp9yeMMUXbULoqqg/qBsFEdjVlLQUZvv354DMWQ6Fq6pnFDaxYkhR2rqoMqtvW+
mB0utRFf3QzqbUtExwGn46tdoanSx/OhIRF8rhA0MfZoM2y4Xz7L8ORbBcvreM5j
mD4c8DEwICCeS0OTQf64o1bnRHqLhIroS/jLGX6HWp/AehJZq+mS7FGsRIQ8KDrY
cpNnzX1oWc488lvd9MyT8ruLU7iMxUzFWEq1rvxrufMWB8yxjl8Ds/2pFCTdydKo
44z/OGUgzDmydPKogDlTtmCXa2YUYsSMwVZ6jVkN0mZuk1i5gEx3Ml6z4K8jr6GU
7GhCZR+MUr24m9zbGQo/kz+3UaunVK8DAfLLacs1sMZ9f1yF6jvTGWvgmm8Nb9k/
5eLKyQic0WTI/t6jaif9QPsdz9aDGnmuTZpVUvKTvppDiKg6q/dZxWEFYGIbNY/v
MaJJi+HX0RnEDQ4OGkTSQIEC60PG8zHxytGfKhf6H36SIWgpoKScPqFpd6tfQsMQ
fHpIUiwThpx4mmes7fd+wu6RFwXzLKAdaCqcWoS/0KCrIq3zBlVLHrJT+9Mtvct1
0wj6OwdPasi+DvLEkn01lcmRQfY3wFDUNp1nuDpu9/Etr/AjrSyGMZTM5cBeSIj8
P+J26XSRdJsfPdA9/1yR9YdlQRu3i0YjXAMUneHJ1m11uyOl7kKpSh6zDVyBcb0y
T7cILeSK0Hrwn59bR4gX/nNzq3DlcGLr+jr+FrBbP86j/5/kd2uRZiCeceZTe4iO
LdKSV5GL14exRuj7+4PkL3lLTsZk9chsvlxdm3e9HsuWpjUyYthwdLx7Lzy3R4j/
XJWcxRyVECGch74tx1Azy9CsRklKg8jhcWlG7LZgJIjXY7uj8DpBZesSQFFI383m
G8udU9KUKVfWCIbzg5uOeZLDVZrpO6OIEoImhtFVMiyrs0+pEQxDMm/BxGcOD4V8
FiYvcbho/v4GZUrb3+1EXMy4UvA1HJf4UBSC7vaCNka23nYMMiHjfAzoVlAUY2fQ
UzHL5pwwBvK8HYEGVgaMhEc9dWjkVxn8krRej0cRFLf0zfrgf97Nd/IPbnKic3gp
D2Yh+XDf6OnzZT7iMW6+0Ek/Vlxwc5v7SZEqWTvRMoDRhhzWuCBrT6vj+VAtxbSG
INxrbqyWSlnY+484wO+WEhMJAIP7ejhox07a8wVwNTBcdPBpoJ/oc73YAOdn3LJl
YNMx6kaOmvnkFzYcb+ydCOhtyBeBee+Gp0MN4sdtDkLk7BHUelJCKhVAFt+G7GP7
pCei3MSxsQvdXTXM1eOBrXGMOURdnBA1OFJRKwdxJe8FHjM5jXnncFIlyB2B5oty
8gBnc0mglUARdYRmFP6Op59u7zI37fU457hrPfW4VbUnAJoNGKo5gqodwfs1viGb
bIbv1mQADpEkk5q9IYbS8ZPAGtxsTy/BFTB3mOZvckxkrMnzpMBzM7P+MeuE3p00
xaJ+aFmrlT3leU0iKDyNLRN2AeOlOsfkwmszfOmFigTWQUdLy5znzZKBFldtossF
E1Dc3tgp+mQq6/7J86otjSdQIGjasC2Ch/6gZ4j56cpHRgpBdix0dd9phC61z7Ii
zDiiqStE2Xecvk/zqgGEIC0wybtgFi0/dUSNTLgqluL7FQh0JNLBegallcblgRfq
K6QSZ+eYtKtsFZgY4ntZO4iXKzmHEm/aaWZW4pn1uxZhtes0p9LHLasaJFo1ognd
Gl9RFGKrK8vvT2qn0rvbLMNsJ60H7DhBhKPncMohqqRSN3cPR3t9lWIyxNyAVUmS
15nvYnP8PE2G1RS994MSqkbR0GkaPM3iVo3vzEfvFeM+dafdjaL7o+KWw3MuQXaP
3wjlurAzej2RrwsBK55beHPjoBw84tYyUKKC9ekrf15HDDg5XMSn4+RxMYjuIzqh
oA28UqV9Jvf5NSiubWN+MkfZhH/Mlecp3wRERZAAV0io/GgEa8DpCA1eZ913BKLO
x2Rmpl4iP7u0h2p4Pt6xiS+80OpJqnsMtm0anHQGiv+RNbhjpKNO+2Zv1VJYCm6W
Pm6znnjzTUb4dzlsKgJNbX+XRZdAfhbRyG1GyJsX2opUFiwuvv2ZVPNCMdRpDCuW
Y5E/oZ58Gv7ZEhBbZ71colmRdi4Gcq1XgB027m0m0g7cV8vG2OzhdcYgWorMTX1c
g11vN2eFKL4YdR0XQ2oqt4eKow6tfnJUHn13jMTmhsKvwAU8oebUxzhTqCHY51f6
elks44Qo46qk4pmtFBr8l0f5NbWOqQItWmZKoBrq0SRcXh5sTIi3qfX8NxGqUcWK
M3QjIMNwH+MNvGJhsHRHhok2fhrUPGeobC4ZYJTBEbM004ksVp1n5kZpPgF7OQwO
PoT9ALyKtZqidK0aoG/9sf3n6LEUH/zBEz6P9BT7vJnceuXELXEIdo2dApQq8S07
SgTj1GbvMf3dZZIOKVz8U8bqoiqyAhWAW5Qrwpx6KnNqg8GmldgDfwxC4N+DrSLx
IEpJHUi9fbuyUugGkLXkNYfkGSMZbnRWRdoGSL5v/tTMxQLR7GFVa2LLBY9LKrkw
aHSWedjD/dnR8nPEWRAHOsZBbw1nY2wnnv72/dYDBxCsNSJi+fPAeD/Cu7Tlb7m/
NWUrTfUpttdcBiQCDBvT6Hyzg2vn7VZhamf356gJeNM9tfTY8eudyXezYBre/uCx
ULlZDsx5j917/x9uKgZBkjByfJXSLzC9eqWUyD4doSRLSY0O71rfd85Jt+nLzCzJ
Sbd6FvsNpwessry6qWIzjuxZCcBfYklcmJ8iQwVZhv7mn5r9N/6+pi23MNBFIERr
/fBINihH2WktC8hrLVYvTWVaBM2XC6oDIs/H5QRn5qnNuoKtM6CgLsecpsSvSVle
XDqT19HDWe0Z7PlrNb6hDaadyC6HdPMSGgu7HLydv/lSpOtFkp8bWLRkN4SRraMK
YKDf4XO8hGN8h2PP+HqB+AjtL8f86kq7UGWDH4Y9oDPnGfGbeFqkhxsgtkzMswKX
+HECZIGQ20u2Xkw2c9dshWFECJVXeSEGLPIJG16i7KMVHy07oYlEzdM1g6VG5Fs7
bLHukJs5HrvFo52YTYoCKUmpFspa2YQI+NQDR3e0gC0r3GaZ2GR0B9N6JxPHdD/8
UvdXhKU6xMtbDmpRY6pd3X0V8VSMQir/b/jNVUIMxE0YJNa0tdycIBq3HIViT6El
e33sQIHJ4/xMImYCdwJprlJR2kww9KQMuEd94khIPwzDCx6LYMCvtOCSHsBf3Kiu
TxyD0A0YRFGw3L87EV8ELIJvghRsNy4UMevJEO1ozPtw68R/mx0p8Cvk+hMiokQD
tb2MlnyingGvEEDc+ZASeqfVR3jWDLa1QD+shyiVAZfZjiehGd7y3F3vTM3h2Oco
G+Yx/FAG55gyz92okheRsB2YWXQHhNFdUb7Zlt7dWzNSUIOYiIQTgHoF1HQ0ZULw
AaEPqxwslge4mPt6tp8dH4Cxxg0gW4pWVlUnEqdJr6w47WFnBL/MtutOWSA5mOwX
wEg88tH0C5ervGahFIjcpa1NQXUcRspkkJgRgbMTjLnye6UGEcr3+ebua8r+mnyb
vSglc4+CnFVWfgaRssNMymtTYDtV4VXBs+ZDS3hffFbUZgtWJr766YSAR9CclNLg
NoaiHlRpdzC1QJ64Fk6TwNFw/2VLspE7T0jxyfT52CG3QIwn6C+Cn1DI03eE1cER
m6YntJCJ4G6FZe/uS3WZN0/DNWQ2h/Y+kPjU/K/tnKGLFuDeYLwogrAhKLPFW8zc
ectv4J7bKZi0U/JCNxrIQiyWsvnSmO0Qc2L1/A4eHFaHhIzUs5ATRAGGkjvEAgto
2NuYsLVsDnnYBvrrizyICSbkcZTUpGFJvhmjKZevKMtdVZTsXyBvdhCurj7GbSlJ
QSNsVL/lS2T89/o4U4EvMj22147Ij8BcX2P7d8iy+83ro4EmpCR7nVWh/izu4ZWm
KsKbEJI+DkGu5TOm2xhgJugVB2Kk4FB1wry4caN7+TsFCLPQn4dK7F9tIDDe039a
CzaRusVxUmvJzo0DDHjfOzaZhWB7mcZiMNCbQdYIUbZvksQgL11QV7er4/jp/O3y
vXotT06eVuJ0v91a5yNUFyuOfUl4dwGH8vEAz8GW73kAZUu+pMuwn40G1HkyYynf
42R5t+jLasI3QLOQl1CCcIKJJ8r0lLW7UXEQ0GemKQqWaSuB3nqiIsExYbtCxj9y
pTd05dFaMQEo+j5emuODe08BU8SrIgGxcju9SlHHrfZ57Tx3a1ceyMrZhZk8JFNG
cNtY4Xro92zZwKn76rLZEkdrl0/AYrVUZadec7vLKAi/eNYkudIkTrfIwTPcMi1P
O/bZR/0j2HD2C5GRQLpVkrHHsY+ptwK0k3TdQke4MAdQ3B/8a782L8QVtpsv738D
B5edwIUtDkax22GSERPl2/MgM6hUxc0hIKrE98PM3EL5kPcSbCqy0/u5eWwF8RHU
udqDfrcTDy/Dfl7DUIdTwDdyKlI38yeyTIYT79uHw07fa7luxYcmYX9I1lW5Cnv/
Ycnok93qQuEH8tevbLOE2vflJEiYBbExOq+uEw0jd+8FYxdfn87xOkwAE3FFjNRu
Xn8vidWWgyroz8z0DJmbRFhKPWL3o6iOUSyxkWotqLea/UJ8Sg3OHAkYMtV1MzcB
obf4h2J4usMqLTAHHgiGD7TAKVPi3TcFzPvsa8jGdOOKZKYPidq1kZCiG1kffI3K
pvXl7yfZlz3aJ2+2vZaG9yg07JuKhTSqTaLYj0YMD0WdmvSkwNay2DQFepHyF+5k
N9IkFFr5/ezEKro/AhSshMyOdxOH6cYZBvDr3PKpiYOHGlDPQMtlGb2C8v3PjQA4
ozJXCSf2z7bciQ7KXT37lKstS2o7Ep7slmt+d/UuaTJyXkdaIYGxC5y2UYeOzT2v
0c6F8z7g9LzCU9WxGd0lxBORPu6SFisXfT2Upxy2emdAinADjMjKdH1XpxJt3gRZ
Kc7OpZrH4GI/uzqN5/jCy8q6BpR9kelFna7fDUf2bJNgieMbeBsbam4LjqHnrVHC
le3rsPhKQn23iBRzkIqqBQOyq31rt9S9XNU8XWpXSAyekFNETnMJjc2y27JP4O/T
klmUgVaKKCh+bsuEwAcQz1gSBjOtrXyX5XBWeYPsgYIboxYdvrGTW6LVw5XZpkIP
Mmgsu1tjusg+ChwB8eV1kpLXkUCMMU5GkOKIqb6ErpLr4HlvoIk6uvMnvVkthyFk
9X2i8df18GXPO1je+Ndh06vQuellc6PnZKxP7D8U+G00jo85tKpk5KE9w7fEs///
9TUHYkqJnIz70WHI/2Vzs4VCyoUXE9/rHWyJwRWQjGQ7JEUVrt16cXSL3VR5BWxT
+1EBHKlqGU3kdFRf2cMqq3lV5IjHarzOTGkXTT7sp5peYfWnveMCFarQpJCdViOd
SgBVwxT9Hso4k9u4cdn5PyYihz38hnVBVlhbsuucS149HlrMQ7tl40fKovcOKLNT
U23pmalizng/bg/GNF9pyDWacncSGwVSXain/kEFgbUZqwB8mcVnwXno0iAwUvVM
HUskeIXABC+CiW8LmFDF9DCR2QzBmHYo1V5LwVX5jGzkT9/67IAENfWhmLjcRh0/
8iXhbuSlPEchzhxaoLJrR2c+IH+Gcw9ERd2dIOddoq7pyW+uZCKuLqwTthHi4oSF
nXgvV8RwlQEAT1nWU/ZwEfjvPQHw0kvrLE5nNh26NadqJoHDEvs7sq/fOwwjBA+3
UnH2G8Zfo7fUHC8U6uGVCal1znhGQF5KrV/14OCv5J6nAhHAFOd2jpX2B2WFbx96
P04e0XAuXn8YYRcWP2AwYL9YC30zmr3QlzwUCUFiFJdlnurs1ClycwkgCrWOA9Qs
7aV3qS7+qGppvyIcTpb0jSXL37WoBcmHMqIzrXaNNEAZvx1DdYySi8sxf6n+9F64
hTlaS+rDBCTN4/tEk6fK9/Rc5miGL2gftG5cPzC3o2D4LiyWxZQEA9a+XctEDhku
kplav8aH1/uW43RDDjwm+L4mC2L3QYokn/c6UWNlQzo3BwNO6x5/dCEMGXHwuOZR
OFuWfqqeKRwrJNMmAJ51v9TFv29LavGFX1sZ7ybOdAN3rJRalTXltWERSe4EIURY
RZBzCI281EI8KfRdCHqqQrGaulMnLgRemiZ1qJSeCwx08zG1sDGx6TVwF60CJ0lS
7yx+1wLd+uTrP3GjKS44zr3A+r+v0dkWpVIlaRg6wsrt2HAwgXSzhW7A4YMFPkVB
LmPRf4KVipx76E4WqhwfV9GC19ziCneG7zp5ozc5v3ShgCQC/Ni94yFETR3rUoV/
ofWHzOC1TJPmunPKXTwp9bFwulzvo21SZYsMFqVZF+lC2Z9oWwWkjijTllvR208y
hPHwPctKAqhsrIlOaDRSqqNBEpFNJX/DJrKvyMrRW45x08ouoiuJrtpR1kp5B3Qt
JLz6fUpQ2SPc2gebP7ExiFpsuiwRgfvqzwnwcfLv+P8ccOxRMCJmM5yrYC4xgW9X
UlZiynH1SKzfosklD/XLgE3SPmjSQbjHpEUIdOmIY6gw8t5wonfwbGVerh9F0KxZ
3oX383iykVkgvFTgumxY4cCJXA+xabxW70QWoh8pX7EUfqYw5pQFtDpFZhs8odCU
O9au9F+jiwFEJrvKpTNs0zp/3O43qi4fwisULzYR/j3tJ6V1gjKsxeqnj9bc6Sc7
Zazqgg4Z6lMzzmirfu6QgTF2FSp6qqklxHLvg8q1Ll7R1qxQgn9VTSdXEuWvwn3c
hw/FFXTG8ffSz4SZpLkT4U5URi1M9+DkG4MC3ww7K/F5dhlhlkvcCcYLyhiHqw5t
scUe+/5VcXL8EOZ3bskOxnn0BIikcYzuwXcXXbHW6WYd27bMGngEnPYN7WlpHNnE
+gK1f33NeUYQJm2qmwf2/p2UrYLRJS154zlaW440+1BFwHRC57/ViLM3i4KGEHU8
R98mB2zlfuJIypIjiog69ylGsb+VGl8sJZ0wjza2u36OtouwfT9s7MFvhbpMa9kq
B56o3VjoV+jFQxgt6tI615eSfQw9pc2N7EwBC50hXPBI8+bQ+XTxFrFUOrDQ0pKi
/2h45ENUiqClvyqJQxH9q+Sw4qslNBDNP5CKrHSy7/8vgMs6QpRw3g4YBqcXx773
ELTqi5iDcy54ZJcVVa+q1JGP79F2BGUx2boFv/bRh/L549E/VvIokp+Zzfej0KNs
Ona5hjaTsKNtXW8fph0O1P92Cx2V46wBHAYkuCOSJTUsgHU2VldlQIymYLoqS4RD
YAthxn9WWKDPkJoUMHtQuYqyrONaGIf6/+wkPb/iXVFWPY1Yhc57SE6s8LxcRU5/
yG9DM/02MCmQCpf8J8rQj0Xml3WOi09iXTpkjonljo1+HW1ysKNOVAagOktAPSvE
mSnwwjUQFtehvNrnhhtVLbk9aSOLC8uR1hVkRijo/CkJ9/6vFao1z2Ct1ZZ+DfX+
0z/aA3wbxJ2cTbf9EiRKO5ErsGxdOt7yV/42bUqD/cI1G9b8JRCZ1XC2IRhRg4cY
yhbYQyGCF1ANg7eWtjnoZuNdpa9AwhjaWVr7hRgyppxeIX/rYvJtvjGPnZmMjiO4
SYSy0vYFgB2zChnfDPcRFL+2b2rea5U61AbA5O59j5qBanksArlRpui4+XNEBjYX
JcrlZ6pe33CBPeUMPyo2X/CItvWtKaKDdNeOfikdVdPvK94k5AuHfUSmzMq42qFm
GqYdz0evKoOYVPgQYPGnwf6G7jVoboRGJj/6h3AhFpP3TUpmT4qeA1cifw4usEy2
s15bzdaqkXbQgrTNxypzP80rBZYlHdTnxVU0kuxOBOi3wxz5Qt9kc28Qbz18rrjg
4PXgBNpAMnScUwmOdM1ys1LhHSqdJLr+yYRYBzLgcJO+hPuCzfxGZCEaF6KPhk/z
G7g0r5wpXPNBrGzL3OoP3ze68E3raS9nwHUtISQf+BhKpacw3hf1NaVz5OmX5WON
48J1iJGP9AF4ClCnQX8mllrwSzRvDbmYwNWYlnF0+Yim4G/7MRqyPzRArZyEZYkw
kAv2JvkuR/HgH8Hzl8CB08KDr+tW6XTXCYFuMSAYuaMJJGJXyF2sheoa7ZEK7mgD
fGp9KcZx9GD8k0/AADjNmdKwH0qj7aLKqSOqK7GhJIyDQ9Diba4vohLEjxYrJvlq
oMU74+Oe6oiEWqoxxYYxWt00tRR7zx6FbWdy1SD0NnYrAmU78VuJM7O/ryJQcRLO
pwLNJfqrXdJtBDlC+Xcec+rfrq10bzEgEAAP9pWnuhnbaz2i4wQCczyB5E1t89Qu
lwvGiDLo59p65o7vY6oWngwNrkzR1KD8LGagHu+Jt7zbnRM8fn570IPAO3ubPWBy
tuF11pT9k1vn/o0DRN21Aw/1DgsfyOCdrlsluPbX2GbUuHijifL9zPVPnFXayus0
SiiJXt8SyXaBmKcjRU31a09tQH5Kl64InSQTAYkc2ENZQGcJ75GvkhbLNIiupc24
NyOJOwgs8j5y/ELlStoc1D8JxMXZq2ZSZ6tV9zWf3SEsn6AA+W312gpAx3oxGPrj
x6WfjmxpH1EbEpQ4f24z0l21RIjmiseScOqly9YR915Qj8muK5dwi96q5vz27Jd8
7Ln2q13hBW7eEcSJUFJbAzMf91oGPjGgNtH5YKveWV6KOhGVRaxrqDJkRIKYHzQz
9amYrp8V5684xhph0Vkx9hSH7CDtNXGS+xnCWn4tM5+IU5jsEr1hS4o+eCf0/LHN
Ca70PiIs7peIWipIDmzUodz4OiPduIF6Pr3iFSLc6HmZYJbALfEKwBJimKMK82Wh
mtW0qiibukO7BsVphFz0drKwZzl6MAlB67hloIpOLhnYBtOlk82HEb1XiPx9frrM
wF2/zpDjTN56UnVtVK29CmLCTYOQ4ZoyoQLpgk1iwrYT7YcxmiD7yRNHxKs5G3C3
ViqRxlO2rl1dLR6gbkowRrggiy+0vMMUg3/3pshHm98cjxbJhhzz8UUj5dI3AKRh
tqaSRruQ8S6i51aecEEaIefmmH1PMeQ/EjmD+HLB2N/UwevmjME2G8ondMh/wdbB
14mf0wWz3OFD+6+Kd3D1GHK1frPFvexHK7MF9ukv7H+fKbZw8BcNJ8MeEaaqoM4S
34kqosVVVUPVPLB/w0QoDkIOiWyUP0ySvfIsRhWuE6Rc+E+uMGoc4UxMqCVbvBOb
vPp9P09C3B5h3zMGjs3KESC59MPUbuuIqiyOnpStOzJQvpDGJaMh6TkZ/8Pkrd/1
gwAHjHWDinQ104+ScnkyAhN8NSDiZ1fitPhbo4C3h1ifWoyqrTfl62g00UmXJS43
mlocw70rFVlOiQIT7+KueGVe/ALeWazQqb4UIOP+mxR0LijLcDrk3aBynWXb8o8Q
FkLKuxULpTXV2UVFDILmFVjeR/18AVAcJ0+APUmZP1CoEKl3yFLfDSCPcnRykIv2
Y50AGpx2ZSXolt9pa3ZGuV7EasX2JusRhR392cVCkLzmKkBRnI3ccve2BCIs6NCS
9F+KDB8/nHWMtxOdF0xCP/7XYynpcE0uaK/s1Z/caSJY046XxKGM210A2NykKjsC
cS0jURGjhBvg/dceuFSoVYZ2VfPTs4q+z18JliFSfQx+KghtXMYA3l1XnWjmKT19
nN9VrZkTxVHYDhTgAoE3ojdD4Cccn+WwfEBgvNjOh25W68TlzAwjePENE8Rwp93E
tZ28Jdk9PE+OAf1R1/KrjnteZ2ng3N2I9poDsKhhCx8cmX7MQCOAZy6INNT9Cofc
ijLy388uLIJd4IrFKE2vG2xmnDCtIeY4itUs1AlQD25bNL6V15Cjij8fABEMOkBv
Vrds/snXfi9eBGpwGIw/gOYKdfb+o6yqyzd1sViVVD8k3y1TxW+1tWZQXZ8eB1b2
zab4IqxEPnEHdVdNZjwZCdgB/jUmvgzgHaPH3CnznDl64ScqATMKJ2saZB7bBgVz
ffp6evlLObsuKrxtBLMAahrq5OLdKE2lLW0QSaBL47/dXJc0XCVhlQ52dAtgCfId
k3DH8ya0HxGOGAx8/9wK5o7hCYxO1qhIkyXxfxsfzB0zmr2T2egFpmEBZMt9SuwN
Gzqzglkq1hyR3mEeJPj3ZJuXIRbjv6dWFzZ8t4T4ywO6CPCOY5dg9sqrl5gO4rIe
DmCxSZ0f+i2QXUQiwm+NvywAA8E2vCRbDHANGTjVvawPewxWBgKH6ziqF5r3/jk5
DJjJ2YRO+SY4rSAMg5Dwvq1yyEUKKzzzFTrtJTYzQgZ5Rw2BTClf35dwzx7cPKD8
yx8ihAz9Xqas0WgFP5ekN02kOoX+QIX46PhZigOUz0xitug1oNSZmrQo6JBc+POQ
cJLg7e0/5UXAHpl8VjQnWB46avgCzNqngNbMUxfm/He50IJrx1fnytAnuEsPU1zp
cAYA0qDfiomfI9+m+bE9OF8OiurXJe0sAWIBC7Z1XtvxJtH3WhhtJjjTS+FGFMG7
O3O1vRG7dQrFkOwm9Ria0lawWJZYcaR4nmpgTdDyaCQpdl3TYkwnk8slJwTD822h
fgXSkNvX4oi/miFSuNNapfPIG3S3ArhPvhcc9K3MMMm3Sxo3M/nUMddwCLs+qSqt
UmyMKyu5nE17GeKKRgze+tGY0cQTqljCZEep3Zl9c63ozx6qUJFXIRGM71fFimLV
Qrm6+c9CZNuhGHI0o8aCAp1m514VHPa8cuuhnRCpPrJiJ8K+yo41Rw728yq1zeHV
COqiLZyMrFPDNecqaQai9QUY+AVpiEdpXTIGsD9h716RRbRWEsOLb1UIxi+o8QaN
oM68O9Lc2sRxtOByFhgXE1AyldgZrKkgu1/+RNEd/YwgjbEAgpWwtVGGF9VlZv66
ixNoxtnE8YQAeDDZsmzmHSP61fBODTBtjMMrAQk70+a2O3w4aBTTi+WUEOw9t+U6
HgbdRSBcQVKoMfvG5nucWvYdrObrk8pZ264CzDK8gZ7ZB5iKqB9XN3PFowMopsNS
Yd52z/Z3eBYLc4u060WBy4x4/P8KXrbmB1oI/Uawh5Rr7wJYTvM3Dcn5WfpeSGsM
T2aNrun8GYByhczqCvx5oirSwGjld8AzcKshv7s+elze1B06ote6lbXMNPClBNko
XdtHRNcf7L8ZkiO0uYOCN1CDM8r7bm1atsDmYru0YXky8tG5djcJcp0KECPmC+BP
nz4bFvMx2v81WM0kuWIaUPBmV5mQeorfWSSSGLzZtSUslV85euUzdvG82ZQ37gb0
OeVoattIwcZKRMCt05NbcpkFCKtKDFr0gKcV1mSZKf7ru7If1IvCFICtkUuyTnbB
OQ8+nziPVgSZRMDM0nd0zx/Up/73PczUS3r333lkGavq3prt3ZbR2InC/ZPzxqm7
JRduZN+KxdVVWFZZOMZZiaIgHAqChD9TqOe0aRGhpF6+MTxqmW92epLUMggi4w3p
WExySTNE3QTNwpsdpJxXIuxjYJXBRP8j1axTsFoaDu0VkFRqqH98GSZUWgfv6vXs
qdies0UFyKTJ3y5z46eNrgbPXC9xGw+F/4piIp6i8T9iGtfiFIkuWJfHby9Cob+/
H52tCO+8b39n/xru0XFbydLplaZ58lxS+/kXZGAqBYtbbM6DmxsIIhWYUTmOgbJj
3DgZi7mOeAq1QcVHTIacLxCFW7HBoUrpYo+QkvQ+kQzenjGFSsVfHNSkem/N3NML
gUvhWtQebH2NXW5VZQH3hdlKc8rlhR1Drzakr2CtQjYBZC5D9Ll2AdP//cPSoycB
aZSgesG6xItNIqbVGr88ZSgUler5GuXfomSIWbWuT04RHYK9bqgFoh52gXylEdgk
HtDJUJFXha9jLPk1Ai1sYym80K6KJ3O5PMhfeFTyE4G4LgI01DkQCn09XgiPbB/C
Ww4eToyOYW2R4dDM2MduGpOIyyH9eBMBkeLkPIRcZWbyvXHf24/xy93811+WvcCf
xcZ0uPl29Mg4ovPXRlV5AAfOryfKnErqEX3H/OPk5MnN16vTNH5eYf0TxpRyb0nk
+NbO7yu6UMbtAxWfaIA1qpPOmubHJ5wm/JU9cgTugW38Kc/QPkaNGiXHx4vkPmm1
XUFvqfDgIBMJ1IJiZ2D/MoxSleR2SDedeUuvRTs9MM5iZct97m615ro1xW8Zc9VN
3HG2j/rfzUQduTvxQHjbYkCPWbDA0mzL/SmJcVqjLPMwacpigu9h9IVDKKERTvUD
BnxyR8p/DzH1Ly8iy+2pBJNViFuV15jKVqgpV5C1JvYSzFJ62Fl/MTzG87ho8Y6w
B0LECzkhJi11mjAqS3dl5YI/kTg/tRnWNmVj2QkVvXE+vYbW1fUbpLj1H5nCIwdK
n4KhEOKhc9lW/MUmKiodVYwZUuBj0oUo7LIEAO4YJs4s30a8iF+4GstoiH0Q3dU2
LiL1Ov0nyolzFGNdYSViKZ2pY5TZYNOzDjhfDeq7/a8piVPVW8BXesL64nDRB2qb
f5sgXeZUSFZaVJwS6R/tfhdY+FsaxcmeTAFdxFGSwnIzPTlTzAnLFri5EK0swVOR
MBW0AD7+lG2OsXOdR9/azUP04c3KYB3KNKrY4E08774yajbmCP634vOl+aisZvch
uaFCG6btQ2W+zFewD1ePLyLTEPQK3U2Iwgfa6meC7zxbQOQ7gTIewINs+jjkuK25
X4nXajkfinFVvOVOAZla7dStG2RUY1AjLs2rMKdp+bd8Sx0fgjvHHShcBhtqjQkj
mNQ69FGjQpaNarrVDlqSP9EocHynlfLzRmPdXmKxCeTxpD3phkiFiCf6jlLEx6Hf
y1qprTRYCINDyE7E3K1YHT9Z77bud/kj0NvAU0glDVOI2YylC/tagBuKHhptgwpI
AJvugmSpaG5etl33yfb28Kgd3XePlzXbNByYS3qQE8TWUo8Ej/Z5EYe6Cxa/rqq4
WtxJgXSb3kkZA1Nng7I9LNochz/4sBf1w3cm6U4e99/xkjVr+V1dHekVf1lYR+0N
3f0mx3Ol7crbajI1pEqVtV+qGYUdo5SGCp+ervkaV/xslTQa2QAX0W7VfIIRKkDx
EfCcG8AVM8FgcwIPGpq6ND/MIOASAnGFxHtLOquhoJRJFpDD3TTxi3qnl0feTzhO
5aAFebOjRkEF8V4NOEhlfDf94xApcqUuqinOXBuTzc5kWkhQWtM3Eo7L+z3FMeXy
9QzPbqduLF0ZOutFYIZjeYXFL11FalVz8y1dTM13cuoNkxTvsgi1zBJRkRZ8Artr
1yK5xieU0mimvgZ/9y0+C6nE/xw6cBGo5fz0dK4nE5mpGnqZiY7BS9lwQ8cYn7dw
6i5Zvv36ysWcRhgFOPIZs6PCNw1PvXBNy2lgSQynK2ZACyqsisnNDKPB39sDAZNm
j24M0jBz7eUUu+KR+RbwSnuSOJTps4oicOV0m6lQJarFJVVsuzD+JfjsHJNgC2gF
6Q/olP0Pz9jdJtxVfyMUCRcwJ75+lfX4R1vEnLopue1nzp0k44+lh2a/5CdWXpnK
8NKPn9wZEDcOiuncr0XQAFJ4hQXeg2tqlxwJ73+gm1gZ3dJC6TisTFIurKpEDlFG
Sw040ktb3u+QCkLMpGxpcL/kIDh10Za/qr4mK1sj1p6xAFf1ieVgvJomH4ReU0vJ
3TXh+M2tZrUKRyoXhf3JzyaDjuLlYIynq9uQ1kQu4GEI7rviawalCTw+h/Jr2uTU
2fTHHK2hOQS/RgwaBTq1leqh8nJEJvUEzf5iPOol9Old2C9+UkkJfZcFT4UsTNnv
Rvo0lAG1xQAPOLSxRskvPa+KXd5L6/BWmMBdf4mUVbkmWnL+PWrXke2+MD0dCQIH
r2L6Dcz7kzAdkOQRoqmgtfyFmmY1gN1Q7znYcVmUsrPK5bmmoWilW5+7culvHfj7
3LaTKJ5dgA6aozpmzi7QwWkHwsy8yHlJRESkHXca8roOcbPpHJn+ekVsAFtxxH0O
Y44op70wUpLL+QGmOADctae/Bn2hIpzDQfjNjkhOLwYYjIAqmiQtSKa8TTe7b25U
Nomcctb8Owo2eJ7fSMTZtzkFG7MQoyJhdzsShmeoOUfclT4KQQr/k8XaPwMoER1s
l5MoHAQ4TqYWGXYgK0R7sG3PpnpQHedYUKfmPVRFBjIxmUrNoTtNC2/qNaiglBRf
LT2fbOsRro8YtlP13P7rdcEuV6Mdnb8H2/GvugIuKb9iifHl/r/d5OXq4pLQUCp4
rkC/xO4y8fI+q2K+oLLWZ/OmnSolZtG/zcbtoKiSDSb4WG1C+imq32dgd9Cy6VgP
ndJmfi6J7nPN9QSHujJCLjfYM+6u1LHpi8S/j0GVP2OfvBZs6ufodbbpcOM+obte
4E/pMEXngqfs7Y17qEJtETRtDmZGJR2cBMxB8VtlBcQJZvC7CwY/CPCQCWWiBwTv
EKS/tXqSNRedkOTykMOromHj0vpOIGpNnaH3mZYVrhbr4XAiX8840Ed55k9qVW0f
LjvaRb/8Rh32L9WWK/sEhcB77W/21VlJjAWyrvfxKx6Ksa6YBp55PHyp9E7mGRJI
CDfJ9akcNb5mGhGk3kt6xOeEPsD2W1mzNmk3Bwid7Ar71rRxyflYRGHHx12BJalM
opyfVUlIiaopRty7oH4STXdpXoExfBWb2KTSZ6fPPAvK7sRhDWhtM1IjmNBa+D4K
sKL2T8PbNG38hTS9ZV0IJLerPLONgj8APYi1H9z59NhZXEKjWFDepMI/5ok+woSi
29Xq0MLwPpwUNeYfZSN45+iqHLzCvbmukFX3G6pRB1tsJ9oQHNP6xjg5I6e1EpDV
lns03jaBiBEJyg+8QyJQUjRg3zNhrfrKgeJoz4R9PKbgqpZfziTEkAsPObfvr4OB
JVb/T7jOdbUS97399J5r3LdNotspx5Bj8aEv6tQkGrFrlwuPnLGqKKpq9VNJHHwi
R+M5doCBoFEf6T/+I/Z+QVl8DpX6Mp4dsfXym19R1e/1+UXI4lthfuxsyJiAU97D
Ke2C6m1iyptuw1Mi+bBomMQr+OlTlO2SpFmdr0b4f/SBGxQJ3kimgaXVONIXEvCr
KjMb2NiyvOWKzjJOakKSegMJt4MfkK3xnejH3CCKvJeqLasMT7y5ARkgOsnblO/O
IOD5yaKYcNc6uHoBu8tYJqgcWw3l0ZnzPz2gD4yF5Y/uPos7dT5o1PwgJ8q4qqgq
Lzwgv1fFlhl6sP+fYgDnxsiNQlLH8E/Y/DTS8pyHFIkK/SvTLMmrVdsdoYaL1JkA
V0cfzOcKZ0rh8bqAo9oMVDYM+cz0uCypss5kCCz4R6KjiGRlewFlvqojoNJ79fLb
7jndoBN+IuUyBDCsA5CYTgSUY1bakRNvhs4NiNg6KBDN9WW6ZvZLmAHvHG55KV1z
7I7QL1Ex5KLy+Agz0hutH95o9NEzFNvlC9sH1StkflGzkRv/KMJtepV/yvspx013
3lx5POMcHidvQCHrGXPzm/8GAyatJjp4c7RmDOi39OWrEEbiQ3fkPKAYfpofoYra
1imAEmsJykCJHjayXmv5Tpq2sDvyoytCGS9gisxTGFpqDyY2N2CxZrB1qEUkWAQq
B8vAzNbMxKC+CC49mTKmN+oFJLlVCBAkDkj/GUZ1296rPLVZxPivpEPWqhQDXDXG
wY20TVxqZZO59uSApfmAOjWXmz1yGQsYEmnOWcWXpZiYy4rS60ThigoDn12a6V/d
3FXDbR6PnYayahKs0Jp9b0+EtkJaoLacGOkXLc2uMK36mi+7bvQgpPCqH0L0plTf
JrleqqQWY8wPcQG5wiDYqWeQ1pXflQ/w76gkZ4zZ64+m58bSxxcMtL+uq5a+BTEY
NLe3LqY7CFbGojDzTjtaFltq9VXrnVPX00S+O/Rd8eMWr/IIPLjtBwzKu2SqU00g
a8dwC47j7N/9RGioQTmT1YvajZD/6K7JdB2fGyweb3gP610hqCMddbJtIBrUnSVj
c5TrADRxuLiB1EX+nnwnajaumNXIXVnbydoac24l+ut8OVdmQpicE8fD4lTKlQKV
q8kzHVlWibGHZdHZUq5OkvCRbMHvlW0RhqpO5S4aV53GEAwYmaKy6+lv7NTd12wK
bHp35VTArne4Vu5TmqHcRRH/VEC7bktN9xTa4WhBHcsgyn++J0uMVdzFlWtFoX45
KHsb+y2ebhgoDMdc5rRBlKxZc7YT35xGj/okB9rJnMSsiRZrX3o2achyYKP/LvJh
Q9xPf8EL79XYFd7T1kuF5COgB2hyOITZbTPfPzfScP/TshbiltBrnBCFlg82VbDR
vDLvp9a1WJjuVTWcsGmOLrNvlYy4JBeqZQnhABJ4ifFBcLjYxsHSIXKK+MIPIhGh
oZhV0ZvL9v/4b8qm1m7ZAj24PC4fbWHNrM1Mbl4Jvb66AuFMGdHpEo6EWnUChwVk
4d9daX2lQadC2Ar28Mja67xuMyot1GPjd6SGRiwiFptvDENDefTT3y6t8vW389dp
soImztD/vZ0QVvHqec6nN/KdMonJr+0rdSBP7eU+iBvPKHdpDzapHXT1lOGbrZss
RAchn7FznJoayv+A3gb/HdPMX+/TLJRFs3qZbkQsG+tMx8OLIZ0aBNMihJFeXDGz
CYPHL9psgwEVo6CFM0CleiDUU+6uLMPEo/+jPkleKVWxn9Ni/letjNW06x/Cn9WO
MWyZdWRo+1kD9GFDbhZ0Rj5ms3jXCbM1I9s1484kBW+QjLvreRUy9TuJBScorZYB
SLXpwbtjbcCn1bkW6R2V1RiTTj+nlE7gGeZD6GITuFV4Il1TEqk3f8Q+72sdi3dC
9/vwESQolZtdjiOMwzv6awpQfGxhGTFVWyRr7dl61ZYBnCFMrSWn7HYz9ag5eJaU
NK6Od0IHejaa+p6oFHKYQiR2UeTbMNzeAFY2agwk0TIX42Gc5U5e/Q5ZhHoHoApX
BnvhpdhbGdMaKIFhEMX6RPTJ2cbUUi/qq+3Nnvl4lvXyFDNx76+PR1n41ibZancp
LgmMUSFp//IZ/X5Z5FaadAA9u6YWGY15iE7+4AtIYFztiV+t+6fiDY+htPrauBBu
Bula5C7rxLMf9UQ8ohnWXP3m0hHtE6eE4w4/35dwI7Lp+UQ/jE/NIkr3TRWwCVFL
/l7jkqudIpr+6jhN31Sk7QX0oIpbWH/tdMhbmN5ZQ91b49eos9DH0yoPOviDUnCv
m/OIKGpQpBcqn0ycsB75xGFHzxwG1+5fak9CUjqJSjlGyZC5knC05MlufMUZG2l3
OBJWo+DFcXoxWpzDTzvgjoeOEJOMJsYl1/hKBYCVAOi3CNRRi+o3fnbmR+Z5uwPL
tKQhPtN8gnoCbagEJCMgJ5RySIcz+pkqEYBS9RjsnAMIZYKxkNe09xnCoo/O14dx
/KpSLVDdp0RzZB6SAYTeeRjd0q5JeZwsvggMD0Yjx0r1jKKon2EXnK4BC5PifmUq
2WoWtoohz+DVQ489iI8twIid2jbD+o+6fHf0EcTFbWahx/FeMjuEUrWHs9VIH1Pd
GEoBDrUs5w4AvePGFjDm3NRPnEeQwgU7f41oYNmmmnJ+yiTp4U03NB+K5cODPF2A
5C8br4rMjiOh0mtmxQNifLk7l/6ppBCa7wB+ITd+yZw0cMWW8qrqHV2dmM3Ss2OX
vS+FlESRdkQT6WErQVaq7ueKEbaWyXLTbhGZfeDEya18KZcWqeg6zdQp+xz2vIKm
sHMWzQ5tYVbyKfl25yyxqPMpDqrzJ4q2bDW9Llz7+6B5qz3JTieMUGHgNP2aMsJt
jjbK+0eBKZ5oCYqOtfsDHEmXkhaah04lUkY1Iy1vbqHcjSwRHgC78NgyaslhhZg/
o0Qh7vMJYEpWB4XcakGoxSyUuJclkxAWzYatOi5JUvI7u3urxJib14MZrvIUK+xZ
8IQ5Pc8hWDVXCidiNc8TpxnDlhBKvDUJuhmy3PE0JjCBna073fNzPf7u0G3oXKrm
z45fTDYj2XqXx54oQTWN75ze10Ee5EFFDK592Fx67W+9fSlO/rZzFYb0cI4tRDKA
MwqbofBXX5vsWUz34XKaX73w6jzvpPG7kUTIWiSe4sfpoeaU4ypR0HufoocBrE/d
z0rkpM7huWQB5nq/AHZlpOCLf4eSBPoumfpF6SGB+0Ei29zbwXySTS1duijdI1Z9
F/jiHaXQmYXPIs0UQevbIxicIzNCPHeYLDSZcpzTAKwC88cWRRzJwIZUeSwA2LBl
Wjvly7NB5PjzHiKPgUDuIfTrvHf9x2xus1pFsEgdW9diUarVTWp9TKtnvRdNO0i0
b57r+2UNitkk38U+skBTojU3hp2IQrfdSkR7IQVDczMYq06trdAjdUikM2l8mLLZ
7VlQftlRW7lTFGMTabLYTcL/YM1XRJV1skbvywNYw5m8lvEQeE4mDgnkHcktlMlz
JsL0T+3eD9AbXzQGJVLspcNmQSFrDuWXKsQ0eq5W58topc08giboiUTUKMESN84w
ob/y3Zv1b3mp3XjpsMm4sFW2ST5JwQhrC/DjNFow8ViDoAswJULXXd6GgXHbpcjh
rB2cOlN34us1zq6L6UF3x1rirlMocUvCUMfgSnZWZXVBKZ8ipGiwLB52MwEaQpii
pKGJ59U4ACs5l3oXaoqLHLhnHZwOrNP6NxL/AJN4qTPxQHcncenEze61tGZ7CUvo
vQTiJTdPLBNfllrYHrtMSuCDzW56bWywAGNSFCCCcMziT4RNi5tj5LIMQ495Y4qL
dJmH8gX7E14vRYM3FhOdiipS/lUgXBnD2SPmecTfNmEpPDhtnp5ZXDkjGWNIEnLA
IrXqEVF/Dlkt1OGVJWNfhoPn9WBHIy+kgXqye99rpdMFkQLRD4ykeFKOlxpJTX7p
unGfV/Gv6SIdlk2JDcnL/iyFNikzpZeC8PhDI97i7jGd0eI7MGSGtzQdOWrYNo97
MFqMnxDkhx/HC8KovUA0ZFjTWR+LormRCLL/uD9Ilwj2QHZxLqz/UfpRepIOtlkg
2aRCk5t18oVmlqFkl+17b9vRFgmULkT8NQPbEzomNy8koeJW6n7hr4WPS46Ay0dF
qujh5dimof6t0LicmoPTDvXXkctKsF/uH+KGsqpc+Q+LHc7o+K2+mQ/MTCmEkqSp
EeA3OdaXzISfAb1pdFrKJtO652JlmoT2XOC2NUyb51sU0uMk62YOLdlg7XUd3yi5
TgFMXbX4INnqj0dMgu6qOrxoOzg6zFp5SsJfNm1aMqJyUNbb/ZiQXX1yCrMh1LPt
ZvJo82Hk2Z5f6S//T+1AjhRqbzPhUF6/tzIbieEm6p4Rg2VFZOKiFHZ/UlkgXInQ
R/pQmNpOaADKBOq5T40qGWYTxrqxgTy7EQmu+3G1wW9RTJjAAI+pMg+wfjoN2Hza
7JxCikd5ui7/0FmjFwENxpDRxuwh1y9Kail+7QpSnN+YTVuI1ZBnf2G/1d+SPER7
N6Bzr3cbpON18x3tYzfhLy/eGSZNhnxpcAtEtw+EQKRizek4/rpibIZfbg7SEEVG
yFskj46NFDeaOV6HxU5Bx9n77z/mNH3/y9gbOfsbPDQrQ8FtfjmxSwvoIaMVmUaa
OyFAtCg0RHSGHtkcKThWsHVccpcxLhlsS3VuvSlttCmTR5U1HRl6pCGFRy/FNvEN
rbxD7Nfswk6UqPWP3Nz4ghrsJTXbeWciSvVs+FfVs9GMuox5jWMjyi2xloFRCRIv
imTMeozr8gNVZS33kS+zJPm1Bz+DE8bnFcNesKQEeUMYdmyRhayFmJVyi9nuxRR3
SNmHipKSHGRRlA4eSpotHHhNQtZ9vMHMEq20biL7meOPPwdR/19JvmNJ+NT5HGuF
JGjkdWDsRolvsSetQPv6cgxFJNVaXxx1knIgvmm+YaAp7vgntOShaeCPOyUZRcyc
WeLy9cgDwnbSNtBZtcRzGba5l5nUzcfCA+xbYYa8Vj10gk1JXKBQ4NEawnuC29l6
mesz72iZ7qevjF9DSgvrpnq8xFFcqf9QGPylEEgsU/Epl4oYwPyJyRzkhS/+PSjk
S77yzrzVm+VzswBLAod5CtjzlWX5YpNNy6QmzpD1JR4Wk16HMdIxtOU2oQHbftje
W7c3lO8W/SAMJUHiveIu0c2iB73yDPQMfYUw8Ve391Yj22gkWGZQEQDhiK0jHdU+
f3LO3DsMQ0ibBNxe/QdO/yfXA3r0zX0i2kdmai/EOortEE5LE6TNzFz9+aeM86lG
CRGk25r0wHeoexvZcmtl8HGrb42GFFPveygVf+CBJ1OHzMngA5U7OQ5KfhhNyQns
DH3f1SY7ukCSIpD/6oC42Cg9wB8Xo1O1rnzgENHcPW+iFG9KgoLI+Dej1oSgw2cF
euypaJ7MwoDp3XKuJ4lD8zMWJXNjv92KZgHZp7cWBN/O3gq8hALARo+g85uoKuXT
s4Nva+mIwgH/F+7hiM01NHO+zInuSpRQ+e6sUiMy2yozCjCa52d1VPwBqIqXL8ZN
S2Je8yEZHJ9OpFGoA4RY8s5rE4HS/Gg9OuPP4w7hnPw8R0tSGqzBwB+9Lg3DTK9+
mWUBlsosLkuBT+lhF/aQByDOxU0AjLgEMmUG57xAwy+fl31W5SWg9/8FisyBjeho
1sSfM2ljs28gl5HFsqITB+DaC6EOLE0ohjYF48KukmqIzs7yPAIwc2CV1pEP/Ns7
0IsX6ubtdfGoJ5ZQ67SoOtuEtqXrRwc0mg/lpnRJsX+DPyH7MxnNqr05p9VVSdFK
Hwlndrnf5rNno2O3vB6vtnuwtNG2TwFX2MArHWqlVbC+CoaMHo8DrF+TnpIxVEXE
J8ExB6H6WMJcMhhr5rIxJdGt1Clrq7ntWORPY6idDWCBCDXjGM03BHNzGDATjse3
5cmn7zrgXy9aYvNjBiDs1N/iS3v+Ofv3Mxdke/WmpStITcd36/wz//a8xIuCHMVD
OfbvNI06CeL1DV8gKL2zl+wf9CYxEoGswsSX8Zxhxxxiu9q0bp33kbiZocoyDJeN
LTu2B6sQC5z8maDsn0BifIcfAGTz42ntHs1kpX7WiLScTq2YhCyVkF1gkm1Tloe9
3OZC3RRCfJQLZEItH9fjimsXCJ/H3bL2dbP7LBgm0VhNE/iKgCTDuvPT84GeQT/H
+d+ZqrHpSLIqT9Z9WAdorJTtN5Vg5MWm5WfsCd/kxRVrcz61djX/GthlHykMaZcp
xK+vcMZKrvdMv85+WLBuaVjUxCbYfp6GO2vaN7Xgh78ERBo2Rr3XgGFfTzHYwxoa
vdya5N83OL6zXRI9mNb3u4mPMbWle6+SGgHbwGVVzkxiFE4OFcFPwpOAaN/fzupX
Y1lEISq4IhaLC9b2ISb3bt0RPb6uWi6uCF0qAvZkZsu+I1dUwVZGDpZ0XuDfsxT4
vP2lKRF8k+J8TRyJVnSoWDgPuxOxKFTb3I8Cl7FQGXgjQmhlhNstzUa2AIT7UH9Y
3uutk0aV6k6hfTWOisvjDEkbHVFohu/DUpSQbYnymk8zBid8OHVQSu2IsCX2PhGJ
hBESAWTKD5ZMwGcoHBcopz1/QvL5/hQF3UiWDh+2B6tu0G4fdjtAdh+mcizWY3PX
4Opoon7OiLtL0M9eKjGkkZQUw2WLpPvrp1D8XI40yrrEDCIFMi3Sj1a1KD0ShCdH
rqGUhys+tb4H4ey9vf4EStEDfHs0YRjDhb6mKMqcKWEBGPMWNAheq9QP9mCJj7gs
9HYhdT/wWQHjzic8YCoy1OPY8CbVXLesBEvciQh+h8CahDeNBizfYbl66oNwO36M
Knpsf8ct4CK/tr4d+V6T4F5T+Q+g20tBoFNIS2gB4xIPMAptqfk2J4aZQf1s+41O
vYoBoahlgXNw4ZjNF4Mo73bmApcsiTZiR7Ta51eJ6vlo5fbGjPOX+LO3UO860ykn
k4lztnyjfyVbNXZdyjhvdUab9vSG11J2iIQgFRiRi3Nb9rIDhf6TsvkXP9A8/CV9
q74J9UbWkGd/y/gZPGxS5NaodQvlgZ3gXCrQOPP/DPxamoMfpsqxL1oydHSByIEf
jcC5wjvB5Eg2Gp2oSb1n2KF1NF4XI+Rdm35LkD0GgVFiNdNYXZwNlQI39PywjOuF
AFutNRaQ6r5ioegn5u7BL1L4HFCFXt+5x/MnVWt0f2M35LGetvn9j2BN08FbZRzn
aRL5YE50zYhY0+Al/Asvn/cMNBz+iylB/sz4G7FxjIwPteOqxWiUsrHsQbxZNyWO
Am0qATwjkHGH7JvLE2RYPPMTg8fmvtYo17PnitxB3tf/exaewKzg6fQyRUSVXcMT
JkAxVKmRjk4MA6/S6kbFJrOXHYVwEh396aHw5+2siInkP6HltTsIlAFDTIlW3vEP
epijcY1n0R3pC62HkNnkCMDXXq/1/6Zkeg60WX5znZgjMLxK6BPtDCghYGy8lBs+
QAuTZtXvQXNSMfIEjbxvJUurNofCziXt7PmM26meK4fhmOtv1zZX3bq2pGeQ4wmD
c0Y28L7m1gB8E3SiuRGAkoWK2FekMmMt1zlXymn2uT5hcOi5JY+XHS0xTHnahchx
EVeALorWQfus6klzx0bDiNG+alBiyoduo/rYOeRzkA+EJWG8PumDlf1xnu1cKp6n
YFL/UvMSAug+ppugzcF25fTi9zSmb1q9RtKAsPqa/s5EtKsLAW2LYu9r5jSIVM19
+sQkLH362czYDoh+PvMQAgvfIMJnX5XaY9lOfxgwDAGWFiPLM3QyCQIVSTtCQoCg
xU5THneWFLSgv70m56VlBK4+29oFwH2AmQ9zRyhROIBPuFpznWalTTH1oNObbe/Q
6S5eBFDEcwUeSB9M+tyWUAC4iBBGkARkbtX3RZJmAu7wZOtxeeRzz8QW26JULQJD
H8DrIpzFPnpSD52QGRvcZ3AV4wIpuH4oFVx+19kDdPRO478F0NdXrJb0/qbR9kw2
NPy2Y0OQUglubIswHgFtThnuTNhPDWn8i5xWQIVTk/V2w9lwxHzLfUzKuH0OcnDU
O8pmxbdnfwdNoO1GTlfTxGFyS0ma3UHG+Iy/5PDre/bmk4QzIe2cP3u0wNHBMDyg
egAf6X6pmB1nBAz1jgK3SHpTFJlW6Bj6T0EiqFmy0WypJMtsVMxK2VZBlCJ8RZkH
ui7BDLS6wPSWLI6/uKXHyafH9xOqjPnQhbZd0vz3O/yDA+LBLRiOLtbv3KZbuoD8
kIE4b9ZMSpQhJsf0bgJe25mLU1apI7IrgIQ31kPVS75fTn4D2maRq0INxKGwON+j
NON8S4s7fvuQ7yAw5W0kdHd3e7hKR3FJNmu6nYHBl3x6vK6WOiMnqgJ8c7Ebffv1
cyf7X6/QSf9QhPc6PZKuszOmvvAzZYHlanXYQGm3FMqef77Kc1NnX7NTm3G5Iyi0
qDYLMQIJN52ieDLlyzgXE67JIr9HhhZfWykpDm81rHK8AtbdvHKN4fsaOj01ven3
Oz2WqUjRk/iAMzDsazGAaIZ+7n9zx/EXaoEaVE+zdozdoeAX9rrpKfj6/r0ePTbO
7lJuJqm2HisXYXgGpHu/HcaQ5szDpdh8J1pU3UTCU2RT3yjWwWwUTIriJu6RHE/U
kYld2EZ/fVQtThkMpkhWnVV24CcgmG7r+PPgW8dJtbJIwlcVzopffhZXFgCDSx4X
/dy7mjpwrCIxYeIazKcPnYtmNnsB4GMBQbEdSpb8kgir3BN18xIwSSjGEkTku9JT
TK5ICyeuad3nkyLCgWh+6BmgBMNT1plISlg9lyIsuZNnB3qEFdjIGx/dYCw+yzOe
FwxJG5tZfzfMSxwL7mC8iDOvu8Ke0yLdA73bWJwsrZOsHy3tkqgZcLex1dcbdDVp
7K10KoW1s6uSILhaMvENnCGCPYYzjmMCOaTIGJuNKqKcx+YLFREomdaVdJ/WZq0g
3Y6jxcErWD197pCBEMocoSvtH4amM8gWFyM6qWqAYpSNWYlT9pv3pnuAMrUHQghI
dNxWmy4SdLNi/734aJ3gD4LLyryP0aiHDYjB0bIkAXWddMxY0E5fZVTunJOAzSZ4
5gyr5QyNpMBgOCtjqAwpeSBc74j78mKrSK187+hpXidXe32Fh7YgVetu688qyhdU
VaREh2KGnh4m3tU/ydRiXxf1496CbxzqUkiJVxb3GnS6zqotC3ZMi3rScW/LBjgE
2QVxAiePC3o8pEMzfZmPKIqSACUeI0ys0piYt7Z7Pr/aPBJhtAF3Fn6wOuspNptu
ysXq1JxlmfZ1XRPKG/XpW1IAxcplA/AAIBxeQK1MiHeRFpGG2vBN6wKBowsqSC3f
K54ceUfdJCHjcIRC5RWx3nkN2vWRHrrro/eiFw5Terlc/cKkawxNzKGGh19MXiGt
YoM4jCQQdR6IiElnNxi0q1gcmPMAtQw3IVu8nkbus0NMq/p3Ele7fehr5oAGsR6V
aDZgObW49DUD6Y3nhXYvjPTI+TAFz+/LNfHQzusgVs8sZGIav2S6L4uyRswpBC71
Eu3hDW+mKUOXeVTOdJqIorxZ4o4zXv/jl/dvXWeV4OLo8LozCuitp39h8APfxujp
88cUGKlWdpwxjefHzVtSWm7oct1MGWkt3PIlHrOYgQhk07NIDVtVDEHuHLPZDfBE
QE8aKzanypDsqN4EUO4ufA2TDqk1wYNxhrAsZyVDn+J+zUkdYIOnFHV0XrqB5SiO
Bn6B2Ngw2b0aweGuwaapTtBPbzvwheuC9CyJlnOAcOxIT0bvZ8URZP277MiwniVw
x92aU38mc63I0eMDMmqdoMGujA/QwncI9sGnOM+DncftKhgRFXZeoPIJj+0+A1WG
cS4R2f75cP0MKY80mdIJ9XXU1s/oTKRDKYpJp91DJ3MUqSM/n1i+NO35y29nkuzQ
GheT/KD6hHq6h/39rlnaweB4GAIjVXDsVtOUjKGdaLvi1sawo5IC5zLnex82ZxD2
2J6O3p+JBf9Hfdi1+PpSDm4GmR5t6JnFoIjfZ+J455jV+whUx4dMhsQ645QfDSEK
Kbs0qTpl0tIso27Qnb4DNIeIZFdBxSWJ620wAFVOZxYtdylMCSOT1ThU40gphslm
B7hgzutGswJ28svB1ZNvfXtN2B+uj11VyfY650BcQUSCdjnr7zNL8xQP4vShjzq3
Cf9TZWDC7vIgoYVcyGgFFd4IFYb4RQmM3lQJ4pcnN6BEtgMrKIpiiSLY5C24qvKy
QtSlsW1LgeqeWtlVfh8EslJ5KADaGguUnI+pqBadglimKVc5gzxICuSqZyCqZMek
SN3auoVVD8QhaznyioXFG2TWzxSrPBuXjKOfzo4NAJLpUFAUzdq9OG5fq3ehnwXN
qg/bqdofg1FOc1rBWP8FNbLsepUZMUdInmYGx6GQQjdGy/NdtZqLzyuwtqF2Du/6
SgyPO0sP+MuxJjSz8+JNLCJdaYuzTLToAjA7fIZCIIGlsPP8AIIC900TrQ7LY7HC
/bVPxzTDqXSAvML8vo8rMcxTHhbKeBa9r2Nc48RDM9c35gwpabOlVWZwmMWDpzSi
ebU5JYVhE9qoJyUAElOhgH54WHb1ras/SJVD2MGra6QF7tt1Ru/qeILo1HFtFqKM
s3u9bSccfXOqVCtlSBxloIy+XGnZYJ6HeUyrRlmrrTNhhPgy0ifgwIqtoAgsBQHY
bTpKoypd2klYlJnvFm9Mc9DFOdnjfAOAKzThtRfte2FCrWUOiQaKT8t6P8JK8Ae8
nicoGvslDZcqT6mO8OTByvoFPjQqqbxGqVCKwGcTR7R4DWlwm7cZz70PL//Jl9+B
2e7FfVdWuMm/ARrvn5wMZm9flkfA26eCct3l2oFLGy8E3mqpKD2esrJaUMwuLnb4
Nv9phBSI7F7oR/SgUSpWAj/fEb+fr7gPVWYJeY5ggrokMjXvGdaxNg49TssvxM/c
LjW7yc09zkHx2X+FMScydg11mJ9Rzo5MzyJ6KV8HN0YLN/pYtazpapzIY3SQq1xF
oSbP6UDUqSAvXN/XdVwYjZQymmuWDGj+K9bhavfE5Wt6BTuA4MkXy9FLTBAbXerZ
UuShD4Zfn19JrKaI9/1LAV1QpIKAhZjd3mUohOgKmht8vtk7X2LgidSKndSiSTGi
ZCli3RESB0aTlbhySDZtfHwljCh7itE0V1QHG+AaYrF0lQo3epUBkMT6eVRpGD73
ri8oVvLuNf9s8P9hhov08DjPSDtkFYhI8DAs/RDbGw6ObfzReohSeyEFCY6Ov1TX
FGm+3nzjgpPzyLG+hNk6eQMz+T1hUlstyrvTG+4YqoPeZ70EWlz0xsexNQ4EJPVA
qZX+9FXXTYD6M3KBTZD7cYHN73HyrUjLab9BFF3otqEidXlF62yXsy57ro0lDuh1
nJNbA7ovnY4hVPP8YfeV/jb9Cc77qm52RU3lhQFsNVHITKCDrhcNWa0a0XqwsD+W
ySOGmRclbmwXzdHkr2Y6Hef858w6S04MgbPkOTPEVS9NWVcd7puxv8mJqhg/qbUY
gqB5LiogJ3jU4zXb1sKG4HwNTt8wKa/0ZhbF5T4dxUYr5INMufQq4hgl0RGAVldu
o8quqiV77dAQpAUxJdJ+3EkfPa/UpKY7QG+VS0e7oD/pfK/sB0wE7gZM3rJ0rhdS
T7iFY77naFfiOYxaUdLN8mCUUti/giGbFtVEeaNhlWh16EXQ/orlSVhmz8vsFFZR
juOU8OOD0LesDK+dZyr0ElKJ7cCBoJWTujKFXJst1fr/WvoP7hnhjO84kiF18+lj
o5PdaWsabK5BvXUE3Cz5x96+7vkMHidD5R/1kccTr9qvOhYT6BcVtz340DeHSQx1
VaSjG4RLsXTAAkY2mnXrX2T1Bsuyk3nncNdmD3TlGYRyz+MjvHT4GqNPJTuPIiXq
xq+evcnt6f7fZfHOnACCpbKvKwQdRgE9jPKRR5aPYQDaj1xAWrfmoXgWOEUCgoUN
dXsn5SS4QbTQsfMCX9WYF6/dhBjL710aG/Vb4sY9qlz6dOXtiNF7sqecn5Od2ayu
yhh2mB+A5z2i9Mvquu2UWuZ6RXfvU9TqVtLlvaDtB7izFDP5D0uW3gkyorv7Oaa4
ibX6pJqLYXX/MqVYjFNAByIbv7SB+ugvlRgpczVJr+4/SrcSdQsfpnQBsDoCiprx
kKvnn35Sg15Yf8SHdQfSa/gukErMlW9in+eV2olTCmZPwfS7BarePvyVjEWIgKFM
WxxEOot/B3eskE+zmgy19wsX++40bZ39xNl3jMeSV54yvYYcJFX4b5CVuFnLMaiJ
FKyG9RYX3Io4Zc5bXOMl++kvJCyfOn+AJQH2TTy4sBBTJ2+CH5AiMrAgOuefj8AV
E5RkcNpPNxwl0kppVyqC1MKmCiCWf8PCqZ6e5v3Ctw2+WgYSJry8zN7DIFkAz0+B
aU+LzZ8MmwUql33qMM6AW0kSC+kZHSXWPvkzzwIaNr6fX+vIzVjk0DHaDPY/bI2c
pCvikFRuf933BHVal4JTctO1LBoDlRIsnUO6QcQV817RQHSZBfH0z6JzhlDkUupH
04/QRBdRkaFiNTtTL55kOpcb8OebL5tD9jHPUionVt4c7AkWBaW4iEZiQ2bcWiNc
0h0/+m4CUSpVw3rt5msNcbO9oOFbSeEoBBdoKDXPFRnzhgNMEpbGGT7RIBsfQUKt
0Z+5OChfyWqMbSfFD+D7A1RbZMQ3H0OWK8fSWY3oCbpvsWLBDmBWRg48d1rnd2ji
MAF9sup/LkpuZbAIoSLW6o/ctI/k7oTiociWtrjjVcU/XcqO8ELeBPADQ/qoXV6t
reXm9DV+yPSLRGxV+Nbe18KVDkcd4ao8U78/16HIBEO00M8maX7eVbhH/NYTiWqD
CyrOpcT4op3Ka27ZKJzXQGBSd+keC7RHhG4cd47h0Ja5JfklGry0Bbd+39660tHk
/+EO12QlKe3MlgY9omqnMMjagzhTH+aQMlPJldqSVqrmFr01gjj2bXTBRgCUYYtv
rhHwtJVwecQJXj+gkgYAO5WLkQHGZk+etp69jT3DI2johwpGWBJIR3NlzS+rVJIR
95eoEDDf5BwqTSZ2wqxTZxR9QjMaGb+I4uiKd+0eTOLVWCS34IKRt2jOxHfTzC79
6po1AZOrky2tLOFTSyrBpgbSbGGdyVPmvTs7Orl4M7NbZ1tHDXIkMMJhJku2/Tha
rYK7i6HUDB/8LtGEtJ2T+WnSD1+HQCAqwL/0hEXq32BsUCMv0Qf/Eog3xhnpvKsx
jAGzB2h3DC7+r9+lEn406TeVBR93m2GWsUUzl/07drVRWpN0PsEBVIfFWJU2sgHl
uDutDA1Yeegdr8QbnrHlOcYvJyfCnv7FSQMx2W9YvG9ia5avLyvQp0UsG1TDEHM9
9pe87iFCqv7g4Ze+ONyFsA7vRP+8pFG/SndRpPiXxRTXplViShubZKzSpbR97aGN
2GSwjtyTscUFdAs12brhEwiwZtb9w1OOQI5iGypJ7x66Trqyk58q4GiStCc6sdCQ
QgdPrMCym0UYJ8ZFWpSUgDP12AMUBojQCm3qWyB+5egYS2Dpmnu6PVDgYsYcdZ2d
KFJOj4HtBFcELq1Lt8cvMwxea2L4oNFGtkUxEMnU1pt6HSDR/88v1FbivKyx//Tz
YkBTvW5O68s+IgrvrndgAN+1QUWYnjJsl4v0Qw8jpwSVGzJfAboE50yt//Era75w
Zu0LR9wA/u6Wjh6LJAZKuOHFXjd+GcuH8VCC6GAHTCjGzpwVHClYI94cTKNRQhn0
/Dn5lf3RmDw0pO9fx7SeU7Lk0vRxftEcyYwoYJKtBQHjnWvae58Bo/Wm6g2fSTrQ
UWie+SMLm0dTyJogZnFydLyuGFNPKm+yVpCgROp8dHWXA8G2Kq2w6ktrM5HSpd9F
bHEcO1CckMGb0HkxUcI/BnOA4xf7b4Dh60dSN7vEpUuRCDyYj8MHKpCW61x+9pE4
j0Z+dtP/scrjzxkFbV5lI0ew5c5+LPFXOk+1AlmmlXoFj50L250H6iisIVFpqLcs
OO1piyG1gbtGb7iyb7K5bHroCyoHX87HEkoDHkh6azWDkwXO1rBbfdsofhO1DmRE
WGf4tyfbNKrYfWQxhHVmp+lPM4Y8gjWXqD7B7LVH0PIaH6QQlehJFHZqSCfdu7C2
VyflCPFQhJPnezOviCtPqCDeeqGHUdMees53gvHdR5J3AlJd9u7EDmDlLLRkjR80
fsaeRwZA4oNhkWVQdosL++K6Glgjg7dHtcnwBmraiGXvaWFWP+0pIWZ6JKo7NQmZ
28AO+QaWLYBYd1oZ7uH+cySGblVbYayK/rH5a+wzL3h85WQZQC7kuvOIAk6plsex
ZNOWuY5VbKKIuiOjGKxXyUshnLDbtPgimGp/fbqo/Mg2VTjylpsYL8dycj8hUSCv
7KppZFdTVNckhphrz8oNc5Nc1H+ZmT056bBMnfT83myiJbCXcqRAq7lRRalWM1r8
ugDVsfAhZpgB+dMsB2pK5kABm8vTwho6NZ0ZJ5RdihBEo8ZDQqZykommpVKTqvN4
o4GUjRTX40Sv+v/MEE1eVJ8SMzj5buI2S2aXqpeYYSJJ8pF9kqO1wJ3B/uARdqPJ
B+6OjGqFeuTuwnIW9zM7DAZQ2RM5QbDIq6GHNAs3cY0SU0n6xw53vR2cZPDdX5lI
cO4OtzSIme8cMIj0D3iJGCpiytbz/TCq78AY+BadkU8wJB6yOrq26BYQhrtCY6ol
SRJ3WXgjAJ/NY2UQ50+Vxyof4aV50e7QfC6P+kX+7JZNh7DhaMdOcgQcJUhaSzgo
2bORR4Pmgmpf15yQHbRDgl2oDGtED63z54R35iVunUd3YZd2p5zGUmdWnlvgSPNg
DF37bi40Hmge7zg3cdADkrKF3hDyP1fnY+RDllqOrZi+0o6hbEtQUAD8tM+ew3Sb
L6MCG/0hmp1n/+Tg/df3NwmCph745197o6kjvwvMK5eC+YDiNTfgryUygfd56cr0
aTHlWcVfPshEnI3gxhowHhS/S+wrYLrsPZqAn5Sw1GPNoQZheBThDhjBGXiqQXiV
2myZYIfjWXETG58fkIg1K11BA+rjY32sW34PhgSXu1xHRtng/jAVfGLGq2JaNRpL
kAELFKvGOPxRCvkYbNQRHA4l8sMVxUsqj/Rbt+9fMQmByavc5Nlx3g76OW4F8zi8
e9Qojdj5hnK0+tHLp9HI7nqXRkImafBc81DtHTgKcWbRdg9z0WFFFftWxk7tv3IK
HUaz9ZRpTcBtEmCblfELBoRcSaoNGJQbilqDzm06bk63XsKBe+gAnVbO0a8uayRP
fCkH9hqYhYaCshGCQGb25xEi1ArxPE4She8ad7q9B8/GAd8mT1gRkawgdsQSqkcE
H6hEBHAZF+k1YYoEffDUQsPI6mkINDATV5GoetszEJBhY7J7BzKCV4vNh63satEx
txgbl0CkaHPmCgW+0TnAjj+X1hf8+9mHeD0kLS74381y4RYdbZeSmM7A8FL6SjoT
6yuGJjOBMTvf+qJ3H0v5t/FBegzu1E61dQkcjlZdBaLphOilrFMHoCXdIoz9SbUX
cPA8aM4HClNL2qU01y4nkGGseOlbzr0ZqMm9S+eudIkPSKVdUl1lzp4TEQ27l08k
qPYQEyIPOUgssShHB6WFC4O7Vzd6tyDd1RKwfoOjJD7frNHkKAgqImbiejA/bb+S
3MA9l7jVbtjed6Sqm2bdSLUYz3x/J94ubwPJV6ZTfzmtr82yZJm9qXb6Ka6SALlH
AFGpq2wBl5Q9Z+56bJBhW+u4Emk6/VmNaqBegUA9Ja8qQfKKCNk311ae9jCyzH4p
LZnJdLgNWysf47XTFckYAa6yeW5CyaQev2rCe3Wz1lHoJlWkCFiWosGg382uobPL
TZb+nq70lTTM7umMD/YhrJZtYViQmHibYTVSeda+fXp9cQlva451Y0qblCjKG97V
rOxU74cd52tyGXAH5KpsWjIBf6osZflHKFSGVkvb/84w4FUqtLf/t7p+6bsFKgPB
hZO3VA0qG5N4718DPZyFNW1K8ELBGVZ9zFvqK0Phcfy6Z/WjhW/87u263B+gmhJ4
qq7DIVHrpMf/+39dDr4BWcNvIjHkJQztmyus4crHobpUVlDwBiWU3o1frgjlWYEx
k4zCCucDIQPKP9Su2L7YwOZjcWGr+3U7+Ei3MT85IAPRN3fSrYDJwO93rZIiCZa4
ZHOQ/op7N7Z1hx5twNJzAyHzqB227OOo13tDlRZQU6UUssRIxqhC1AA/CDXcnlJb
1UYEL6tg4J/6cpn/a9sRs0DpqzXIaphlS7YWa8ZKKWiULdEDfH4I6uChk9PWAWN4
cjIY4iiFGGq4rQGt0aLhQOloghK9lREe/SlQS0K2lbrzUMmedRQhsLczYybgDN9R
bttkwoeyfDxYevj1HOSbMqAk8BC8ATCT8+gXKys4jmvLcFQTRXWLtosxuZGHqO2l
oYkJ8VgBoQqGxAsSJPiqrfsORfHPp8s60yYanQ9zQDkBMBWOMfpVNJ4Bd8PeJkM1
KUffI5HLtdMhuY7kqSvLGEv9mwzBK3Jgr/cZo2fJYmpto5RalGzdRERDjWXknU3V
Qs/tC4LIbVbkqV8qbZjPX3hRKHRiNyeOO9UPLbFM9Ak1F98YO6LXvMdqsxSj2OAT
qVWIz8NCsLmVIasNtEhWuseqknEvgK66UWw7qwEnzDae9rUz9x2hd5J5yNDoBRh4
IrEn0WCYYzNaYJEM90mYfD4qjBFsHw6jlp4FySY1+t7Ae/ooJwrY61QLPWyESRpC
pK2OyXErh0a6I+qIqQkycpLj7TIDZvzzs2NdVs2ACgTZFKq7WmPDZoWUfUgmB4MG
xKNhSHYICCDcOjBWTblQoBwF6S1bLQC8oOrtT0LLSxO6zJjvsxHJ57IvYy2lJdUP
WgUCOCv20QM8T/g9LQYdSHb9gxH/6CVLf7vS8qxYkytl4kSq13RyPptSiZzjR4sM
2LSnhOkGIIKBaXibzPwdeyiH6K4pEnCOJQnwwqFP3IpEPALmBbvcBocb3YxYKnD2
0mxufKxwbkVpVcZYEG0QloelypQ9AZwj/x/cbuwGI7zK6l8EdyNH4M78vfLzx3Vt
Jh0gmRbeORnxj+e9akNLYmP6ZgsqInyIqhD99Pl2Ta8HH4ZRXEjRpj7bDkwAzgzB
QjSawAQIJIKz6OjnG9GSJdtRHr9kHbRvCrJMYsWFan8o09qs3KchAgLy06j91Tqn
sMoPaondA5F0Gfsx4Xd6IUzv3A9CVPa3yqN3ems4hK+4qUNE+n7H6PvVotVcmqjo
REkTYdybwOlCZ8YjJAvR1+iDHIpMviyViuUlanQHp1woXerZpNDCQWfee9R5J7lG
WyvuFRD3svhucGDlo4tsA5qfc4SePV/ZT95CEYcUc93rs17ajSaHF2wEFsCPKI99
9SIsOP8qKxDEY9/437ms78gWGE642kiHbVEnRIIfcge5RQD1a7eQWGuTk2Qrt3kB
nKF9aqTMaHkoHv9w7EO8wm9kYdxCLwQTVK/IQFIB6FMIR2UT3B6hv6nDG2GkZROW
m9iMJeISZOTgrAcZOQe8MT8hE+aGF4caIl0a8HVtRQeu9aeA62ywD1z7Ni0fdNkO
4YDQ8rFADWP7iy73dSCgCVZEfBEOIqL2sf6BFUNLmwuWC+r8KZw8CZqxCCXOlrK0
juXk7MLP8Q7DACacHFHtSZHmMLeOuPqneW3MDJZZRNS6/CDuLPEG1Bb9vnSk57qI
zCKKTI8Z/v+Lmzdsg8pDKKtqH5QjHnEvKn52ck8ORpVzfN4r1MrKoSj+mCkGlzDb
+p6mnRxcY11S6NqixyY1wSS4PERx+NROV1BdwfAncI93hAimAjD8uCdcOJB9J49e
ZN2v68NqLtfuoaHKWXeA3s+d1AkYBtgtR+gCmigS4fikseLbtY4N63ONzviMZfD9
Vlk70WbUwehALOtqsu5M2CJv8qvcXh4RQNaBR2vsdajTXnjjf678/NFYkZyNcnZT
LBQ1yqNLIC8MclUt7TgBkH0bDPdZW0XMvQIk1tcJJR4giyXpe5KLquvury6VJz+E
esBf/31drk0UkvL0DmPox43rwZ5BYe8TYYstJ/sh/oQg5ZqDSfFAlRqyt30NuCFC
mwSx3zurGtpqW6cbJzacLmwO3JkoLODGTycId6q6jhglZPrOuGtmcFxgz2hw1eta
0qyL8VvCJ4wYM0PChfjlxUE9mOGVgHrxzM/B/p9o56CwBInlfYD92o/9jHu15Soz
waZu6mw7Mhw7wYVFNeb7TTJNAVSXHAYy8tTuLLm7EVWUZyp5tnwdTyjKvpROUgIN
OcCVJPP1s54Eo83WWVH/KPQ4t3gnV2QsTwzZRHy5GoI/cNPZqBdKHFZAu7dl4KLE
q2puq1BUv7AvtnonU5O6YlSGulohfIf4EV9OEBCnItsSF/bPeuU8cBmEZcrZWfiA
ZrF5X+HOnV6FZ5kQwiBSJq5YNJTB0IEYiML9UQogY9/PCP+qci1wUvVXCJdPZLyn
1/xYicgY4eNMSiNVoYhT62dCoEElKBEco0Hr+5HQfPnZcpzkEmjtEXgRPUbR+bD+
3Bw3Ynwk2RANbphULAm6wMfHs8kgvi14+8VqfCuQxrSwc022b6MrL4c+8hnwR4x1
9aJ9Bhcq/wzIQ3XtRqJYYZfnQ1gPBL84K04Lsx0Rzt8YsUKIT3TjgemYX/iOYL/P
Li6fNPp4KWcBK/DOVecwgD4qG8eMQM4A8V11eQHv1gh7XdGLA0T0kk1Ye7n29wTY
lxF8SATOHiIRANc66gB+Byug2aRyterw/FKnBYHw50isLtUonYUZPyCwnNqmtGKD
6IovOBw9KKXKr7cazCi/kWKAyYVeP7VNwmGuwjzde+BBF2Du9oftiYzmhvKOKmjL
VjuYIOn6C4NHjToCTCTpg1ThuSxMQg8C6mSgWLqtPa2c7iXyxzJmBX6dWTQ6q9o2
Yd2GYrm0vzhWfX6JFm7y5dVuYaK4zfZGhwudkziS+e/7o8p9tuzN9F8ejEl7kh9e
DWZRBQGlzxUe4/dSMcB9O4X8TjyEqA0YDgGzH0t+JnLDtKohwTO2iyCmgoi9B/8L
uwmPdFC4wgNW8gDFrZ5ulVwypTPG2zRScls6OZ1IYC9nTBXnMTkbUc5vS9zdee5q
yXYKw7KI3bU5tjupGb+uq+nMdeSf8QQy7WteaPY+hBqlQgspRHI17mEumjSsi01x
RoF40OgzKJ2/tA0Lka8G0ob9oUqjDlg2UVJs83TNIplmT5PM2KamW3E4XGDN+KdU
zkPYXn0FoHE1zdKPdYiCf0j7BXPmiHbUV2JaRCp9OgF+Nw5/8hkgfXCs17uE1XvP
vjnlMBUh+9XHzc6RNGFvW5Etz9SfH1/CpYYeo/iawboL99tMs0UNp6ebGHrT7F2s
Vh1RaNv9/76SWOBeTjTv6Wt+TUaSDw4/jtUesbaiYea/mltw1S7H7wSjMLqIucyl
CFpSAayI+4Gnl7MfsK2IUd++wAu8IaWyT1JpnBw4swahPheo1cKbig2SKp/7HkZl
PTRN3SQZF0ktoOkGAJFUa3buixsTGlNthzt5fYGu78Vlzl9luRSJFkT3klR/szGw
SadN4ie4/OJZVdMH+d92ED5nE8skVd1bB54Z9P/nMdIzXN+IDeZTk8AL1UQxS4xi
VLLhrd4EGdlU1vpxglD8aymL2yfh2VeeqZ4WxMt8peC0g6/llTLDi5IlRfWP0JDX
HI25JpAd71a7E6EhFb86UP/Y16dW0uMjzAHt4w8TZ3/62MKv3tQX2Zp03UdbxfPw
oaD0gjF6QYHtJbltD5ZfPI+T+wbDd4AGDLaFg7j2Cln5f4xBZpCGmUvq9Y31ZgFM
pDpWs5EunkKFRTaeEOQ7z6OfvCVFVoy7SO2SngjibFhh8SdCLaYn2YJ4XzkX0ReS
SQ46vgXPLYSil1MOAnYHpMni5JTwTNALJgjzOuazOzSUeLOPbXQmGyMs3hjU7xYM
68rfSzsyP6cqVCNHZiRDPhq86vyZGHZaRrmMIgGtelEtfZEcGSJ9MULnoJEWnsFD
eEPfKoxxW3xL/w8vgwk18whcgFeZ0bnRHMhUePvpvxAehvmQMBwcSNtDGZu8wftM
8iF4u4vf50P55C6AB+kz51/LSs9XPxMj7KCb5NtaCcTnIG7PPdkvSenAWPtLWUAY
T+H2M+G8wPpZnRjmR9I2PsdWl3xpJMD61COhnOgsJBNRnvOEFe6V871ep4ZGeKop
0zJ2Y9SBeCvmcBXSSBUqZoUKFhWzEm8yC8v/pxn61hja5aJDUis8qHyF7M+YYz/m
qv2/5Q/lqfGw7TsGpN96GiTrh7SJR8GPKzcEKSuISon9bP9QIxygr4RCVMhOpJr8
yUJBlJcxfQCqvnTdFNJ0u0FfljogusDzxYc5SHWLLpJigs6KuqqBcMaP9PuKZZgH
jR6sIya2U+NCm+5V//GxjTjTUzyhkSiGw78fmBbqDxHd3jmhK4d8NcT3mP+gZ1Y9
6VLLieXT7tcrXXyW3EHEcOEBtbi2FrFtX7kTzwkRxifQomr2aSKKiC2gAEbmrJI+
H+yNnC9Dli6i/mFzZRGguH/X6UXJyJZ6oH7gUCnsX8YNHF5W6+faoQKGbQwUVqdf
VgqhH+Q0bBLSxEWPUKoajZdGRx2gz2gShEWtjwMmYfbYtV9zRlKuMTzdwedcW5P5
XblC9i/5g3tmkeKW9DxGR5IKAhgav4wh1dTasKdyhZ39sZJifRvp/E5Bdsxn1q2+
3tq5kcxUo5DQdXohPsBFMeXhLjMMasDGS4IGDhy9GdFuUxc7wR/Q/oAzlfDnR+uL
3UP2J5k7eyfSNhB+Kg4cHlVQpLrDgpwEvUIlVs5vrots9aF9ILH0SgDcTg9s1nDs
Slw/Nawa082+xN2zrjuOJmcTQbsoY0SSRKPik/9/meg1SV5y2zLvI9lnCOqk6hvr
S0JJH3Is8HfLKoNVdKz5J1IKY0eSiEDqMX1IDcP5Tsr+4Z4d4wN1rdygdFSUWe0Y
YCqTaFAbdAxaFg9oqmb8DTu8k4dyYvUYxGmCbH+50mKKTulLOpR4fGl5/mCYJWwB
bPXaQHQOK/wPhmM7QLOXaqxEFA5TnN6xA094wuAkVYn+wlccgp2qxOmpRcaYllzA
BgcCfOoUGC9UCCFCpOSqddc7oA4wvtXL0Klg2G8k2Z+0BhOO/1y8Evzi+OyZ43wY
J2UToEvqXe0pmQwrolwsukOcyF7aJB1K9lS3TYehWsrJ/cT6n5ePLJ+NyAt7shhx
evA5ZC9WsBIyCR+O00Qy5MS5oNEceUc8Uq7NkXmZQS9oEJgwdAR07tlZmRzxKGRQ
qTVKzkBjTEcBxJRJ332t1/p1iuCsKKuh+p3CYdt8H23/tW7S4XwW2eN8GgS1Igll
kDGf/TmXgLfbJEG5equaducIsY3COJejB89MSUOYnT3+MhSvraAVSXCBF+XWcsFw
wjEwq3jP6DUqZTQym3w8ItSrAUituFl8X89dXw1Z10mljYGoSHhVf9FgcmcAjdxv
6MmA7ug7AzwWuboPlUFrbmxAIXpXTCUbw8PTKye3BT1hW01CGC5icNJq9jWA4++8
ha81cN67A/JxSVNPQ+5jvD1nIySlY27ZiOWBjsg4y8D0PfND4UCGgrX8IHuy7kwN
HinbH1PzIgzIDX1iYE71yVZ0HWameFFjzzyQwWNck49kya3QPbxibR7FtCx4VZJr
XxozWfCDlfhv5PeVeHI/d245/aoRKcdnqRuYDPotIqpYOvIfJ0tY9/PbZJzxgaUJ
nmosbDfhO+6fUFAATmx0mcnVshLnZM+7HSLh5FyAdaPj95KbnqCnNor061qs8VxO
zPrf/sK05ItZWzT5kaI7jsCvB+Pq6AhmZ9nATxzvIsKtj/slERB3vdzqnEgb3xmr
JfxiuhL+XyeZka7EcNiWKBof8dcxKBujsvw3y7NZcdtYeYwr/qy0B426mL2Qe7Zi
R+cqQB4L+qJIXhxp/3sUp/2/qg4HeWYveDlwTdcQ43nRK37EQdOaiztWww8u5oQj
Du6t/EgWQlbDNPSveorDPr5jbNWmSfNPt538OYOCAh6Hshk+OYUPFngnRTpChYWi
Z5Lvn/RbLdEZ3h2JXbvatDU//zF1B9nT+TZXcwON3lOLWScjXgUboID8WyjmCr5p
OONFirScbLwnlrGbP0Qwr79w5mNGNk300iDrkqRqMcNybcAPBRRFdjozOs0Ms2n+
w7iUOJ/guly93E/Gnrm4ZsNeR9DaFpbFm5iNniKmgKTZosXYrz+trN2g6JI8kwhS
LY8DnuK31KNla1NdWMNz+f8Zt2yqVJ3LO5STpVgS/COkH53qV0OYLP6ODjAmx9J+
z66kNaY5L8l3QVwXfRQmGY7jTh8LUob88s3tnC1vUBpL3+asfwAsA63B/f7cfcpZ
n+HU88bQUFBiVeyMXj+rCcmrWMuhBQnzl/1iPNtaDZNwyuP0SPIDocRwJ9AukSOy
EoyTjAFv5nYx1qCb7J7FrT/NSdw+u0wQ6hhTumzAMtVfopozYThkN5gT/EYiG0k2
2kvDTzGFyz+c+st23/W3/UVqDi/thOtFXpXPdIRmIhcXrYit6Bqfs50hckNEhZrC
I7Ap4fCFDpdyVH0QWLY8I1u1jHmLsFZ//vjH3bzZQ1adDxXTRu9FpeP6eqYQKrZs
+mxIJCgD51kIUFLPaiHbYlcp0ETa0ljYybd1byEmTylBkxS9WMI/D0eOJ1pBFVUC
04YWPoMDZOxS6ZSTTa2dWUz7qoTLU6wHfaE1ZEku2bdjZzgnaK6XWM1t2Vd55WBt
SGU459e/zGq6tM47LRsXUMnL3QtgZBerPq23Sr82oP57y0GhsKMUJBKxMY71L79F
KqK0PV3BLWAYUJ5I6IDfLVSFh6HrZgm5O8f9PKu52MOSTq3T909oab2wd/Lqr+Rq
bkrlCIm3YC+uvLsbUNIQZaKJWJLiJgl68mcthrwNouP+waCrAHYlOKW/g1Jm42dE
be93Tw6cezyjNGxEfEaodqq765sYIlVVoImpsynLKvgILbFjD+f5KTRtfU5aCJSW
zNI/X52jO82xJn5/wlE9GXN7wePyeBjI8S2C+FNEyiBa1VuxEpvLmRCaH+i39v/c
tU4dXnAqRNW1sSHMuwnxWih8NviEA07m6q5u3g2Rzf2qwO6LuQp67TSXL9YpuHWR
Gy5iXnnyX1xsERnfW8SSFNT9EXdAZKdNmQ2bDRtBlqHe599yuo0PTWmoUFFMSEAj
Qc0h1cKqf0UPXvRmL/YAuoMzfWEagkR1ttAJIRlJnX4Wr5Xwl5LpEX8QKFthXuqg
wRjiYUMdlBLn1rF1P8u6wxjAz7gsgbIznFyOrWR7FoG4Rge3qQUNm6uS7OOfOoso
L1/Ph/b5EAOg8F+8sPC2EgjUhwcGK/jylvAPAUsdLshsdIzkk6BnNYR9PSEIry+u
I1S0Ay/q1QDgVM6s+HFu+5rxOuk2s43khyn2Gcp70+Tj+PpAaRMncV7ERmpLg8Ij
ceCNNIKWDaXJB7CnJWFsr6ch1RC1i/z4vPs25z1UXAl/v16EPXwhvb7+N9TGL1r3
yBwHMOKQpMwJgcyPt3xCDVVIAp/kpstl9ZTVVD5AQroIe0RtFlkqsUkPPtLZrURf
cq6YFp0xooFHXgiO3XmqCCZ1XunYFoZQBKueSnW4rzIzQxgwA6oFy8RNcRFD+eYP
eiCxjE+Vykr+lAVvQlhl176cqckEQfd2FO37bLn3LaouINr3Td0pNe9xfsfH8OrP
YKdPQXcOKtIHy4IvO8T6gkUHd8ZcygvUkOMpU6RVr1CrHvnmwTpZkHYS5VHZMEHn
C9tIJmnF3UbFml4Di5zmz4gf1DD9cL3nz4MTskHTprFTMPdiCoLygzFfsdSQNOH3
HPrdFsZJ8nEeenNbBYvCLjFI879q+WLGZwey6wYziyQ7qj01HXZzD9Yclsf2av8l
ZwsUFxCVWP51aMPqWJRqi+PJZ9G2MrptpVd4O48ZHwF8satmvVC6Pgw61iDokGAb
XmQwBPPdJ/oO3/pydHTfd3i3Kwz/0sxUYU37BMRxesU39APus5swnMXwLm25wkdY
KcxbJw887MTZYamo98jeW7W3OEoPLmXbt8MmhmL5ikwqCItDYhnlWD+N5WiUPuvY
Uj0+d/eGzjOnusOp620cM8uqTB6pUWMP6mwTwNzRbVloYZaWeyeq2pBns7Ix4KJ2
DltGRfJSqmaCo5NQVl6FipJBocCdhsNrJVVzMpBpNHyNyQgRhlJfL39D6aeoMCbc
Mf+fyoKjWCFbmhIEjUaOvLoVRh1iIclHf7u62ZxZhtzEnpH7+QhwCLaptoBeSRud
nEJflMxEFhWna42iU5uvuZx5ju1Ibuk/qqn0tL68T9fFiZgNhYs1rzJcaP3I39ku
KWEl0muN7jO1INpCjWYOiKEu7cz+Dcz15w/WqnUw3bYSpse4UX8muF1z73BIChiG
UqplLrYzcrq4+MoYy6UGWt03zwiZtJFdJ5wEJVxa6eeVKyvmqF1J2dG+6uyKqHjN
3j6wYTXQmzOiFt0Sh0jvtwD3+i0pU7a+007wG+E9QEryQZRD/nRR7jIdTvFTRCkd
ng+Lhv/GDQRMV8X3dAl4ov/Bw+0AmkLa7R2Ur+E1LARMDlR8Mbes5p7USodUl4Yv
ADSlvhIZ1xZ+Eh2e5bBlc/vScb+iqRabeaueIxxJ9wdtWZpeuOfLywSusPnvYWxB
AN2bm3XE3DoXYazi78iwsU/vuQOXh/S6TNYF0HxijZ1240f29PKHgjEvy8buADZ6
NfWc/RuGalVn1OqOqOztdP5zJQdRACiTYEeXm/G2x2AbS7Qam0vjjJtHT/xLYedZ
kj5rN5a3I7tTn742fuLkf3nNqYCLzg90KltGtnXSJt7dz3p2GnczYwOUlKcl2QxI
XyLqj71roLO5vXiKMB+eftd7BMGjFbGg3rzkuJ3GC6i6QnQ2cg5jT/ddNu8ufxn/
QghCQMcbFjjOI8fU4qbyvrsNBl5+CcwCRwz8qyB+e9gf19z571xZHE1EPsPlA7iD
Q8mpaeXwKfXkulhcd5cxpnCPbKR+nK+Tkkb78d85OschMPVTL3UKscuW08Ep8MrM
6OJfgveKU2lr0guwZ7QObfwyEQgeaefr1EERGGsoa+7iymTY967yuOmGoaSl8H0h
yhHgqdNvoFxZc0MvBkD+GwyRI/Vc9MwIdFJDBvoTgGbnvXq178EUus4KG4QZ409W
vE6eiDkxxWckRPXCm1Jz9HUczWUqtrxY0g0f3G7QyM1AQIr1JKzJwNVOfWBcFZ9y
7cEdfqE8oor9SlEGXe1MunZEfQiH3Y3KHcmcUbBkEGIqNBzA2T0sZGbm+B8K/830
XrQc8thTPByqEkDsKZMhjaRJxEbs9xcTPI13fBUyn5XJV0QQ3g2CIweDiAeS7CEo
q9ob0pv/a5IZhO7RzjQbzFbqKOjiutloxOLsICXhQZKtrUOEaEiQ9qjZyLQi0Bw1
ZWrZgaInplNpXU1K14tCplX55PNPiEZGTVtkzYGL8WlwEuuco/WI9HsGpL0mGhBP
9vauS9CXEatmZJl3iGXEMqcmAbsPARPRtOlQD77geAouzpnGF+S0FjV+LD8/uf6N
Zii5Dg8b+63/2urexWZdDlLJOhLjtDzhf92wcPbt+AfLqZ/uwshQS7/ekfsX7v8Q
fvGXCaCoI58mAbB7yqY6xw41cAwHAfarsw8iOUfZqFPkyPMuRaXjm2GGOcHTWMLs
awtSGRrwVlAqN8TaMdyo/bliLNntrIcWNF1/Zvod90DwH+eOFjvRfwp/nh/P/zKd
5MoH7s3MYc2wcgxT+jIaGXhudXv2Lf5t10jqOdEw6W8KMIFNonucYyD1RgOjB/Ae
WC5EYOzFG+8dVwYdFjGcVU6yS6tFOzH/4Wet+7RnmQXzS63G3OhIdVrjE/raBWJZ
rbeyifoNHEGy8CZHjJzaXbH4O0oram/xoeGiAmYpdKKfOlLZhLhJS5M+K+hR0HIX
9FuYDoMy4wHleN4OKcZusk2aKlgk4r2MiSEFDETpqk2kHTT/goSSMKIN/mDISuGN
faQPcaj01q0l02XSp2xoML2hhDKF+BWKvtUv8p4NIbnPZzO+2Bq0rvOGcDf6Aq0I
+cvXjTfSfabMl0xUfsXrtKXRLsy58gZng6DobgHa8OrZy4VDaBVViRzKuavWG9LM
Ebmt34NGpeUHWbfcglVgrRUB5RZmaWkPucTE9mX2TyCztsz5psGssFueugJ7ZQhU
kbL0clPrAjNUVsgncmyr3J5Og0dBEuQRvUpio75F0ZSNYtcNU/pJbIDJMyacZD6C
38EemCagp+w2ZiwOCoLT9kFrJxJkRT+pOYJeqRuyq36CR7g3K/1XExCgwS2jAvFZ
LhXolGYt62pLomet82S6nWkFanchBVPiK5FfDXtZAY8yfSJ/Q4s8dA+/M7SHkCEe
iyBCglRflCP2QvpK6bGhAZUNHMZbEZOV7UZM+Zzkok049y6s8h21ZUA0b/llGY8N
IHvfrGLoPSOw0QQz3/Ojf0QYtkpob7j+djeUmSpVdE7pOaK4YysMru0Txrpmi09A
V5NgFaSRC4/f55wzUx5xwX9Vt0/VsPUgv9sIY+yQWGI8oGhGF2d1AwnHTrUro+Fu
1+TLCx5xvQpOFZ/u9BfF+bvZA/uyJTWzYhkv1+xUfU/+L/gP8CCniXkqVvCtWKjZ
RJKK3tz9+QK5vbWwshUJrPyXNRriYnLEs7TEg9EI1J9TbCvqIu9uBGTSlO84wTm6
C5AnjHG1WO03injreMtX8ShYLi8igUwdeOkrJKd0lFwxkgOSFx0PBVlwQlaa3GOp
imwQxrAcZlO0N1G36c88ShQziBMcIVs8GuU39m/eo+HcQp4GNyTw7JVTYPKuL7eT
XeWJ+0A3JE3/bIvMqw/QNtg/FgS/4s98ELAli8bCl6c8O2tSiHU9JCWYCthPZ3Ny
NsfO6zg8W0cWXnSDoH9X1D+7IvSyvvdIguXbmscDzd+yPrw722Q5dpHFXlwPJ1Ne
fWGDAhj3uU4g1gnRio8tkbyZ5celGbwSbiSjm3FowvBPx+DJMqURPZ/ME7KVS6oD
picHoESEXPj4csb284JwaQnmrptccS65lnQ7fsdV1n8ZgR8KLQRkUuAyPEh2wmg4
HYFSat5W5Oh2a+M0Yoaai+JpZUmz9qJAkyOaq/Dm359yDirvVUVeQOdarW5OgTZg
8CqYBqUNcoZlnAqeNtsOFzH7HFD/qtAl15qawfThxSIv2n1bhnirgyLhQ6dj2rBc
St8tLOeZf1j+NaT39bJsHX4b0IsMHmlmJ8RHpbPU6QgtvA9qvt8T768lCLOQv4y3
jgjW+rQX5UYAyjfpb1zcgyWJ63SXry4o7gjnoB0/XIcON8ZifHiUWUfIlNY95Og5
Hd6AWsFqWaEwEUljwlwF7P+gvJHxBiPx4tZI/ZswuOO2AN+GSDxTrAkIaI9/NSxl
KOcIj3wOGofBXNdQan8kInE6Sn/MLbBa1c5qvJy6ueWAN39OGICXm3hRY313Wz42
G8I7syCpUrsHFO6yNza8uw==
`protect END_PROTECTED
