`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
73MDwbMTd4lB7XR8j53ZzVyQufuyPyVA8J+RJOwncTCmkE47oh1pcdHrvYzLKlOn
xPPnfbEQ0wAt61OVZ0m7lselClplY19Fhlxy6wKEfApFFGHNlPvL8MsdWyXn4lbF
Sz6dRQvRKmic/gushY7rxFZSSv5vPZiyQaXHkfaggUM=
`protect END_PROTECTED
