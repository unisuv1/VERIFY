`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iyCsFBWU5FhgmyJQBly0CnvBaLlzp70ILhMoILrdIMuMNTt4z7EuQjOO3Yc/USH6
9RfohOY5RS7vZ3QmcdkCoPl5uAUpUbZ9/5DXA4/9fKh/ZqQYWw9V2KsVLfy3DItf
qLcuKYPO9xD81NcCpLQTBOXZbbH9ducXIsHG5ofnlSIoXRGPWj60HW4Ijdq5gOYk
6BZUjE7CBH1QMJIY9UBPrCs85t5ybcc0dH1EtPgPUYj9zVOlBykvJVTvutYfY5ZL
41OCGx4PhqCzLaagYY8Tb2VL1r8hLXkCJgQ21XZ2yilfl9Uzyg9jgkJNoRWMJg9+
lcs8O/xmmwWfa9j6VI2r8woN8bvcJQFNkzVVQo2GeNLrIMKb1tjeW3enEsnzWfVG
N68zZ+jhalkkhJl+vBZAJ+h3rqYHDpMsoiYA1ywwU2QBnYELEipQc2crTvEaYEqi
qQwrzCBn8TA7s5A+D+7HkK8FimCZs/i38cdlSOZskWG+8bBmV0a1xCcuYAfr4Pns
zsdue26UitGoEcGUAfWJNM6+4+7WsbRQ804zLuStRxm1E+fnmunw4DzhST1LBVAB
2bOP6JxRhEsrouNmQ+8Wrkg+i6byuUmm/mNQ+jgcf7P+1uckmCALetIQEqQpOii7
89a/Zf21dU2sj2+roEGT2u0prrGlmXAp7qCouzxmielseEX69aigLK+a2ZSVimgy
q3lLp7Q4C0T1tRjSMO0ohhF4JefKLywQv/6a+Q21cXjjaCxICxemUQrzTuexFC9V
ZWqFsH9DeYTvpbTlGCs/oYYm3YbVasGGfA4PA3pwfW6jfEACXkvGRGJXXLeC1Ap9
V08mq3zozZHTKKIbw3uXjZH8lEYj9D/4SxK4h0UlY7AjzFU4qVdUNzL4DlJJDs1p
IUNOI3m3hjdMQyESSCAX3LTAyA2XNwkeymMAnrL6FXN8Zqwsttiq2bhtD3BbeXHN
rk90wzpaY20tXSBUptdTc4cJcMr1CWQk2Cb+aZ+pWrhXa+d9zbZ1milp7r6dEDYs
hz4wnPUMzMC339zkadA4jywOBn014cwE6Qdvi0kb2pDwIf3IAsL/PFhwKLiGuTNy
LtVS5lPjlZpFqVnI7z8ypchzE/3kJ4STzOBaXm8GSPzK/YsIoEcc6x43qVhoyiSj
hODhmsYoosb6U8PFE4jLWl6KdJWLOktvth57lGIFcJ9V7JdRpldlOhg/7UgW6awY
YlMloqPODv6zA2knJGBhVTWsrptdUdfS17ph7BZKS0srBaOVbjXX4oHSLK2M90g9
rlV/V5AppruOI2fmBnqlLAWjbsMZceUHNonUE3ohULLw0HUBNUy2Ox2Il5Bf2Tp0
Z9htte1PyhjQyAw25Gyu2MiVKQ0J9WVP9EhPKDtOv0GFPZpGIshqn3DIcYIJKGyt
qmYYslzYIfjnf4h96lTtxcsj96u9QgnGsm8t/rboWqlX2Yqcnrg/UN03dtXsdOVj
45HuQMUMA8eJG9at0KWsMIopHpCcfn9uoQrlqfY4IRERIbsz/j5CVYFb6EDghs+m
FGbY2bGCUI4Ds/x1ilqgmvjrqNlN5wUk9cZKcyfOayE8StRT9BJrl++Qf2KCR4r9
NsXQcM/lfXLxMm7jBSNfqhKrLJUMWN1d2jP6n3z+cDRJn9c95ShW0xYZ/7PckyqS
rLQ5YXQLbZumJ8APWTiHB1xNx8aAJPLK9TNYn8pG4/ZH1UpEVnTkCPurgBcnnzyp
kog0XE1+1QPFL0Fxu0MDufd5N3ZgY+xAL6iNysScTNHpc1nAeysda99OBOkjJ+Fk
DdQkO+iDFoN3itWbNci8QJaDcoDennsW1JLSeuJAK6CxGi7i8W6e3LS4oSej2ki1
btkz0RBfx9hWPdsYXHrB9FpjntAoJbFomU4fKzdyuguvQM8s64GwpDbFb6DHFlPv
fMAgySPhWDvfmG6OS45y8fOAEuNgYEU+T1DFe65xQDzguKRDj/TZLWTVfO2HYo+y
366/z5vsxQvQyk5D5/SnTazQe8VdjlOGqeDAnByDjiBvTCzpawkCs6/oe1Y5L8mY
Zh6w/6QBa/1sRF1olzj7b9O3jwgzTTeoogmN1qbkvFhmxFgmJYsxqE8vtraYpnIH
ETIpw9K2Y3tzoiRB8E/jq+2Jd34+sIrGGCnCjyAeSaDnhu0kMlEytbnYjgX1xtHi
8EM5h93zlZHflPmkggVaLzBCnG9x9Z+QnA4Wchv8CSDSgEkhkrj41H0xT/+U06Eb
Pcp3X64u6xwsXMoUNaHaaRx8MC7FWgdTvYrZjPfmQ58L1twrSXgXT7pszfOM0/3k
7Dr/C8bUd1FDkgJXjamOpJrz7UlpIxUgL7kjR7rC74Sz2VFFkXOnaNWE21vKyGGb
e+iAXvSqD8Mdjj9oUgZ3Nq+yc4+Khp0mS/5uAP19EMzBu3rCFTGcKTVoNa7Zq3sB
MfkZ3MFkUVM1UaH0monEXtaRp6vm3kRReNoJQvz1VlmopxdmZRRLRBb/QHJuEOa4
vUI4OgPvQQ2AbC34SzEmQjxeTOOEq2BUHFpcvjlsIqXW6XKYm/xmoQtac92oPhvX
in4OEg9xcYQesFaMWXf5JqpHSKpmXdSCn0mjYtsQcwaME1Ms5jeC9X3SmG1Hjsa7
2tMyecP6BeKpBt15bTdzRfE47GOgz4TcKfbvYMLXE9YI2sOvBaS7zio2/shdZfVh
QmQTyNaLz9+MqBQdE0O/NrmrSbMg7iqE18dKCRFJ4mldCwW3I6VMPI50wfHwHp4c
y7WDiaxCutxzL86TTE3ABvDZTqZ7nI05RDedI8V+bgCukFO4GR40EKFpI5ITHmng
KAy2XRnD0VXxskVMU4ynVcE6q+CZ9syIaWJdHOjjesuuiwKj/zJ51MAZTF6TFbMI
9u9BflUw6H0KAcRkFzlJwiLHO9uRUhCkZl20GOC1Rdu7TnZOH8bFKbOS9e+ixFu8
fAugqCyDb6Dz4dO3pdc+BZPNj+iFzE07jz3/HaC+1HfJLElapm8Pkj2veO9y2CID
uWMuuM/ANvilqfHzo4RS2iKKUYO/R6hZdfnSAs7TGUm6vKSmh8UKmn5yJB+lrIdO
26woUg9MojIG37QqDjZ3UjCiNSjcusX3qavZ33BQBgERxxH6EqpxcM+ecIGKWzzj
wsdke7H+lIH9HCHC0ELW8njAAoqY5D0/UjkCGpeyUa8L6dEYPaDVXyEvcdBcAIbp
jx6XtsM3FioU4TKQ2v0EJvI59TEayepc4DfEy5euRTnkEVRcn8M70YPjtaEF3dPU
7LT4bv2K7rdcBn3UldzTuWZvoQobHKIhqIKOmoY+ZABtoIeu+tS6XItBaY6dUfrl
a+drxlxjD4bO/vXAq+CIYO5ugLuFfFXAnGp1Epi539U1lU+LnAJhl4XcYYccMSsg
B8p8nc3pocEcYVkEf+h3XgYfYj6Jg1U+C0sRIoTgb67Wtz0em82ZHFxRslYPjye5
IrjDPAF37lVTjBK9mZoVQZFWQbwLsqBcyHrJ36dFJZQK1OseXPegMICpajewJSq2
eJ0hPZECPIVp/BSPsbnY2fjSvD8r0imbWvC8sWVlWK/UdXNWLnL+2lzHUO9b7tOS
v1s8uFcqCrXfMiQ09G1UXqM4AbDHnyehchO/kxXCO8+ttrDf4Q48jm7mZYZiRhZZ
MYfa3tZHXJe/gQ+sC62fbg==
`protect END_PROTECTED
