`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8yQDMneBFZcnQFLvY2fmR62pACt0FnozxFyQIY3WBXQd/4HrMXEW6kxonIoQV1Bc
c+J3GOvAAQkTaH2ZfNRtuDKKM5yVQsYy6X2jkZbM80tRXj5swEQv30ka8KLROgHk
xKigb2umKnnWAOmdQExmgPVNlTybaJnXl7fbXFsMlzGjK0r//DEqIIBJor0OXpHA
+mQZPf5LV/GaseL7OekIA8eGH79ZOcdtS/8+whHtcJcTapSkzvso83wWOUwyJxWk
rcPAvmQcJ/p7v/wVTZF1XidzZwNI8d9iKQtpR8lfmAktRrWsjdYRewbh7TQIW+ZA
lCnnn7xLvh5TevbQCPdi9z0Oqq9BK1GFaRo1YaWeZT2nSkfRay1EKiON5D1GtcfK
6o9tnlTXibffXCeZmqAdAlrm7sBYSxXXQppge3MjkFZRXcI6xBNI1ERzVSKz4oBW
`protect END_PROTECTED
