`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
h/hQIibt+pby6lMSxcaHEO2of1w8f3zrGBqKAXvO9MWDHBMzrqMOa992lSh+rDKb
AG5PuKKRCkQ+gPGjciIwrA9RNaEt7DCPCj3zs17LueV8X0TftwyzYEFAg9ViSA3O
VI0qRgA4XooXiFMZOU1BWNsNlGronLPCJ064O0NB24CTMeBxfopsHMdjhNDDOqGP
Av0DmcBuak0Zw2JHnaPlUdjtOmb3m9RezL7386QPbToR06akoBVHr7IEihB0ljVG
j/j2gdU1qJuNMET/ctlDms1vWds/SyYFHMTW1Bx4Sgv+Pn5tNG2nWbFfAJG8WlcP
r9aTXdyLsVhJ406f9wMcyKoPufyz7r1cmuZolwPawKth1lSHfD6lp30d7awdE6xI
1kPi4GRDMnA6U2G2QER0ZuKrveSIYoIpEnrdVjhcOrCxE4OBQs/xR16Mwp91mPpc
KAbXhHKoo2UqN0ZJKGzxRP6x1QY+k2JDpwsKPTBrA3vhEhM3Jrh+23jEJ951+RgN
/iMpsh2zjk76Q2DMyC0penSuLGXZy0LY762FnVAHQMxpWSmb5mJvqV0VN66ZikkL
9+TrRpQlECduwe3kNKFuMO9Y/jaxImeVoQFneMoGF6D2NxFL9QHT+AkGJHnjYr4T
gfz/oo2rP0In9GkhXHmeZIVMoEsxwFSEiEQRJSpufiUoIvM7YeVw1CL6iVfJgqhY
iV9kKbdlwpYEzxexRdQKQRnUqYCGFaI9NZVc9NFOcjzM8zv/DPBM3hL5vIvmqErA
r6NqsAWLZNFyXifdRDfifGdK1esHk/6KekF5aXAhzRIFrjDhagQc7KVPyhzpqH9Q
0sgUTsSj0UEKYThkMOGd4thj6GqM/6bFLcBV//HPVHxgU3llTKRqvqWBgUy2O5Zy
FEAKzFevi9K+xRA3PqE64h3YJf776Fu4Wurj2YmjjEWNBRBKGBHX9VSUn4W0Tv/p
93lDmmdxAloQH5dSfFqj8SuekPSO0z5PI3uABxEQugMkTSwJ83reP49xaqHXy2pG
oesEcm3iaLV9I8eqpAGJO2iIQft5WX/N2dZeT+iFhxuOKQ5n6Puz0WBULdKU0C1q
MnyDim6+LIrPybLja3OOk10fuEqirJw4GFdcqmQSd8xM0QE0YlVi8ApP1x2CY3Ls
VnkFb1FKj5FH64R9OOmk8uF6FhFXvp/uS+KLChB3LfKu/VTgtS7/MQ/KT5Th0nBf
sAeIg8Q3iXD4SK+f1PRrTtvwUXxcDkB8vuh0dM+t7ZsjUMabjSieaMYQ0AxZFH5P
KBswFLvmpSGQPt70zcOD+BzJQOK1OR+quBGPbEAntZh8arogtbQJa1M8hbhqrlG9
hV9N327OSjdHPbBOMXJRaaQ/uxbk+QgFdnPij+Kz0ynXNCJpcfeGz3cVeHPYt3ea
qSA4bz/X1IrJCqN39NA6HleM9abF+n7lRqZgmhS/h7xqVSLA9i41fOiKAcy+Od39
MknDiy4NRzNwQTqFkhTHe79OW/wSMx6Na5JPwP1gTgjZLDwJTTSTSpwSB3BsAhVb
QvDyJHywD07caEgsC3NpoxkH7tq3PYJd0zVrMN/BkKJsO/H9CFBhHjlJFBMrl2X6
pvvZpBJK3GD7vsfTVhU5xyoaRUh7ut/KvrmumIbMSdn4bHJCwcPZe3I0MdPzGBre
TLdL0wqN8D3hfpa6O4XlP+dDYrUnVFR7UHl1qD2EBro=
`protect END_PROTECTED
