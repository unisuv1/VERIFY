`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HB0YnoslRAMJu21s3HpuR0WyNH/Ou6/DLeJkkfmDD01g05v2NQTWv6EoRcGe45Ui
LQxDmLAanKujpitXFh68gybTaO1oD/j6DPpr6TrmcY4LvgI72tYW1m/H0ZobLmWK
S+bU12jL3Y5IKuqnStaWBwIpijJMfRfssyDyvbNK2o3EaNBFdNzUKivzz+KTq3Gf
cecQvaTJHgmaviOUeAGCnJiluyEHnmS3Cgs+wTBgDSgBpamkVs3QClAKQ8agg0B2
Exr7oTR4ZGo3nEEnvlF6Gz/WJdb+Bo9ddSZ2jKMxnYKc8i41/f9mCWs5ZM5CsXKp
9nHSpDUFAOFVprgmF2ZrApyAjR2kLlYr/6tL9018JFciYcBvroQcTLyjvqunCBMF
qLgINDtbDGa3y7RCCP1KPcVw/PPtuhQpdgkFlOMJE/v3NRfycvfoDoIAsfHvbVq4
MiIJd3fnAtpiED/SCj5SkojvF5va+5D1r+5jLiN1BZEO6WWB1p9pTRIzsQwSCMXC
yOWvOm1n/tI7Fr/Lam96WI8bGH1ahc0VkQAfx4uodxRSji2Km8x4FpsgJxkbMsc/
6jzxH8oSVWz7jg6Q85/VsqZXJPSN9OpVzaLLjUWZhIA13mIloPJ8yn2RDf0W2jYW
X29vuT7HuNBdR7Deo1k1KxcS6i9RUmlCsVPPTY4/It1gyeaNoeCs8cOwfsRSLm6t
1oyBPDXvaNFMWsNAbuX/mcv/bIA4zKNC8xjIsVeO/kMauG0bWnHf6BFJz25PihCd
ehUdhpxcqKUzzj2vpIxUT0Buqqu4mTqxKjUuWg7WkyK888nbsgEjua9Zv4Oh01Na
OwTIQ/zYEZN7I1T4ivzCYrtV9tCclCAHmjuQKSdLXqfBjlHhNpIU6sM0NNpgXjm0
3AeG/b4p/s/lTtXR37QlK1KJPaOElPW8t1SQnhSNLdGkvVcgWR/5o/C4b/ooYBo5
ea33h2sgL3M6XGrUdUhdUXg4AEduSbwp5Aqs+HmNWL7Zynfb2vUnren+QziGQ0iW
QxGkFyiC7c+g9gsr5dN+dm7tf5E9hk2JlLF1niIwCKYvYZnOFW0nHkSPrlZLgfWV
ve3xojNMFbaojRByxarYdKApQV83wQAvhHtpyWtS+Re1pXELoIyLmTAbIibMzGvG
e1zopRViv3359+c+nujA9s2aTxjiFxWBBKOJ8lai4Qqxa+HJxwQbe+qs3Cx/SGg6
379YB5wtxFTmdvTwUbrVe0aRKpYLe1R+rQoKfDI9wAgCCzQI1Ggj4LTzr1xD5+Bh
1ItvnkIbcFpEuiOgQfwNM+r1d1Fde/rwbYUs57joSEHTmKIvKoYeX5g3R3tLwkVw
35UPLUq/lr9julxWjm1JYGaPMy+VaJm8ciwOx1u6Pi/JQkoaill5m3/5jt0Y6uKT
GFwRR/y6JMeH1bIILB03UkWLX1u5M0pd696m9eZbEt6Q4t4hmciruOgBLdcbBLe2
/tgu1HzWuCveMJ8qphWwNllm60ui8CNkF6RATxxID513hYrqHIn8h/ZxDjvkSYMf
vLd4nLXxcgcKHKNnWVLG2V1RigeDXo/JX0LWU+89f4Fpi90gwmQofCt/kB5Kkp1i
+hiK/hcyyBNzz2rdAaLi0bR2xMucS7dv5INdLaF8WmYgrq0TJppBlnamlFliMgKW
cPMIb7h1BXKFKbX5uF3w656RAGG4kM8K4P0YyOv+dRVgwdm0Z48/iak0FMH3pwzE
qtueLgqGPOB61fEX9I8+eZPej5y1vnxwMflNKaz2ZDjKD3DnTcV729gnpuPFDmmL
GdasHp+8zD6tHVQFdnVieInjxRhJQb39i+FNGMsgUliI8BM4XBHAOy60TQzDHkeW
j5vNJnfaxiG8cH79Oj4KGO/CUpiZITgTJsqvjXKdEtWABdPoD0AmzfkWInIRqA4L
vt3Be7WjZRZhkavc6Nb/VudtgUSuSdQWXPzWo9zDISP+nXiKFapg/O7qaWtp9136
ISCFfHhLDghyy018pGSPB36DhDT2etpC3kQhLhy74QifepyqZPgEWK5N7TnE5ep5
TXGQBJvOshj9MkJKJibEwZf2vWTWUCQKnHDZl6sANgiCU/70JsuMxFRHdWAi0zyg
YOL0TI0yqIYP2N3Z11jbdy1Jxp+dzP6vrcw9tub+VeBkZAEPAnwPv8o3U2lwsWqg
sAVrD6gFeHe8tGuEkNm+g6XYJQVf7QqCaIvitayRhowTudXemgMoDdHT7KR3HqA7
WSF2AEN9qOiMmVdSYtbgoil1cWfdI6iM+d1NxyDMH8Hh3JwocWceTTzvzvGOKhmp
cjLq0TtJi2A8TSmTZ2LAuzYiFKzZmGNvnqqHq58IeA1nDSLl974RGCZuoms6t7IL
PCKwX1s0jyde7BjpsC8oHuX4kQbkWcc3nBi82Y55h7zAsQQwBekT/lurIe4gTcxv
F/IiwWEaPchNPqVVlCFyiQ1KzZ3MTv+xr59tANdwMzX7dB9PFR+zKd0Vj1UXrzed
9yDjo5VmKRIPX9IS3JTWbdsGwmg+KRbWNEs2Zj1W+NHPwMZSARAlRNFwmw3UZS/m
Lk5Cv4+Xdy5wh3IZsJaSYg0ZEU0rg2sk1aEHdu4ngIHLMbIaGSBaqXUuFVexdD1N
KVPjwsT3obXyclplQ4yQL27MvbvkToUkbcNCT6X5f5l9G8Dj23bQOHuSS/wepLk8
8cBENSdKYKUbd4kEpBXc8f9YsBP2/BUBk+jAvY1eMWNfobVlYMv+br3JQNz8taCY
6atiqJ2orbbk4w3RcjulUEBXYUBXIRZCr1VBG4axUxRMruZKjvkjNryAD7pDg60p
yyhEf+RrsxGOTPA3c9pWAj9AunEBD48/Q0aOxNlDMVlcRkG5kvKYydMTidjEcLS7
0vFuD7a8uODzvHjKs2Be/1FPKAzHktu6S56cOTPKdpjJMCBlX73t7rgwrVpqTXmp
iw51ZljJVPIplC+jzvj7Qo6qxALoMf3QhNW726b/RdjCt1kVJPi6IS6xrzY2ljXd
uxJFHPmdfhwAkTs00M3vUKYYTqN2SHw1xt9gL9fHbY+x2DtvTxYQuEBVEntt4NNW
87g7l+ZB9QTve5DfZ84Rl4xrp+cjhc57N5E7ldQmFwJCv/2xZCcisITcAonvsBGw
yTVryaBopF2g2SsBpRfR78UI2bMVKOwfb+lseKvppOdSVdoujJF8o+tZcAGTL+6N
gTEOQrRieK19NXIW8bIbiN8sdcndoclhXnXOmTg6kdFKo4FlY1GAqHHXSrbqkhpL
iNYvF41DxeRrFoB9WKrQNl8T3UDJUC+dO6VXjyxN9XUMTrVyMEhq39jdW5bRZNOF
TT4jdzFdtr0tTNysm4MAW//yIK4Li+NjYekZyjQboX6d1TfJu+AH9DBXo+bEhHFD
+PVowKp8mx11m+eadYCPFMi2HvRaazGowjEZdC/1yeA2Zosdx/2SvIK3H3ynUrKV
eoos7G0v7d+qa4qBK0llnjptmPuMWaTGvZHbNCBE7xKvlc7Q9284hlVmBIyqZwKi
zfkunSLh4Zmkuc1SGmGyKp6mkwS2DoyO+RREsIfo7OTkaW0N0HLz1KgsqNTeeP/3
wE3purpHjWB+K21EMyC47cKvVpqyVtTuBNGPB8JYgOSENSJ37/LPymzLq28O3dVz
KUHRZ/Dr+LZ5FLY0JnB1lcVrSLOqRKW7qoNErD8HkvYNTAnxQJKHzUWcwmHaUlFn
mxIcXYoa/GsxvTpW6oeuZFJ7NNNN4ZCfAPEHpfyd2d11vJJXWrcF4j3lwXY4DOGE
PBcU8jPZ3frHWEf2ldsKEae4Fi6LHOZYU4sAvJIvrv6EYVxIrw6RQperzZazuc6U
FB2vQZYuFbLc8/iQLyfmI3eyKxzzxghge0zy4ZYZCksWH5tIovurkAUKlGNS+NYg
h5YuNaBhIcCNcAH4DRnTusqaGdHvxekwu5ejMoyEOieU4dZydUUDiB0jLA3E0NoD
DoHkHehVqeN0MzdwgGWdidZgfto4/oQn144ZuZd9Po519YV29zrNVJl9LZEfA220
PJvuoKYaG1qXjgsYdSgqZS9qeDm5N/lCy6ZT1jYRNTOC3a2JkNPiNUP79XI6GWyX
m6JihQfeKHuLCCGa2eavMkw5ZaLZwWy9QFzr57/696Cd5r/CsjJOEHtQEtXnJhYU
W0a0QJqB5culaj3Sg/PDHbaW3AZ26tgpbNJ2sj0d3IZ9IASXdT2idFiPMbJgZ46p
l33f1k3ifhV2v64SjQAqAsAMPGuFSt1GGk+5YBmZWeJI6GVKUv9nAe2shEHbN5qL
Vk3XEcAF3imgEluV/6mF3lg8xrCw83K28E9zcQFwG1GPtT8MszR6EjvWSChn+7/V
xif3o5u45Wj7d0wy7gg79VHt+AJhgzIcA7t6Qn2Qlecr8020TEpTeff9o0hLvyY+
61RfqNYmYJLisBZZa7BxRgpzxwy4v39BMkp/xOTqxlj13sO8kvXjLg87bxD8fRn9
n0aiYlqldeDE0Q3i8iM3iEiYDm5qG77JDX6y6hafA4+VEzYCSauFpvIm7aJp+0+I
6sE0sAAFdZhTT+8TUefqv4TBLKAeUyH19tIbAjTjJYfa/pzrbKWUcraCpactpqrY
iS33SfslmAS8P9vAN8v5uopowCG844v/rPs5rV+YmSrxxzpKX7LNXKhM0emzraDp
KwfKsy3lCuvrBu4ACLOGc11ElCs7bYvcXxGe3zHJmhKvaV85lC1Kj6LvFid2OSbf
PsrvB7n+KeB0mhKKW6FavGg0jvJxAEozPzxalTmootHgUs9QXi3/qBua8eZnQ2Y3
3fyGsIAj0idrMXGXevGuXg8yRlIcJGEcXDtAst4wptUeCeDDXByk2g6TbJKtnDT3
zKiMBkIfD2KnfWPeJuK8AvhCEQNcXxUOw4IP8uIUOK5DBnjij1bgHMQSlzhGGkL6
NZv6KO/mbrgnd1VJtKe36RG3/mcfgLb3uYQe6BnBUo4fIqxSfTu9r+xT4/INZQj9
OuMty7Fwdx9+NaqQEbP/mDpZS8CqMvI/i05pYupEnFVRW/5arXBzZEUCc1WPAiCp
q5fkBZqB4VGs09F0n9BbqmFFy4oKk3Hh/OTPzr78ZkmSvhqZZ+VfP79e/ZDDa2tx
l0Tmlx0CiS7wVcno7pheKU+wNVy/8BKaDwo0ZK04+9nD/T3xouaQoUm7ZEeVf0/s
gJzQa44WgXTusFbMgSf2S3PAV+H1WrXEf0tNxSDyhgE4XH7AA6oNTZALH0mRjwtL
ZsHjJiL9Imh49vCWoaPBmQ6X9oinCKTMYtxTiX87y/DIdxiZK5U09gWV9EBJAnlB
iFcl/62E71Kse/tdwkVh/KZ6HtLFfT5Jitkrbp2H2RihoEY5512Mpy5QWhLwq2Iu
kCsoktulqb7tPGl4N6Of+ogD28wtOChB41bCCyPssDH1O2rpd9epaSr0w8X6Guxw
0Haoi0ICZ8Rbm1k3AxyhsGO2Py7dfe2mgN0QuVGK2gWgjcy/oh05h4SfTuylvth4
Q64UbFpTtT/RTDu1KvGA8c8ZZZANdul4fFSMFbOP5ranzT+4Wi4B9OlpKPCPB4t+
0DB84wVZziDOi8N5mLDC8X0bq0qZurEiDS5rf4M8G9NIRU1RwenF++tssSLGyJv3
1Xe1cCF1HKbmrSNK02cPjyrZWzdeXXICDi3gFGCJcG1w36mbE/lznQIMWamNKu7s
GvNmnJAvv5lqWFbjKxKqu7ySiTL5bSqlnTbeWyumWMc9kYgBnB1YdDO6u7+LDS+2
tAB1ODyP62LCmZWJCnS15F+A78gdqTddeLAqnxqQbAQ6TrQoelbfVRJsUAsyUR8+
yvl1buIi5rUfW6K+XJzrKPbP6CyDQb9Mb9DO+HBcJAmnRio1pmu+pmUAjmHoAwFO
p+3fuiKenZoCoyQhk4veX6W3+mCXSYNFJumGo1oefsVUjGy+zIUh4MS2Of8jR0hw
Gzuj41CXlrZLTYYXWNXVIU+q3IXo4FsyxW5snNxZVR927eqw9oE3YrN/MKwFzoNj
kvWmb7fHZvKDiiprTnpAOg2daE9E8QqsSJiha+kx2+fbQwXsEckxTml1up/FOCvo
CdtIKq8Xh/siHeD74kqHQmUrIClAR8v8dOjGy3J7XRXSIYNbJE1dharVjHaApYJW
wWafnuaEt+PLoEcNQVLwPUous59XSAj14I+fA3fxAcPUhCme7vf9NmYdqxTYLdzk
mj5r2vyuN9VTiU2aGXeAFLq5CvO/z7+zyeck4KHTQq65EpSAL5ODP5Z37uq+A3oE
rnPN/TONVNpmXGoMFeVBphR6VJai5rc0mCXo1/ePdsZmmzV9qunmm09vQvBUeF//
m3TmCDNDaKR0Cn+RLTW0r81sHPchyd1/xFapywkYU5yqwxPIm4VpYWD+z13ODqV4
+RbYGtjrI/dbxELIgzi1+KFzQQkBY07hNhFMOwNzoN/mR9OEoK3kM666/YeXmqrG
SXTuDysvdwAK219pqLLP8iKL4qGGlhyXoemlTfnPa7ufawwQ/1MmeGOr9ws3O64T
M1TTwOvVmMqrd+3YhhLlv/CFtpBd+wcEfBgwBzRfwzuRWRw1OHp/w6iMTAlcEAQW
L2C3eLpwkAuzDsefNcOiac9SmjNmuwIrfe7On/UvNtuDB4v5wmXTh/JU9lgsXL9z
0edlLXa3Z30RGCuoULsrJGfnb3Pb+XYZ8XdhT8t6hnv7U56fhPm63maPv+EKvU69
gjSaSDlVTkd0eNukcD6essm3uBS7R54ysrn9gCDHAvF7p5NSMBcGcyT2YfFtMRFi
XJ8RLFviDQ0czPFpbvLLTnh4k/V7ppZ6O4HY64ktht3gyEDegMEu26apY3Wp9fpl
yLstAYZljI6Gis6AuXlkaygPHAJ7Wp8GtDQLa3XJZz/taUCt+EppYb6ZLvKM5DLH
zdu+lXZYN5AxgpcTbAr2hWx9CldUPtN0cDO4XVtiN3JtuESwK1VwYxbI9x267J8a
954/j/3QkvIqOMULKGex1mOd8IM7Dz9Bi9t+T3qOsBe/YS8O/BITXtEdidSFhNIx
cVFR6MIFUf9C+y9eJXR10P46GVQyWBgoc/qU5FvrAn1ebwyCa8YovjqC1HQcxN23
8Jspqt/YsrtcQIMaWfcIw0yBYmvtrgH7XLykY9FRvDYV/yb1I9/0+2rzY7yuHegM
V4JApaHFr2PdpABLCSIKvRR7Ic8e0QHm5Q21JSS6CsccGkjTMQirIs2ExqSHhg2C
jC/2HkXKK0cMv2POvd50njQut5ISh+vb5haLtLpzcePnVWt7sX7/jtAyHZ8/43qy
hwK2wb8w+hIkx392lU4ZcVWyH2D4gjBKP0GMzO7ZcKG4HqNg+p6WsJHRZgll1I2y
8CY73AF7St92kRg49qeODfCVZPw5i/2BTK5EcjIr4xOkkWB5m6PHl7/zZwlUf9dn
kWZ3AvdasvKhw7BbKr9SrEaciYRSvXO4HnnIRF5OPi8a/WRrbs2PZ7Om1IHOXbmQ
NIwtw7y3O71KQQbihEssAOOwE2xLcRpB8WGSvUMI7bK531RGBYUix86TKhWxv5X1
BfzuOTRRlj1eca3bsNn61X+bDRdj41xuMtzXWorEwEs2KXBkAywMx3Jwcq+vYNrs
ATrH47B/8ShJs6h9L4jbjMHdXFQqWOfObL0TTdlc5a4+ZwLE1AIGMIDInbNeLNkw
kRh7M171Lbu0IywFvt2CeC/MjRpW+eLqP5g0H4lNMgwlzzt749y8EYn8TQzvZjD3
KgNUyzfP9/9Njg7CJvHRSpu7d7jV+fVwrM1EW8yetroVM4RBxPHbOC7Ukqxz+edw
tZuDIaHwEph3SEg375HRPaKlaGGCPSalgWyW1iHJ9pc70U1a3rAeFfhhRy01+yuj
Ph5RIzSu54Crf9rFtqDO8TX9ibniEUkgKjh9YW6t3HMKSznJ+UTUVN923v3s6qdx
YmIdfpFyLupWrT+IFO0Gg0fwMWKb74lSZ9cHCtFiRfbzIpM6bxOHt/hry92mac2r
P/OP1tnRFDs35vVhEALpoChuRQ/Y/xf3xbGh54InefBzR0UPDEBSrH6wjEgQ2IKI
9EJSAvAZPobJwI7uVOcyqWAh63GSW7Jx6437uEW0/QcmmwDcdLfcN+oyUNBa37Nl
tuvGqU9N/Q57KHj+wpjYv+FpdFU38usZvCdlVIYjLfQ0baBNz3EAVm0nfQa7ZLdZ
MtbGwr8S1rC6GQmJf0tdoAr7fxClVBZjUVie40znNh7WEa6WtOg9uiciv5C3yro8
wqY358ZcMcEsTihEujKb3dOriJVKDj/drcSeWQyoKG63RmQnr6cJYzPWXF7rNCkX
wZfBYzEAk6+y/GeSX4T+iBMVyCvbiDadYgKbmrmlEKbwNIJqahLNpEmlC7/M6WD+
tWd4M5Kg+o453Y0zzjNerHa7s0SJ5jMAcAaLF9YmzZGIYAswPTKTdh7+RB7EGLJn
ysA8EPhv4SsKOdL/TBtKo+5D2jxOPMvADok+PueRMpGFtIxoqYVMQf9AxoCiFrKR
a7IOyp/+h+wsUV0xFl1GhTz6uR0mdCjyPGXcXTPCbyV3QqIduhl1rPgZWxj/kBnX
twcdWjiV7lYAPh9VLLHNesiToDdLcljKe+k2htGh2G3mhJ9Z2F9CwcEa8EKIZr0K
7O/UlHY2y+YjLztDrkbYwvTarXryEkVm/qPzRoyge0Pt/ddFddVGVnP+zEf4zcyh
UU3BK0tQuX5iCqbty5UesqIZ6zYOSiEubcmfOmqtXwrlvWEX2axRjHagvWhfH8YG
NgaMwpjtqLQ39xrTtauaCDHTTB+b3gUN+3sZq/RarJEZrObDYkHSPBKrxsSK68QW
6qFxOjMI22PicaXfkauZmV8KjN73hFy0k7yrYP7PfhxPgzMGwnRC2YmhZoxiAp6W
dL1ZzsFzVh8E1ZUdhCPgcDeDC1uA1wLNxK1G/LYZCaMUUO6P+RZ8WLXYio2DmOms
6GduBRrsFgw6hPCWyttfJ3mQbVL9a3iV6tGPQajNnMCMUambmSJyeUoi5OdNZF0C
ctZmt8ZmdbUems7NEHsJDCad+FqTB0kwi90OujL47EszJQcSObOpyMMOhSNyzz77
WpEel5Omq9aGmZeNjeSeSoGkeMyHMpaJ+pPV+376XuhRCS0JMHVjhZ+shMkXT/kh
L7EsWZCE9u4LWLX6CSYoQNwfZcd/+N1xlHh/kftvXhZRqjCUIk4ivKTVI/EV8frN
xxLzgFErOLKxYYoa/TtrHC5tRlA8nryRKz3fawLLFkvdDu2AIo1eneSAtoOdIUQP
bWN27e1aSWJxeAWOWaTOdY6l1qUqLyZVKEiSiYUl3HXXy2Sx2KLe/5vgwoUO4ka8
EsD70xUi9VhsJslAfF6jyrFZL6OjAChG9lNkwAurf4es3DtIzAf5krbpT2NJb2x8
sFLcQqp9Fr6bsWduRy7H+cGIbQcuSrlCrju7EtGY9ID9Ol6TKc/t8GVbmURwRw4M
1QYIm+irDD7StjvZP8k/GJw5hDBFClzzDNnWqK/RJUTP3RjWnFxgbYbBVzsZVfAW
h5qKn75/X2UzWIfOEOvoUA7F/6SQiPrMVJjTEKiyGh0r1Q/rpH9UqTu8WMGVMXcJ
zXWA81Yenvg50QzBmi3a9A6TbcuHtj3rIcogcatjGVN49MosBEN59vDihoDyf/c4
YbxYgYhXGH0oQNNSedmU/y2N5SFi3rSf+lUE0McShVCNlvUGdZN78jfsWSyJfBO9
LtQqxozkkhhJhT65PoDkKf5EXH4kCl3KmHus/VAy3of+P6hEkztmDYdosryTPaxo
EPBc+WL/DAGUSRZsxggGWzZ07L4xYWynY3QfhYv5zYetLZdbAZS6IgUVCdnJ2Zv3
hlEbK8tbqTscKqh0iPGVNOQnmiQqFq/olWtp2roSXY1Vx53szO/vHKJHk9kOe3I3
oD9uXx6Lb0AjyDzyamkI9p7UjHpZ2CPYokhEhR56+Onq+oQaHPiMOUxr69v8/db2
px1ts0wrGC1J7/eK9so8O3/ghRtHSZsPXI9lSXVJC98s1JiFDxsVxFphLeP4UHCU
eaDGqVgSKD9SeZOr8CN31pZEQcSe42Tid53h68lXPZXn0jH8OMfm7zH/x2ekNPUi
+pcjpFZwZj7Qpx3xxFJQPnEiDpl0OBP0St0S8DpJYneZ2WO4JIPiQOB/Bt5eOq5P
AfC90J0DyLcgCB19oU0F3DKmwfrCu0Alycx6E2e4WybAoyDiUiuGWm5ZqQ0kbgX5
T2cZOFBiQOp5F8zUKpHPj/nTaTp7SYJrblgozHnY4HPnkmGBrb1PgKh6gw56jX0/
tnWwD+Lee4NZsvg1bSWOD4N1TqGPRpzxhPWTkyZPwOBAR+0T6c/GPPeegOlmYOhL
Od2qRnQZ395BIhPSWqz5ynG9QrbwL5srNKU0282jij3HTqUMG/ngumxX4dCblyiK
zpbgA7WwOKgen3+cj1B3jZJ9Q3Oj7eqmqpRu6Mz0vz4GmTVNHX66UOBURRbGCNGr
UIl63KucwxegEcZSuo7uvfvaLcmqXHi0C0iNrVPL33/xnLYd/dU0tQj/SYFdatkD
+8+2LimMAlgOyZXrfCW/ognqrpvi8uyNz4eFiZ6bYCM8lVP3AUAAUdiaM3xPnYbf
iGlzdOIIVl9LSpmwCWtJp8ExKMSpFwUyNh3Smmyf1NaayH2ORV6CvcENmtDK9e80
ELrtnr46CMtAI3wTxc3RSKe4nr2a1u6pgbL5GT+u9+AH7jm/2va2TuiIIpFvEa9O
EHnXVjJn0UIo9002B8nRmcdpUNN70M5DS/ABNUFTuW4RWfHlzY8TTv8C+Au1+ah2
+Epj6LjnhVKL9rv3kQUmvtufZ2o7VB8Nw3nfMF1af2M10AgbjdXkte8wl1QuRN77
CsBmFfUziPWNa6GZMCkbpQJ7kOVWl4dS9VbfCcTpdrc90tC6H08qmoB5A6tUNT0h
xt/lFrLvxeecV1kkKEqqrN+2MuEnrkDideXS6p9wxc2Sml6vFUhXme0uH49x83lX
QW/gx5VwdqYu2LTrjH/BtHlRD7v/X2hrZc4cDL3S9mcgrRCaH5uW5sw+GaRisKKb
nRtPl15K/GA2k9Bou5tr95pwzQDJIQRMxNmAiYuu4lv/1lTHal0ExrQJ2MRVirMB
hFCbwDrjx7RXww/2KNO6UPw/WpsAPvj+PaqHoXutt3JxVmu3RhAasOg3w8eVZZZl
3hP+qudaLtgEyeCFXIVchA5Bk/Cu1929wbFnltEBHtNBcdOhxhhWBoB83H4XKkDq
sZvuFQfdL5fV8TwiJZsBv00l29PbWZaSgOKlnKuRTMi+XEqfWkkFEAvKPBlhqSmm
0pQoZ/B+NoylBPsYjzX4CofKD8fMr0wxXIAVwOTh6SyRoqAZHHl9GzcREOap2Qbq
YReRcOmJJ+jI7R1TPCi7DAecP2qi52PwcMOiZIgqlUsySgR5dSGWlzFL295um/3A
46ptwmoTXyIDEElYMUnir1eug68NyBfREd+Pa5eUk/aRGBrZYEgD8BaHXaKTEoTF
D0cxSHxi1mBtabBPt14kk0iclArZHbltw0bNTObkq1uAo28Ei6Pb9jpGvIW6k9hd
hWxRzTXtb2asBIo7oq1o3tXfDgTdG81EKaSRyqLUaE4YICM4tKt1p7E5F1l9yhFy
WxNSOFi0glrOfCbghsLR7gArVafC+ibT5oce6DlO4gWYTtIDFZE2YHrJHlPgNhAv
y/o3itdSZgDDPogtBMsc1lh8pkVcPzxijdHAaBipOqzfi3/g/ZuzSuZ8+BjnG9ev
PuavbfmJCQt1vtTZoOp7NuM6ou1lzJZ8vASZN5TjAafydIS5IisusIlkvmMOAg1e
JYXUWbJHEFxl5ISHhylNGRHF3RWemj4f3uYYdfmLO7OCNZA/LDWbBOMslZcmJ4lb
S5ShXfIFFWZR2Gp2cTxA0uXIpE2KipU9UL3TVVe3K7XBDPe1exefW5R1tw+Zx8NS
2ZhXHAClZvzHz9ySSqfaXNHqmzdQf03iOUbAU+ugback8T4nPHHaU8Jb2DYXu3C2
ZTlStArr7de5xHIdjfPy2DQiRsTg4YEL2TAdqzfaJTtPZXVaUxK5KvZLGaXT9Qbv
aKQxttbYbWMdOapZ7+6o9ZE6aDONznQSMpJZ8kZHMJEueAG0BjSgcf379LIautod
tEUuwc+qt4/7VBJ9L96r5taYKQzocIqV6OBTGpVIe7PUENeFhKaPKz8tSw1NfwWY
w46sNQ0/2nXB7cY2pPtZ3qAK/UePMWCmuEiJHoblDCQDz0/1z7vYlUDUrlr6/CG9
37l7Jy0tH2n2sEcaK18moZvRdXEGnf1JQgMK//2WVpRk30LQehouKOjoWF7FQ4hz
bklSInIi0rLh1dwHdx7uzVD6qSBVqEs28ZJhapP7Kw2TMRNYjAI6i+p9/W0QtcYR
aDtZarUqoLB63Mjs4y3v8sJn/pF+3VXTDASn7gnRLrI4ruWNZ3kNcGL0sG3GBA45
AbswFdMH5DBbMajIEGyCoiMWDI8aQ6r5DV/iOu+F4dmLfZ4bJDnR2rwAkOe1ySkl
SBfC+ZoQDk4O2rpFwDzRMZSL/WnrJpmBeMtpAODwnfiIE4Ci9D6NyS3Eanu/F7vT
Q8Jt6Q3OGppJzijYOC2EnVQ9+B+u+sCU/cA5DsunEjXPmKLBUjvTATkSXDCSGq9F
HNfiCcRkInXzpuxDpEecoC6cgIKWjfiEz/fpSLyciT07osypR9EFqg4d0Ao4nbem
tO04mccdvt3ChVgUMG6Qm90l3MXPxTGETkt4mp7p6Lhk5thUCEukt8kchnaOji6A
Eoz+MxA2CTiPJNiKnLP0i6wkCRDYYVxvmqVY7EA9KPEVIvBSnSeQeBxHF9ikJV8G
/Kpz28DQnldD+jdLgOX0SS8NNIhcCpCfKbMX0e36IfDWnQYzr3o7lu8zo5qwnp+H
fYIMhPo5qGdsPZHbgbKKGn9S6CLYrtora45iLH0qZ5vFcJqJVgaNpYUsGSt+KxPk
1MUjJPXCVAi1D0F5CInag7iZxjCyMjnW4pw+bM++wVvDKqWAKPm0T1+HwQkumNyb
Qj126Sol4bUk3dnA4iykxHCb78BqJM4XPwB9s3m+SccJ2Mw7So/iTaixFV5aTGz7
Q4esDBs1nUzPn8+GyX3M2SNXb2SZ0t8kyJ/QNHCiwpEg4RRGWkkAGtHU9mBhq57O
qchfx9MXU+JIiIQdwAWs78gg6FYmx/zu/BKm+ECubXeJxTb4vR60iv0PM/IkZtuD
4oI7R5dFt+QWO13pxZU8eiu9g/0gxedwMLLElyxc3F6kEueuU5Gq5ihc/VuAWXg7
uTokkqPwdqo/i5M/Cz0f2G+kiDdquQC0563Dj06V6wTpn6l24tMMmHTtBkUcnBMh
OVa+Y7mYaxMtvDEF1bgtA9/ALicaeEz5HKK2JvQgNx2MPxNefoae8yaMzsh/rc26
Lfz2b7bEEx22E4YWOldyzg2/Ax8BGxzssRdSGdsYX5oaP6SC0Zd6ArWJqPKlQnyG
RwhqzPd1dRgtz8yV+/UJJb5xaPDm1bbpk8PAI6zdLHnADwCRPJnJwJ4smo7bxmyB
yQgmC+U/7hAoBHS0DRjJPGo1Kye4mdGdDii3xUIcwzSJuKTXttd43NobKGKK53f4
1iMq1BWR+EgAzFwF75Vn3ZRB9rTfDL3eQFGk1vOf3hmFezBgXmONrqrOQHn/39Q4
th6SugHdEqQ0MHYwhkgTPXMHfL1s60Cg9mOULsCiYytERnFZGOl5yMEU5Xdp1vpX
O+sp1go8/xDHuCAaLVausD92t2aGtSwGiGGkZ2+xxtHsuMA6stf5WDB5fuOZd8bm
RaV41uGTSojUCuWHjqsS2N8f6wvUR+3ry79lVw43amKZO3W60j3RV499fQsrUTxE
t8AvoAvqrnwFNDo3HLdFJXF7aaILrQGv6DVSePYjCnA+YDKXH1ZzBqwDlJ9ruq97
+ff4m6GUFA3s9T17YfCxP+b5lIwOY+rHkuyaOZusMiILAk0b73lRq5IGNpk9Eilx
AUUYqXkjeb6JeFSNlVRxvc8A7GKTDEbWvMGLqB2bChG7Bi8k+lAPDXDZmGb0PRP4
1vjNjyFKGNFe/USAJFX7+yTnZ91fr2Kt2OZ3/nkFF8oLYJPu0B2aBc7ZF+4zWmOR
IfFrHM2ikgT2dN6NYdrya9/Ddab67Lh3STwQYkGL/wNiyjzUaPdPQC0+TthMGCmR
crK5gqnIW6W3lIMGG1oUIqSdqubtzSe/02hLavaNuxgj7j9JYw6pM14fFgoQW1zP
1YXdnIUMJYO5m7K3WUmF7lywjwMQ5TTMX0xDBfkBgiC8ADE1S1FMcZA16hqm41mx
4IyIaEilufBNuWJMdlOZU9PTPZNiW/9ju82LdYURWU0iae9MmDP7o0Rh9SZszCOP
UE3hnMBhyCy6EzAFAyXrmgisDnmGkj6lfrqHzo85FOWckn+G7C1dfqhJicFbHdU1
62QJPPC9zUA7HZE4baG214obgjeDxyxNyv0xGAUyD7sj9NvYS4VuLFeGBIp8+ln7
Y1N2s/a9kZIZxJnbu2LPeP3bDcGIqK1OBB3qvgZWePsphM4/tDXRoVcFkwFBCzNM
FUm4tW5B/l4d1vls8kFgg/2V+dFNSjUoPwD5SYEJFD7vboLKW/9FBZ2+Q6L+KyhF
yQeAQ+3ZVwSOIQcl4PccfJXeAOd6MLjkSwohOVz65c+swwJCnGFNhV3DME/FQaLh
gze3Cj5t/m8x4PfR6l3v0BOH8E9DLBJbJeS7Q3bHaNduurzztYaVZm9ZhQKrO0Ie
w5uYxY4r8BDjKEB0NS1hTafDwGB8f2lDqPM+mErxUAwbza9LMOW6gCwNmkoWCHan
NAeZu5LXKAQzxLA+qxi+NnZJTJPNzorWvkpJOCUgQJHUuaJaz6J6eYq7a12V5bHy
K0rxgrkYdayRy+m9KXiHPAG3iZlZIJPOQY5eWBnAURe+RhkA0wvye1RuQA2A8EnY
kj7m+ghrtivUjUs3o7PS6RkkpaBGRNh4r9YWlyXZdHwOJxT4ebSj0y3l52vP44PH
Rj3ZVmw9lo5fj8GW8IFByK9zLFZC5YeiJi2bIsj7bwVmuB8jqR4HMMt5eWL+CDXY
UMZJudtZbYVucoJSz8w7VuMK7WzYn+13jfYuS7Qfah+Jt+WzFikJQQviJm6XhbAV
iPsTK3nDOmt3Dv6XYqSae7LX+mBrkEwTn+asMewZ7ZJpVHPbgklezM9Sw0Ey1bCD
lzB8EQMPX50cFmr4+YOJYNZF9IbHoVWM40uimj2Im+eKFTzJxrY7B/rQtYX5fEmp
Rx2Ynie+kH9IVdvWD7ZymnM5vjihXYpKM0SkrNCKMwBKqnFGXABChyQuOmPMQODm
9bAisFEC0U0sry8QtQj27lSSut0r8s+jfF76qfyJDGBcmc6WEsUwjrRCFMRrc33U
R1wm3H26nGxtt4qh6fouCAw8MBBidSaB6/u61sTVx2PdAWtz8DkeMMN/D0HqJA82
oBSgMThaaUyibAA9dcCniLLEIcigUel5sM32q++efYIvBa4wmEDvKqhmqHsTmRaS
U/5iLGHI/pX5pRr0xem4jcMYfkGqwaNK+zs1nVbDS5IINAPZLrc/52xYTMu6GrXN
/rkfcn/T60FKwk5TzH1QHgcqo0ipbfHCsbCe96StwDOqecN2GdzPl/qWJxHhQM5L
HVJjx2HCBwdS51HT+Ta/GtnFR1heZtr7a62PZFHqq2yNjWbN8jur23rr3SEvl0tp
4l6YKe9Gul2hrkacknBWQ0VUdJOrc0dy9WB5cQr32g7grF+m+2jYyG4Rqg9nOxui
chk7r36aucQ7pjI6UIqaT0UX6Rlg9VmYGwU+Sy6MLtlOYqI645Ga1DcvNZeHuk7R
F7LKfGVXF53FR0dqoNKmye+FbZqA41UkKejVEq91L0R4KscfohWgKvtzt7jPJddV
JWQW2mPJRee66p0o+BPBzvmDTUNKR93flOe2Qw8+zoN8+VK4jTTHkuXBZtps2O/m
OfZQx+zUgONsveIchpsDwlxB4+f7/wI5kTbr2EpSWatG6zpnfTs5D9lp/uecrJat
CRpHyeZHMbwkDSK8zgXlYplbi8H3Ia245PhjF4pYSvOBkzJ7p3y0BSC+GAkjkxoO
vYH6DyZi2/1wSHUTW4QKFwV5cTiDoLHSf0imYc8fpUGUj9nmUqFitU/+D44DA8UC
RD3Q87+70ov4H1g4PXUA+f+UomXbTke7BC2NOpKnWyebrGVCvgIiO3HgHbbq+Z72
EggvXTgE0PQ0QyKuqVPmpXX365w2Yn4eXx9ATB4XWMx8QgknPYnimSeztYkBxJ+r
82tc5qFTXfkJYhUYNFlIff1R+/Lwr9foXxbgT1lBBu9wpblPBJlc9UZnAAChgOgq
mxdjIfkSpXIjf+hwKjLVLuk64r8dmD6lnyI45W2ijfxWtFD4HSXBWwXTrJ7IOdcj
5dLG9xZs2HBUJx/S4Cs0Eyu51zGD/Oc6QrdIoayKgCtBhc/p8wQGvHd3nzqy8+tR
KieNpq56o6NnCbIHI8ZFJ/4G5ol26heXYAurTb0VDGqzxtEc2p7iXoIoucNTp/RR
8fp6BfQWOQF2NpIoPZTzmbi0IUCmDl4+kPUgVCZIn+OYsIW03HFlcut1fjyf95Rm
ObDu1HKBpqPYpdXmP0SbviToE5mjOGzutcHhMTGl7A9BgVe0fViHDZssdbfD09Ib
vEZdaj4AjzCGzWYIjy584a7Cp3wEPih2taVry+t9dufhq4eWwF0VeyypacqBZA7O
66fEx7d0MIlhczZdESNZck3fNQXajtszuk3+/UdyYZ/njgcl7kVo8G9HBJtx9+oh
veuAmuLiiq9qfXqH5P8EaZJq8/V2a351QeAiI4UPmoem1tpH3xpAz0W9KFwTmQbL
O4MOwDxhouVJnJYAhXWzkPiVaKur1bK0RTUrCfNNDfezG5ikpp2X/CKsQGRfH/3T
6PtNH69/ByPHGMaTgwCiz7SrmtMw9/Y6467T5bbMMLVdmLRPb6dywYw+mp1CGGoX
37hJAvr7d615jVJAeEKvJk/bJDFIRBvvu+dhxOfBES5fsoQKy6NczRUvt0j7CrE2
q81RmylWx8k9mgqkX0wYHUurKNsG5SfYnFAXg47iMQA/X8yuMk1pQiKkQSBQN3ML
mF+WgMJ1zq9dwVrhrhdsSb/HraOmlV5+6fL7cmoVccbTZnaSvmVte9w2xu2SfI2M
XwGapjy61N5DoDaaP/AvtRNDPpq7KugdLtNedELVkKucHDB0/4h4PnK4Spb+dub8
eF4bfdsdo7f5GQx2Wprgtyhwy3BXC3H04ftts9qACJFl3Fw5R4Xm4k0FukkYXgSz
7AjugfwQ1x43FAYQA52IpwcOikqmK6c7kcWvwLGlzT+qp2AxmiPwB+8zU6E9mi3N
J58LKqNcYbmwF/tLpMXZz7mGx/leq6XiGderAMQf3y1G5iIfOfs7U+m8jGoiFL7X
sg7fULDFoSa22aYsOflQ4/p0LcdwrugwxdT32yUTWR8amShrvfXX3Tf8+VPGUfM7
vK/PfXM6QhQbOe3RFrg2LCddV46+RBy4e37B8MIe+ZE1RGG62x/ahtNkGC3eDXm2
yEz3DhX2jwzVDNOrCN+X66Ju04ps8mQ/R7UlpfbzqUlBhxMW0c7DlipRoi/vOVAn
76OZBZ5vkNIZwCNhw/8t9Q4uBCfwMGMx0buWrBkjwmLtu8t1YOS61RKbrrLA0fr/
CA7WNccxq1uzcrFzFy9jh+06kVdi9PsC9FUNc7vAVxIS3N2eAkCG8vrNzQtYwsW5
mUTFSoGFZxAzO4LjSpHHThefpKd3Fq5UApOPKQc4+Nkvqjg9u6N+NgV6EO/HPpjO
43o30VttoW4uNU82Dn5wnyGGz+ym0WHxudKETHEw7pNdkA6LHu4b6aAGoeyK+keT
vdUoZi0SbvPdBWyc94osoElyCbJsOOeGjKOIFckPpUMdJhGKnRV8GKrwDf2r3Z63
j1jKnjqu4akcH8eg9o3GHdcrASQN0eOeTDkluluYlMO63RNLCWrjMMhiCvHEq2pe
ndSpZPfi36T+neM+GuZpk8VqMG66mKEnoX8rtVYgytrOfWSYgZVqsOtDr1xv5ma7
ca/xipZ4TRNzSZ0n5pQKUl2JX2wZtaxYsFl2cbfHTS0ZQvR7sGdtbbdMea3lB0ft
bZnWHpzL7xnaJrFLUjt3GgA1Xu2OlO7bnbWMQzs0hXdReE63WRZh4kO7NoUCJtBU
RyoCsolAQDWrwzfS6Vdw81nu5ET9B2ynh8liczkzhOMdQ7d11y8xwWZlOctAjC8I
hp8s/WFLj+Qc4z6085nbLnp916lI+4kxKTSB9IZUt0qtByXLFCCDd1by3aH0h8Vl
AdnWbWEmqc38B6jzKot2AD75sK4dOjKDjD/eTor1KpHFi0iDBQwu4epSCnBdQJzH
oakp0Y3JTL9nL/6RAjeEUTKnBZF8WXABCffbwDuJZkS4TXOXJRiidA5NGWro2MGT
KXvATYWiID4tGH+vI43KVCC/dtw3XSWYlzg2a1oMGQm8NZTeO+DUnuAHN/cqEdaQ
eW8PvqPQ6DHGCXYB6MUTl97SuUSUXPYrb4GFeVhg1sEnut1gQWR88gKHr8Z7X9q2
nUGS8tbP3MWadrKseKgvK3uUAgtyExI7YsVGxk2XhAanC59HPu8b6TfRkE46x1Q0
+gm+o+NkTxIA10Ziw7ChHCTF/ljzUsM9X5FKkdsgyQH0S8zV9Ofd/To0rb9cEm0j
oylA4C2eUxIwPeKdvmpGGbvyiy8xtqcMgstz7K0r6LIT0HGTHS4kIqxVIazDCtxf
AAJPXpWqHrXQWqI07JMtabSz8efn4/b7/8X/rgbymZDo6vhJnjA0mTThhJBW6ZTN
ir8SeAwM6Nk5HZ+mPiss/JwGYW/zl6AdrBz3d37m+PflkCFzYvo4k4akuoohRcjD
BPUYOsylkWinqDuRgFjfiB9e39VdgcEolec4XSF52yRW47q+ca+1wtBsKi0MSdZL
L4acpk0Tzpm2yyqFYgNeM8I3U9mFSYkmsgxvXR4rEeiu00yo4YCTEPt992eFLFtU
0uYzfob8LJEpcXn5SX1sANzmcToS6IE8j78/mH9l+5jMGNBnAlcLS2LaugEtZ1nK
WnXTMmD6U3H5yAOAq3GdqGM29SBAFfDOADS0fbkovvIgNeMVq+ZmW5f4UzkCqu5P
5ntRQIL3laG3i+efwzzqVHiYc8WC2jAYVAFVPlB66rpsF2L3mCvzPTfGzavglXtG
+D4gw5rRq6yWvCuKYeH8bpuyZTAci8I4gg7i0Ralsgy2iR2bL4Kk+YCjoUVUjO7W
3oU8Pg3G9RqPFoMrbQfL+GNAqNmjOFCqrrEm1kdcrWJZI60Yv9TD4hgWsqnDQGl1
g7sdO0rAKBq2xBHZT8CN9rqVYX+WE9HCLRazpKs5u5ehI+TSzYdje42hqIjliXpu
VbOHkMuqi/DsRHhBxp8oshpqI3O+yigyZkdAoGYCJL6ar6QbEHXbncON5rpHDnBu
3S7JuUZ9+ECpefWAtGKuTdcOH7w1l0Vg7adX7opBRdwwUraq34XIqibNUslAmnDL
btXDCsHwIqZ1bqnLLWBkRs8zlbpQHIt/PiNMnhwbR9vRw/7hwK62YPc2qX+VBxBg
meYQF25omTnTZA3c90/k/RVpVzYkYe6RBadUch/Nr+AqD8KrEcY3KlPuD9YontsV
DA+FD4PlW/glfE+IaOhFz1xy28zods5hE0G5WlXa3mgzDp1FxVU+KXnojFq+vT7p
eLN1x1O/2FPeMUKbZm1+6XwXyjPrwhyMMfXl7nt/7F46rIrYHrSWIh0DRvZmzwYn
rspISVhB8q/pe4qQZyixCsSaD8e2mR2f1Weh83qsvOkTddHYZxFce7/8slmWHFnj
p8sdjgrxdSGK3MZl4Lwn9FoZPV64Jc72SxiRMj0kvCHATN3MjFiOt7JW1tGuoomH
xYEV1e3scvpTz1+T47kNwC5r1w+vDszlWnwZylkTusHuYsm4LkahEicuSIOFPWFG
bNT7KVpQNsmOKhf7YJZ9q0wBTsGxcQklWLB92jQHh9QnS34xVL3Y2RlgRWrev+Hh
x4nPnCpqIuBqhw9Yqob4vDDiaxF+hrO991kI3ldVfhfzxuhah3ZQbH5aOq+mIqRi
VqaTGtDBmTdhhx5g27c8abwSru4B+0pkXkDauD/RA1Cae+EdZmUuAcqR2OGVkw0i
ew3BxQ2RBgsqrMTZf96SvCqAOGZBA3TWtjCd9zB30ID2eTmV11o2c2zfFUzaxdgS
3ImG5/10bglDzSiG9L1OE7KiehmdvneCM6LeBBC/SqJdsmkhRX38jvAAcU0pxqYC
N8oSuJ2gno6Qnw/QchR6e+BAFUPLiEGdIU6drbfZhPGbu4UHp4DKMgRMc8TQyMC2
0GeF7OWZpDDy4DH6imwOldZx4e1fhmTjqtAzbYEdOz6e/Rjf1Ig35krZQYgEYJyX
2me1LK5miCPuQn4W+KVm0LEW3BJl8X7rTo7hMgZW0hjvy47ywMe9fiZvzJGWklLt
U46ZqIPq/25b2/rbuvF1xy2MrW1isGqpg9ZWUiSvi/B6JN+qs8j7XAKLiX7PP/wj
GjZjWTiALyUT57OaaGVf7siQUUxz1eKI68xuTw5Ad8nbJtNWMjzHY+6VbSOoudl2
BeZZaOH5Ek/V37c26VHVJBe+99pg/O/AsE+b0M6+DGcSjIMzoY3rMuKCkiZQGvzx
jRHEo4Gm2c65fsaDVKZJhaW/op6SAc+XK6N8khl6Z8Z2cG8ABMeyhgx/+olFaWFU
yg344pPOWAMM4PdDMRnBNvr5YeW7U6cAz9sHoinKnRcPgL7hf/pw0h99X+pfq4f4
D/8ewcpRz/05f5bXVWzqMV0abNoG7cdbLEzBX7XLh6VNjOl4DjpdIvcyGAirg1LV
FVJ5+6XBXL7sdH0yIIuXS6wYZ1pZXnCDN2NuggQiNE9hpakARIiCG1jyIxWq5p0v
eYKuYzezasvexhNe9NApv9DOjGruJyIYo8MYq+ENw/mSQ5YIJDCwzNPXtYvuKyFx
HBWhS7jlYt9aCU+u9YqeQ/NNA7GVEMMWKQgSquD//LU3rFV6wPekZpntlYBQm3a5
G/i/EVVXvVyQyvF1EygTLqEhqYGp7IF52v+OcjtiygSPzBkumt5knFYVAEBNMNCm
KZIRGT+Oi0DWd9gUs4WTvG3Fvfawfpi04G1+3LKfM2vTXU/sewnlaX6S6S8zlsuD
BPwCdBoNltpUmdOutmZMraABzZpZ9jkMpuxpESOotQowMV6K9puR9su91qH1Y5ZD
M4l+4jID3UwEyOMEAJQW28yihrDXNFKSg6v1B7Z7KozaYS0f/uMejUenHrk5/thZ
drQha+6IxDA/YplR0SvOIA+tZqPgMn3CcY6qoa37TwtEEjJ/4Sn6KgyHWB7OH1Wc
AHq0iZSKnJn0tOMT6Ry0yizsyAh92NJSkDhUzl8d9VstSKpbRXUWXncSzalILrtg
A/pVZGNV/kAdiLLj1LO2B5DFe8IJrAJSjht+DjF4DB9joP0o0bUWrMY01Gkgd7zv
1jeWZjuLIlgIQb8Bacc3QWMJWtbg2Q+a80FUodSa3DpmEDHzLHmKwEKWelw9UYWU
WorEBD+PP621nUEuKDmE38y+lEGqLfdC+Pe5e35X77xHcfrwPTHhQas16Hf72yIS
AuH8h8u9XuGX5m8QB7pgzg5JlwxWWWyj/lXbJMyB0iCkX6vG7/BKR0F0Uge/e+LT
jp3H/IDGAqUG9sy51ujYTy+Ihi5HzyzIdiaae2RakULZV25GdG0buQVpGSJsFLsr
Cq7K9STWejJ4ep1oMfNv5ukSZd+OXwiKq9Gs0ybQYrIVYl/Hlk0sI5qYt4sduSwK
7WBbKkWtUw2/voa+J1q0TDyg/VaP9xXMbB0nnk+k6Dy/VTxIbretfvNIppfkTFVI
r58pQ61FtMsLpfRhq1JTcKhGH0pmIkFuBmGZ7ypWgZ296Ig005rHkK7du304wJ4D
9od5NIJvrjXw8L4r634OMuj3qSzjvIpl23PA8aqsMNjQoGEvwDJo6CdfKL3A0nO8
Q2MgH2T4paGzxeoDorZHC9R+b27BuPTKRCUQwkyo1XbRNG6lKEAd1CYZmP5hGp3s
UuUFOJvi/4ZDqMsGXEqeKZlK2q3Pn6qz+zJFwnlaJKEf1OdivkyN02t+1MIUctBs
Due+DPFEOLUCvdhUg7EMD6ACRKsKFy6IOxoo1t2+P8e+sirLMFyc0DKFXczQMyDY
H4k5EDWUkMx2KnDSsyYretMc/vsXgCGZDCQnKuXVFuGSlmd7bFOLsufKTmsQ7iz6
EasIKSI5RBEeIOjeyFycZOkAEzdQwF/9w4yq6gVDK5bUKunXlgB6DnNJLEx7uFrO
BxHxmRAOjQQs4tklMi/knYl7lZVUMgyznjWaGwbF1TuHn0zQCyRdxJEswRoJExBl
1nnGcdFyKaRM+u093f3nCucGRxP668zh24vK0a/ftKw2TXJ9N7a+kZoI4XL42cO6
sN4pTAIjrc1QqrA1kB+LkUOywB2dal5p4QoAM73c4wVdBNC3ps5DbWxVp0qfWMkD
IVaxq2Y1i1e3LFjaSNLMNfcToiSLirMF0qVDnYIsnOs+DzGbgZsjSlFTG1edbsex
tinxhD+nnhujElqyuDG/9fZ3xH3OT/tS4oSpdMnck3ljU6dYvzu4lGOzptP3fk5q
++vKq6TYNdRgLvsJwuLWNjQEJn8ZbEPa9RNnwVaxEbmCi5hBRgTpXIzb9+Rx2cZZ
HT5OZ1hVe6CTf5iqGeUdKpba7Ha3+hWvoLcZiLcjoJyUBJY++I6GHu3ssX2Ln4up
pxslFaX8ADFwJcu8N7Cb83MgwMw72buLf82VQaUKFiBzMQwkfi4yErxUBzSQtt5/
XZ+ikfz0rlTcLiFqIU4St4Qch0dHPHSpZD1pTVsfI7UFUPNpQRfCdWslFMI+R8Ov
7W0XSz+/5I9GdHEJ5xU6YtS/qkbfLA8iQemuT3BlAqCy8aIQ/X1j2hBEftqB7udn
O5F2AglynkIpGvQqYqENAvnEHkekzKGS4Q4MCwbG9LcHzbWY6RYLwYoJJwC6+oXx
41xVZrmlBCtRGYfF2oFUukjyJHIF8bJ/5DtcstFvFswZloD3B9UpNYoiqc2De/ba
kYbVeZX+RZtOcs+2t2VnSxuLACaKyYCD9Zy5Y4YbD2hqGDK45SkLScPMvE1QSUh9
W6nIjqv7QhMkDDr9xak+PmscvSYIQplGnoaPanmLNw8VI28zihWeiEV0bSCrPVMr
8muadb1NmE3b4ID4k8nSY/AQo33uNIemn+UNDlUSDqYbx+17KLugUPf3tFBeczip
t1ZH/cAGHOJ85EWqTst3pVgyIiw5wPI1jI9wkpQ03TU8UjUWyl8quUfBeIdp5m+D
Q1uLj+nUsFFlteKffGX31yaVVPAY54C+DAMRpQKXfJjiQouKML4pEzpqg8zI8gXk
KU0tUhD9E5c7XizX6rMOG+mOv24d2rp2Xs/v5xDvHOvX6sRC/kMeQ8FYlGKKb+b8
cVOztrUcxlQxV2APgdIX1RaiNy5E5YEJjIvCN1zR8g59YnNIYOLHhUdeVB1cmhZa
ildSHEnqkBxhmT1ixevbdxIRSnt5aWbxXMuzVCL4OUrj/a9JTP0CVqQjsdy4NJT2
oDPhYlUFtv6A4iHHMZUU5qnGcDS0iA9TqGaqHp7hvww5vi6wuI5EM65P+Sdp3FhN
ab9baclCEYVwYTYuzHhhTgo2uuYCdrN0OHvh6L6h7ui4Rf1wAfAebkc8LZiT37IM
GszljXIVEqKQI4qbhIYxkpKFMm/Wb/rc/YRXsdXpn35VjG1dz2WOod/TStecTpPW
gEvoxDo53Kuk2aHk91CUNXRI3D5V7NlKMvIUFM9ldAm1FnzuD4RMzL65QcY2/a4n
oenHzq5m520naKmKrtmoz8FPxguKANNg56lY6L3feuVOaQ1LOyAJeoxNAytxQs3p
pucyKugCPDfRDhMkNpmEhR9m+iPTWDRrYHAXJCGmY4tym/sVAiDFGJc11Mrf1+Lo
KAs0XX988DDwE9uH0N5mteup2ujvIE/j4QNQgRPuNv1DwH8PP2KNDDxPU8Xz3PFm
+Tz3/G/oQZvUXorIXvM3S0VuK3HB42F9u2ObGaoJ8kD6/+6SDp3fVESs4PI2uAP1
fNr0hjED4zvH9bA3DV7ek1YlffEfbeYdRbE5vbqtyQpyzJi3TGlgkcNtOaM26zIz
pGAZaNfKSn9Lgvy8wMxCRD3djTf0uNFNrjMFnkgsff3CBNiemG0SJ1dzg+DhNaPt
t39ygZqTeq1gAjAIUzPjWWZP3y6uLc1GMWFdfOURmUqPyEoHsEXSmvIkUMk35yHo
T5wHbv68uTSNtcjQNoWn/2uSHMlwvjQb5nznv1ycU3VMx215vmJDs/gxZacH9Zcu
ELTsDiq+w1FhS+TaPGrEZWCzkVobnkQ+g417iGfOVHc4glsdhbRZ+fbjAoWpP2w2
lCBV98UKvh3h8RB75ON0WkFS5jCJinQJDCBcQkb158HxBaShjaFApP8DfL2eMuab
z/7ZKGD/HK6ivq0WSPmu4vUDQgZm31/U1AR3cBNnpVuI7UXmTHsqayD1doER4CHH
Jog5V1PHzS9/DTWq9JeUyLP9hktPYxaplv6vcgkO5eoHSR7wSgDzoaY0/sLhkJLV
cE3LrIJ7tFv/JKTbTx3oEt++O+ExhXg8/Edau0GcQfXFVRJsjOdAdmPKFKlJYRu4
qxWHGOKofi/sQEHz+udzOOq8paLKRP2poWvUK1DIWabzpz+YWmvmK3qlPr7M4HbB
edridMxS2Cts0ZyZxgmKM5AXZYErwmj2Hrr6ITBLsyBo1iXvgG4z/oqtbc6+kAFv
VAcvPt4mIXSGKC/EDqQXFsar6gS0ycrMQ6yE7tV6uq6EufWEmBfkQZO77UOVzfQ9
zNHn1Mr1wj07p/gH+buqMbg33ot38Dg7c3f63JBgmplY2uPutDYpPf5LcYLzdYw2
yWn9OULI6iCGyZG3QERNjMrQn1p0C2Z/MQ85iq51B+y9HNlq69a0zavlAhpqzn+H
Wdufqsrhhwbc0pyT9+BYHvDGgZdpfr6MWCTolVu9e1RyA1bOnrq1ZoPxNFgCFYMU
OgfJyLQNur/IKD235UhQb9pOgkcoM91g2HqUvWCpf/isXHH7knU8AcTcH+fBjlJm
/BInEtHjGOP/bVbwYnegCaGUo3ffOaUZIE4dkGFRM1lyfYLy27ufKfWxtiW6pg2u
qov7tPqRgMpxXvm1pcntEnrfgo5WZCN0WKzYSSawG+99zvc7UbEUhmKYHkmcKUsl
XL1725KdhZlMKOAn/5OiVAswR+E/EaeoZDOqtoGK3/+oq4ycE3QRuZyn+Y/p8/9S
Ldeyq0Mu6GAGEKiVGVIZx4+BASWlhAGIk9/tFuK+wX5xnZ2PCdvklgEMXrx8qt2Q
0z8C7h9rNNr2pHR44fhfDLnhVermmvaDgICbUY8yraHKZLOSwMviLkOUXoMHkKIz
5yLWlmyemtpib3bgLtfh2+96SKmCmTnEgbTopeFLXuMama5asb1Q8Kyi6j3L7U6R
Hk5aHj71AD+CfmaBD9kZQNHDF4ZvMDRgqwQGPtHF2NO60lUIcHGzQc6peKhfyTco
3IPoCozWz0o2/bfhegRB9TI2iK/zjM2Ng5iOUBsD16NGtpuEvHbHvcSbXlLh4TsM
MNfxb8n5SFzEjqs15MTFDaWgQAT9XNt7NlzXzLTJgQXbXcaxB/nlXsb2B0CmxRlS
4dtvnAJBnV5/esaXvYp2fais20lnBeed1H5tvEVlz84yWgeZL/dYrPb6YFTNX170
j8sUZDk8aht662sfRSdwVkOACQBXZdU/23O9QfLAyDMo653eMeOmxvl1sP3owrPr
g+zr2IWgJRrKiXP/x79Z6ODJFYL5g+/meQatZJ5SX184n6/W4gkcjJPv4ZPuAUZ/
PCrIjhW7Wwg9hBtylwzvXXwvIFovBO/2fIlDICKJUAuNRxsHyyOrS49hnrhpMEng
Nm+zn42yBII8NfCHN9yJvZTxR7EjuhD5Yaw4VknL00y62+lYaTeIINdULUtkS7cK
bs/HzJDddxOvZtmXsYBHJtLxuoyvAwi3z6WeEO9ZMUbHJwT0dSkO71xlaAVZx5AT
D9y00peJrvoo1pLi6DyTV+J3fRfAHejsddFo+5mZ2deCHe01qLAdRi51gFNwnSwP
UkMboeWeW7EX6qvScJBmv8VVKJR75EzOAtlsVbdECKH+DxH1kenlGsRVqIK71xxy
8yRzXIdvOfFWNhPsjChoty+YuvuXqcyDOkMBxY2kqDa2aA6i4fYvusQLibAfthkk
F9uDMPN7j83oC0GmMuwcR/lI1yr6tm2hbJpc2ik72qN1RtLVtsengiAMqSI5OGBj
uEzXzAzBe4hzE5/VmenlGkdN83XDyMf/GtIr40fkKQBGOYXC9gD+Xmo0d2qOmNkQ
0HXYOBzMtF+tOwlzUQPWoFcLFdp0I+fYtpO+JV9GiB67bPHRoOCjY+SB1OK/YE7d
0RmLTo6q5YbMauHcllGRAwOPoJw93ItsnwLA8NyhMj/zwMpBojEBfibAcqIhvB7M
r2/qS1kyaKvPOsnP8hiqIcmCZ7UAT6F/tBvtxjBrGayJP5Rj/Vd1IqlZ+f+6ik2o
I9Jj7T+QpXb51cKO9TJ7vobUOS7Ww1xyvwVavz6c7WdiCOruV4jJjkGaNcVOixNo
yAeplN7eUg2wd3VTTaRPRHING5BIThb2BIvt+JmfwelZV8zC1fp/nEHDbyUESOYJ
aaeecrgFiB79Eahc9pGwTPX7I/S6rzuhr4pLa7q10FLhKFNzlWUujYNGhsAz6afh
rcO2mQMC/bQlpYBk6fZdEX7cNHlvReODLhazY3APlnmfdfnjAhI0jXK03Z3eyN8O
kP33GdNn9YxYlqNZiVWFEXO5tl749xoAWthCKYgjFORrrcdIYTEDoWBVjEhquutl
8EpTRAXQ/DSom8dd/QKx/uaVPxk9PQ+pkskYNGczQxu1agxjboGniOU1BjX8lmYO
Gy/Ux/z6HXSgvf4jekA4u/PTso3je8bsO4RwuzGj17fPJPHfNmLJ2HP+akxey/KG
aFNNsaOUStA4zSp6ZpNCx5Clnd8Pvm0erhUyps28mn+QOGqZ2CPx6Jpp4i27+etH
fnmB2teu5XaeYPDe5qHJKB8j9gGofcXs5VmA1BCQUQba8gjitDzGFyFovkEe7uem
2I1OPx4/ri8Iej22eoW3fIdSRuwXcL0g2Z5F5Sazv0aDkqi1NfBCfHa9eD5qbBqJ
3M/QXyGKgjt10EY0kc2nR/mkp66wrChm07divkDKVmwg59IXkmZXwKfpydTlO8C+
65cVl6cdk3dPbRJQldEIYdBXhYdgZ6JFzStfu+Lo95cl5E1W+WuJi2Jw0RSr82v2
pCDbKSMnEX7K5sLCJL9KOW8BuFI79cWWa1c6puEvZfQ3BMBPkWMrW5eiIXH+BGK3
+A6n/7PL6jqUI4Q1iZSZXsTPQf0ycvvtm3OAMr7QQac/gbPrsbUK996UIbzSFzkw
0KlQljB8GLPc42XmTBKUq+3MExNV++HbMVOkzlDyROUje/0IRq/gJl/UFEvpB5oU
IjpWA+H+5GY/XdM4WXCZNNW0GE3+LOoYClf8/ToWIMEEpl2MueNF4wSQlukNL2e3
FvHrv6PadLHfhpEcKb7NVP4mMBBEad8Zpl2glvyZP21XR3WJ7S4R2JIzFAET4NHY
xR0SJkqnhjdoo7/0hbpfBO8QXQ1A/6ep7QNadeOlRDZNNg/tccx2YBm6rtD+mGsd
666G4Nxy6TPnMqkVi0DaprDFeH0E2qpd9oD3oXdySibj9mO0518xJgMn6PPzlDox
peR/v1AZwXsSMj5uVzTRnhboOag88sVJoHAxL7JErr1vsiPuxFUFb9FlYXuxPjDh
ha9jijKIlm4I4f05t6IbwgHYUDqDKCmIXbtdV5cboDRnDKjNECjeTcQPQ4L4vgPU
30ida/ZkpctiYFEky6YVKi3DBYVQ/Rpds6MEE/GpDkiL102Wx53DCG+5VYlkfnRG
s/mPDxiNIz0KFyWRfJRgqxPb5Sgtt/n6t5jszpPaCKhQkP+zyS6hzYs8KMPFJw9s
ZFtzWEobgsRNJZd4rwe5v+JZ3C7fwjJQ0Ufh6OE/dZAdeNpLs25PpG+366LCgCCw
UW94BvM7W8Ss4diQAbHowwihV78aPVSHKg/5HZjg917+KdKQhx2xNYsDEwXlygda
7R4pIhrMV3zEw8AyeRCgbgiMZ4mmJ8TCfhaGmy0S09SmMb6nlBJRi7B7vx/GBC/7
wcMbyPCIbR+lx9S6VUPmxMBnkt0lTngaI0O4dcMc/1buVzB70y+G+9Ss5HplHPBi
pK7w8yLlkbaWduhJ4CO/8MX5SefAbqUlWVUuL5MMEniX3K/9QkDj0ecE4k6lUbfa
t59F/EFVbwJE6tFCmfA7SBvFBtco7AaKXkJBUl9Xo4aDC1DfhRJOjh9iBeaIJ38f
AyJzvGPKqtUds37I2DTzRMyySWlpPoBsSxZl2FIQxjeeWMbtZCIf/4cZXMkEHwg6
c79c7jDWyN7jR1DKEQ1kOYJf17Ujnb1WOmDpTUFMp148O02rVSD0eOf7k/G7fQei
JvIgPp8MwNhx3H6DQ3njaRoGJx4GiHKVvEmOR6OH2WTJItprh8lzHsNejA52/uNJ
xMa0l3vgBsm27ZJcL50ma4onK43P9j0DejYIBssHb7UM0zeTXzR1AzyIL2pqsHt0
EnRZqtH9yiEW0pfS9rkNyrjeoohrceFaRbM25cr2Z/RDBAJilzHA6GW+ZIwdGJbb
6bg6oNF0jL6NnJ3GdJu8fJdqeZewRF3FSEmP+Ik8iRmLHK4ZRYKl0thPM7Mqwn1g
VAtoxKUhAQpWe2x32Fj2Lr+JdEtCyvAkcv2PcVpmw6JTSvsbDuPz9kzVCZkqYTfS
+cLWJCFYYuJkNqGeAmNKA1zQGm4NFrI6DxSEmXyekYTZ5QIZ46WxQvH9f0JZpDPl
ydSq1qLD0DMU11X+K+8tIjC5c5QgmT0dqrj+WafbJISjnJmBavW7aziG1iYUSbAb
DlYR8mDIQQW+2APYBBdqvf9AemZjDlj8ibL5cxbM+duszzw01ze9pDOQ2GTmK2PO
jK/ZpaeJwUDtCBT90hkDQCu9uV/f4+H5LxWQJjXkfMY0z5BBOHXrW55fjV5gvy7v
tOLsG/F23uPvTKCQSj8jwOSRIU7C0sEtPX0odZqwXJXEQ0XquqfdLk/B4QX5Iaqa
c3jQ3u0Zjszj2Ap4p+Kctkykn+Dvlk04oZXoYj3ohwlp2kgw+XZkZfUjRY8YNZen
tCizcwn7qqevoqJzYPkvcZwA91P5PveLIi2mb7CtryEIewohFbdIav2Xvjd3GjTc
quFbiMsiVt+lBk96WHMJA3CRYPdjsGAqqMPz4T0DHFnfLhCvBAg2aE2jaoXWgqjY
U3GGJl46D/z/M4/kYVD05Z469HSj5f46o3/Gh9N0KB4YJzUlkSGOkbN+OrGhBKtx
DHsK86wV5jYNdVsGxuhUJzgBEmLFFlYDGYDY2J4BI8sj56JNzIp6KuhpriIa/Iyi
j3EZxr6/kiWCc3m+VNaPgZnUxFJITDafTX88mx8DyORPOOR9KFSKwbeF7bV1+5UE
XFDy3BPUSVTR922gGsDBmgJnYC6PMAbOtAvouwMYDJp3uYEW7FT5PUjD1eVosnhA
a6YXGndDMxtUzjs1R29JkUtlgT57MLKO+Oe5nsNM5zX6JIINtV5HnhtwvoajkjMN
7T4AEEfpXBncbjCDsRxIdAp8rWcNofEJGEZxuAvP4rt9TT0uRRZf2mZ0mQ94MBBs
XR+E6JFbJjL6RqB8EacQs2iiO2snQCtKuhlf8ZxRycQcOSeINz1J4D1gDQB2pSnh
4107fTtGotOwhY8Dm9JwWXr2Yn/oA3VKIFYCbGX/KZbSCIkyCkq/L07uV3l1vXwG
XlJAIudJN0tNJGBlfmjZj37d+qp6DzJkBnfPIqxaRokxpg9oNhJ86ykm0+o5JgvJ
G7+incsaj37WdWmf33EvsfP7exBf3oH2SCFCQ+BOe00o5vOp/BDCcgHbbiZBLbFl
yMv66pb9EPXjo0q3YguMR5SWf52eEcdwKXi421Vel5k4REObJ+WbD+o0Nd0ghC4p
s+ZpZKpvHVmizrWIuIf/ouPB64DVEy8QBXCE8ozwWgXxwClyxhlvKoUTOyjLTOdh
yU/hIvuUW/d9Z/EBFgKrVUXA6Jbfxu2l4Yq/vo2I/pXFDZCvCTWK1tnZ7+3LY8dl
NHtHxaO5yfKpo+fie3v0vHGkV+Vy+spnFY+wtZc07Cmgz28pRZBMG0z4WAg9Dz4p
K0/+N7TNnmlDUyOnlNtf1TEYaAFZVOVjs0dQzrUZnSwq5Lg70bWiaVTe7pEDEB8T
N3wb1Mo+Vo1BrPnkfXTEWPrriVHjxx15RSx+OjL+Qzk3+2cmhi400qZ97aeihNH2
XsYKJtPDDajgDz57Xc6f3JcQnmdk8/WtC33+hFDM6sWk1omnEPqpBRyW5Ofl+oA3
JD9wIqbr3rFW6WvNOHwkjwhCuNetTwfhR+tYYQ2hP4cQyMzA+Dfnf6jIT2Q1s8EP
ax5+rpC7zXIVGQCG1lQhQ4nbAZH9UW6NRGXRTnaOhi/YiNPFFNd4MLSU7Vr39Stt
zI1TgihTPAuw4O4V6RRDlc32qvaNoMZP4fcW2acEJ/9w5gxzazUaDjm+NXO7ORnl
LeI8+XivOn1AuOUUguKoWzzpdOn9PTOn/O9hFoGyC4kt4dgU0Y6q8VZt7lAhoKft
OLik/WCMAlithuTJ2jFSOPnkg/rXt9nRXZLJwVVHbTDN1M/GSBwAWIzpvtRPiPXV
yCaM4j2MpN4hidUi32Us5BDTzXhbiqoTGjvtEmTS5/fBVq/ed7WstXEesGaFz+mb
BDedVCjcAMoL0+QuNwAv1Wi+Vnzy95gKouSbuC7bY7jat+xZvoLG6aU3sFa8gvIA
IQqGqqFqm3OGfqphYvwuIcWrsDOhhDCl6DPSFK+pSS0uBBedpinGkZtnsu0yQ+h5
Tm2bjvoPPW2Ph6/QdB/jamVskn+SjrcfwiTcXYpxwaDZL816fccNV0jZm9FxKyFm
S70XS+U3IJso4P46w3iWcu1ErPxiwi/QdHWH6g/uFOoCgD9mwUh2s/aC9x3+FxZE
gOh3eDcoWJONm0mDi3YLYouW9ULtGGaAwMsTd9SKmoJsvl2RnuEfYU0S27gGVVDI
F9RC6pFbPPXn2tWXkRTd8Bl5niP8lEtwP4kJFSWS97AxsbrhmmiRnoUp7pjxDMln
i0YpPePDGgVELPtrJavhE4Y1MOoUNd9Wf2KKkXabWOUQsZkrauOZEf29enITKixU
+4GpV4jriDKJLvD0v60Tka/vuoJ9lVY/YYPeR+8aZ4fNnHZDjLXGwBECqWXpcGbN
+l6U1ooxlGE5FNk9L35nSr9Nw4MODhIkJHc3Y5eJMdiSWo0apjvAl2VeZDZzW2pM
7ZZj7HJOIoIQ10YAX0mM/mydQhGjA+MfYU06bC+hYFxUBYZ/DPxzSE9jepKjmuvI
aoONpKngq1C3KfhfSONsBCgs/+RM+96EoBDNM5V+kHFuMPSye9E+C/8Cb0kw1qyT
SiYdQSBmmqEL+UJ68O+KcKVY98a9+fjCbNDSY0tPT5QtAwy8M4p9LNACd9OxlPL/
P03JT5OefiBtjnkudSsrLnvLwB85itM4Akdn09iWh5d9322mbY8awyl1EjGbjybI
aWnOWvxU2gv2UQanfEUMV/+sj1xWBbkIHYUY3l2X5QMMei8hjEsv0h8CmU27sPzA
i2QQ134HitbSjDTcJvBQJTTIapIP6WOOHb91dznnyoWjLS+SLq1LoyA9kCI0Gm0P
DA19VfdTUXDjq49gC/+WBoVSWOyntpJM7ObRecy/04QYi0+aULBFUJ0YizO1Lq1Z
Jw/BD3oBP/aTwIMP0JA6KuOYcPlm+8P5ucVb7iMJsaPe2AyXsoub2so93zjdr6Mt
g/70tCqx1vYlAkOYv08vIK1uqoKM1AwFxJ8irUwc0q6pBhjUrJsQkqZUIeWzDymz
Wd8cyA+4Fku02l0uq/PW2AIhMnmROeW1RH9ElnQdPm60V1Z8L98qKsfgaVOmVywg
MxZTn25Tm7+asRUy92QrrpeCNIGkosID0+rfuVto16jShYXx6046CeY0XlTt7PdA
nV84KlxotNGEOFp0WspHsfcJGefMZj3ciwyDgtkrvT/sRDnd8jDVZngINgEKNIIy
607y4EQ4WFeRhws2wKMZz7i4xxNuyIkUK3r+cfLc/aDOlw5FbG86Zlp4Gx31s8NP
NYAc7jY7vW2TI1I//VZTHy9Xy45qUZJuKa1rlLby78F4DpGsL1cIj9lrgBP0N7nA
scvDHyyzFA1Qv5yw+vWhV7dul8x/FVCE6eKqzeXaRmOGM/KShk72He++XfaE4EAr
mDUDgWcffA+14unJblljnJmLjeTAkhQFQ+yvFsGNWhPwZN3KCRnpEy0GR9x4FwI0
gea10XgusL2f+QVOT/xC4LOoMql0KMtEfwmXPsl/A5CS9Cg1ko4Lzb6vryULeBWR
Eg9pIynhQ8qzOEMVu4IJ8L1W0Zq2Tyj8B02ycrGutuMefECFhtOC8xAdtV4MmzLj
JyKPJ819gpuUpA6zM8/zYq6/XD5leD3oV/fZAAqj/bcDcfjqx1I6WYV5C6bS93m7
LY9pmcB5cpSvK+art46O6Cb3EPVeAaDDXfdq00mKGbb/GArkAO4LHmFbOmR1hYoE
lBB05kKBiOz9yy6C8MKLW7yiX2xkh4xm6sQshwopQ5PaEC2xNy27/hUWhMvDYbk7
656EribaXsEmVLab+mo06ggUhuARfYOZ3vjVxcUYzEONqAd67xvVRta7flVhyJIj
fwXJoF5n1UJi8irfw+ljbSO5tkTp44SIBwTqV1tD5gQTu12lvDbRoq5zIk4VfHWT
z4VQ34Nf2Fsu+IY88GGvoAD8RUR3+Fls/czl6mT8UwlI3YBIvpfgG7G8slkjWcLN
zCtNMfp/zFThkVwJD/DU87miD7gnFnntMqJTLRJG1MwOm8KkgA5qvPueMaU6l3XY
3azTMJTITsgYnQ80HF3gqMc1TAcyt8VzamGamDRo9d1KUCw6lDRS3O4UbzBU0k0G
SoynIdtscvIs/y/Qt2hZ9Cnyd8vVOpBPxOPqL2q43fa8MZZW4qT04mwBG3Yv2Wx2
6nQGmj/UZwfi0t833tCTY667Y5aI8CJq59TYw9yMzTYMaKIU2Z/supo348yOgurp
L++WsK7XPvrvdS3YAkgzR4IanMXHa/kXYC6yyj+iZbvabmlUvWlBzM4QaEtZk+aB
NwuoAi5t/4W2VfIRKpvZ/YzH6pfJULeUncrRxNRjwWNQxjdpZqp2b5xL+YJEre2v
uWF9F37DoVkoS/uN78qCr7tB9fAXWUTHk0odEt9IMX6AE7RhSR1vwpFN5F4EyZIw
q2kkgFAIA9yb/n6i1R6rcKoFOcvmpFAct7cU+VmFzSKVyYFBg72zr/wRtNvedpBf
wDB2iEfLdJdak51blKzTzMKrOyiAQsYmCA8GUaMvd2PXLrHTw7KsYLNSBEf3ml2t
AFsrtUhhrSl0lwC82Jm6smUl8nlG8jiU9aws23/C6Lr7Ra3ryS53Np1TywEWDfxc
dCw7rNJvWO1cofEOeSq+LpfHi4kLvq4Moym/QDDZiGmP0uUXcU4rXsQkBD5680NO
SrWWxTh7BApE+Bxnb3KQrKfv0S7IEO64XRZulCpRENqHSWD+RXWImJtMB2e6Q8eF
oIXe8UiyGZeMbFpfyeISWgOhXYwf7NCknCHbvTaxCxB0JmrGz60XIi0sfjs5Dt2s
xxiw14SYSbRIHgCo3AtJ2xeFBqHAj1XVfUpJm3BWKvmQIdw1mQrv8i9MAz4aEZJ8
xD4hgYXfgPA/wFRSHlzG35MK18raqG6V2by6BkEuA7jhp5RmM4HoJxu3Uqcm0hmZ
Ljo27VXZFWMtF5bET0jfBdt7RJRGSEoG3zrNl4v1gTtwxNf6sZ0vl84B1smlkwye
SlwrcRUzEgQ8hnAvYiekIzl5hw0SoTG1myocGwLyZk4lf0de9bjg+SpstLyq+tcD
Tw9YdBoqPzYS3NpBaocHs5t9x+rVo7Oskxfo81ecnXjEtHOxpoTQju0t8xA/Ndg4
0PHKmNKfByvhq/3gRfP2598zt9MilCAB+E7lZNq0+T+co/sbDaQ/twsE/hkzF+qE
rqwpOER11BNPGL9SIWwus7jbb9vcRRAetgUaQ3tsOzVQCyWHDlIS/cltBkhwrPC0
OS7M8V3UMfK7b+ZyHK+U36h4kcLvNpWHs1aC23gvSQYOy8WEZCqUtVB1NiUiazZp
ilR3WkhGCu9Eeko2A4M2QLPQyKRGUIX1Yla0JU0Lcelz6CSy8/hjmjgZlnzwxyx7
vXVQRAi7iNVAQHRmxEfRfYx6n3uGKh/Ajxm2MeMrVCU3CdhuOgMs4IbglGCHFLsX
8Jb7O2JqUwRByl5aLFSo14hPkdHkZH5I4xAz97KrlaDjfCuH3rCm2SppIo3Od9Hs
GByJGS1Sy3OiKMVCHEu75BGqBatrHbjMwS9vn16uYIx+6Ox9LGhZrUjJFAtjKO5a
mYPsxDMOpckfIYP6Epeydgb7yvr6BZ/DBmd3B8gNXOq3kim6tU6A9+2GIHU5j4HZ
KNIB5m4Prd1mqNouj+MZi+0AiHvePo7S7gvHuT22Y34H1Rk0j921PLxCljGz3x/c
00R0fUrpP4a7VwwzmM9lJsQtIdmADL5d3K+ZwFVyjGtRRr8P7Un5VWPGbDbjjb00
3YvLQNIDq58BjOGCW4oXbVbcaE4de5r7zyz9XHaaDNpfGAa9vcobRXOXlVmdY4Fv
xqSzSyAuRVy+YcxEtC+iHJ2TWF7vECKSP94fy+FHFYv2Df9bnKP1Quei0iokx0Mr
dIwGB461+T4jhmAlkU+nuhnjyrE7/AoXW4fgRXk2ovx6rQUsSkQoFQpO0n7/R4Kq
eDnkPmp0gqBP7yft+FtnMhIpCzNtOpGwl1rSKhZ7+pgXuiDbqVGvy1p3r1RDd77C
lTEBmlpd4kJO0DU/vhXvH+jvCkiqNppak29r/ng6KEx3t1ff7bwVPpNvllAZE98Z
AnAuXM/sFiaCJjvpvgWXfO7aNPm09Xie21uly3uHsvB2bxc/rafw7DGCgkruRGDi
bp9NeYwJEeLHHE+KGFEwL4kYh8FMz6UMzl7zKnD3DqS2XNICX4fgJajX4PC5RNOH
oI7xu97uYo026xV1Ms1f8b1dHEYGHyYjgLv39zzAb1TE36llUXd1mc2hXebNCReg
HvuUvgLbR10weNRoI9X/hHnMCKP65KiMdSMAO9V+wb8WJkMMs8sjgtQRJ47BY9P1
gAKCbpYNp+nhxNdo8MY8tBNOf/V4wUtgzXsbLHi6RpfTwIZGHsdr5moVC4Jg9Yn1
fP/M6vFHBcpB5YpOT/yotoZBTI5aqeYxJFL23wBOdGqnsrd3Y11+8/bGiS9/3UtW
GBoPY5pe4/LGGGKaaHZwNHRSrgJm8ZXMtGfF60r4KDFFkIgVoeyjD2kLwTAJ9ibf
4oBdbNRAhRFS3CJaci4Fg43y7Dli9kB2kl5xjHDVtq3cblihn1YHZNxuJlWttTrg
B00a3Tt/I7P7i/RLiL84oRDox1F80xcLG+UotpuiA6XXg9Gzyk1eKDlOk2m+b5fG
rfF0r8JgJ72OkPuGtlv/igu39vAofhCvaBOsBXZqJ81QvDFP9dA4VRqbFVFrQSii
d7ex3hwbY6eFPc3WjczCHfFVfBRkek27Uvxgd04YZNPYT7xdM7D50AN4GYBnIa0S
Hb7IF8OCKl4PZH8K+AA0WMqAIb+tk2q8noQiErqJr4SVfWA6Bu1uZZrYkZGVGWox
B8qyi8G7Ajt+ZaW0LLxpGKMwVSYyE7dYUQWXjIy5lGl3F3iHBueGQmaVz5hs1ZbL
ILe3VWNAXpy+oSkGIwmtirSLH8y71pdMjU0YDWqaS8dviuHFHpkdsHTowmZ6hBH/
jrXcIzHnUTMpoKYpGLhfkwcRxt8cqPVI3XqXmC1vD6+uizJ4lHZhVLt/c3hGIL8m
a6QwzovZSSGIAxLHo6VPM3Mbganvkn/TWsL4Nc2MewcvoitIUvVUcrGwXat1gFeC
iqi6NmuQMKAAtOeI+z7R9nxFEGzNPduKxFk0wJYd3r5FMVmPP2O0zuueS8F356ra
hEn5iVB8FYk9UHciUT8/8akmgJILMEItMCvBMP5YmLEme3bfNhCpnaJp6ixRMcgx
yzRouB6vw3/i+i0XvbRIu4Kg+5JbKcfJMjGzPGwy4zgI8F5H3d7ql+eAc0nOn6i+
k+EcXCE4wsYZ/dy4ysr7cH4JilS08UQ411flEKwiHJKo1wfwmSRMWC9yQJAc2NHr
w/RQueeOgU1xVbdpySfQrRQXPORUXVC7b+YBYjzb2Afl7Jd3WY4kUBruBqsoh5b0
Vd1AdpApZvUpB5gbApwE+vGil+2LaZ73sfmWYAGM2a+9V7pZYHUbQU9ulL8f6RMO
TicaeNcIxE+7wNHyo0dI8dMwht1SIGPWiOea5XC4qzzPFQI5kJJoT/KjfaqZoLCb
xcN/YECOiV37MzZY5+dqm0l7HESUr24qPSZ7YB63+ZDeSqIe590bfysDhrweWBHi
0pizGA0OfnDKXU+KT4AFF4ING54S0J5ojSdWYxMzpszMgOniP8msLs2NCvj5eGF3
JbATKIDkqt0IGew5rd6+k7bgHYco+vTZuLFo6G+ke4VCjTdxvoAzheEGwDcSAbQs
vDLVmmjDs5shH3jpwYg3fU8ShN9i+5BivcVE845Yi70UmSlF+oZxARwIYiaKrY4t
O9Cp76Ha5Jsu4OKrairzW1lwSwQsUA/96WmMo+4Ms2K6I/IDjr9niCNIqqGtWL/W
mGikKc9GwJcbugxpkmAwMH4G3qii3eqLJKC5G7/2KUEb28V8zr90XX6+bDeqNAcV
J21itETm1Og49Nl86JEmUc3Sqq6j6D4VRIfY17eK0aaS9hUUa2MzU0zF3+13SyJR
SibbFtZv4OQtKrY0hFqKIbQbr/xWlWMfIW16uR8yKtl90021m/VaR0VnK4FaHjPs
Ci7fmumeJH+FpeErZGkxHn0OGqKp0zynhafOweUZxyvATNTJ04ujoV3etOqxi6Zg
XK3H+ynD6LWYWjXlCQf6NQFe+tnRHRT8eHI4BeatoSewXYl56ju7dvs4L4QGl23X
U8dPQzb04uxzgPiOqnN0RPjzGUipe+2MZ3W4nAKV+e8Fi/2/hkTUAHP+jhKUacpr
W5FtRDHrhx8TewIeUBB/xz1QxgibDVXte4GCd0kxl6HDkAjSHx0dUirgrWhZtTNe
jLeMxza38YHCwDZPlnx2x7Ct8rFORg/uTR9tixX6MBtwFo+14THfeEXbv3BQPCls
C3m99IU1mAZrmxjTL0qu59tvR66j3XFw5dk8hd3wbgGpwK3wq9tC2PTriWahzEbt
zZV+ob8/m94HRkGofW7Q2DB4z5u/gGoZ0jiMNTov8R90SBqJ7wupKXpOsIRwOg+v
5l4wxO1ajawn5Oh0qYPK9t0mHqnRLPFbdRNQx0EzCOjfGwKZuRQVueYmNf61ZNzi
0W9KoUk0hGEQDBNaQrnMwfnE9hc/LGew+C64vAG/EKg4C7t5JMZJzTuU0Rq/574T
w0s0o9IUD5Cq38cH5ruX0+ja54hpldlsqhO3oGp2Yzy1kJfKAo8ClXkKfBKFIslE
FCYOz/Iw+9NCn+fXGbIeeEejZTAO+0FzNvh+ls8pThVZ7mzWtdLUye0fWn2Zr3Bf
2rItXhwmUBOk9kPc6yeElxS433KWqbJ7GguLaCzT97gPWZ63uyoh19m0HF+SRzio
af0jRTwMltuyHyK9mGmdL+Mv1aYbyxEf66iswiVj5tuE964Yd1bJLadFOI43VCPX
OabUff6Ry5OceZF28WmtlAmQqQXbt0Cd+C7TJ2VKjBQchWYktlqoGzTneuuL892b
QlYq6ryNC9mIn2gBPsMu309N5j/29R0zM4pvJuNah/zGzPS2v+koM/d1eb+kjBkH
VdoC4C2szWA8HWp9/FV9J6k8VjrxiTWTxsJsTyptLj5rzb4gZkBfJco+AEu1Bl5g
wIoGnh+fwTJGOGljkiGNdd4LesvbMaoeoTrm7/7ZjxOHo6tqjhjIa0c2Uxbpw9ig
sQugzxHAXkW4dT6RCbMEFlWlc4z5dWL3bzJBVhqaHLbbollJdXa/e6p+C9OvQzY1
VOARycvmE/sTHcl0Ox6Q1rHjyTVNv7GgSRqigV0EmVu/apvPnM1uHdbDDf3XYbOm
K0XYzVBnttUt7yB2WspglveuPVsvX9kPAb/ortNFG1I798cWR8+LMHqI+wcHfxiY
v8tEHalWaO1G1I9fO5hxA7NBXvm7DU8cmzU6Q8u8xjhBqCa2jo7UEOzpCs7a/TOo
rP3mPwVt/V9XDfJGrA0kzEp30nqdVSEeErVF8qlQKq/pKWe4Kl+WWVjKO9yNfj6Y
cMAhagbZzcw3OrTcIhe57Xs3JZ5AuSjTowzu9P9oD3ADbNwINCfNPjBd3LsJDQZz
2GAa0gi3EKWc/9Q5vDFpwNa6OstpjJlvAqkemY3dnv+HceOKSCPTrjApGBWldrWi
5CWusb7Cm6T/Bt/huN5yT2IwK+jNIOgKaTEJsvo4pFrJfTxxuIa6l5BiU8JsjdHA
NeLNAbrpc2mLhkWY78+yqAyA0RiCeFqw8r9qNm1A45XIW6sd54lVnih58N7E6VnZ
VCi0UR4eczl4LLTxlP8l8HYwB+4l5b3F6PlrqLDBPtqxTltp9JvabLo77OmLfGCD
whhWg5A+RKxWpw0yLPstttSKxu8i9q38IVWHZErdXuydX/YNRfNDttFHG8FVESFw
miqyEGYt7RfCA++ASx76AB9CH8f7fMT53KHaY01KR/EwJ8ydfp2Ejk5iuWENx+U9
NYiidERRmOp/2/r9O0k0GdOqesByjnM6h3/aeBKmhrESIcsD/N7ZmP1Ft1Qjc7OW
ioHK7EZyRzpg3y/BQsMEQvrD+6VOrX6HDtK4CkJLi+LTX+E/AxY0qG88xgg0zZ9c
XGjdwQmNVRLmyxsnEYE6CmPnT1OMd3WrLUnWzv/gS/PsnmCn2pC+SUFYrLkVaWe7
UfqQ0X/M57fl1atjmXyonNwMIRgJDupm+dZsEbWSvRMGTLcaEat6Qj8qlLKZxdXf
Fiv6aMXVrT+0UeBPU8K0jOW0rhQ6LluZrFkIEmf3tYzYEZPyy4LMwSnMeI3Xje/8
Ca2OKN9/aisQkr81lUIhbuPRt2PaotgYiJkZhB4NrV0qbVaw6OjgMcjvckqAe7F1
oOkBPi7WNTAQhjyWDSZjK4taAQnzStTYJhxzSWxWaqWPUOoWxxdnfoCvGVRXLvvK
sUgsbkJ+FLAvPGSYZQWu3e6Qa7RVjycHcu7uQsiMeI/tAgH0An5a4mB77tzKTYud
NVgaj2elKzDUlzzMdhCBZzGu8xeZ1PNtA61+htS5AQXDN2L2W8cPGCU+NR3BpKgz
k/b1tkC3Qig50wjvLrNaPj09lgbv6PrwodlKe0OazCBpcWYpW0TspTwWmidLgg1s
ynnu5qt/HwWEPUgZ0jXAhe/6+kJuYeESy3IZaHaiabgGuReRghUroLrUqZ76ie6U
njExIF/1QRzonZKw3kLtzWfSQbREBZud9bg+eiyRgr64aXjUKLz+6n9DZR2gS30r
FNsEQ9IXK1rmvUUDK6rL/upKZbK2XGjur0kuV+b/1JlfGLP1FN60TYqGdkk7eELi
uRjEM1JwsKjhydZPhf8MkrCjZZKFlX7Hh4Akw7AsDGfkKNaOnkDfgzmwAJgT7raF
HDonrC41l6b24XF1AtLVR1Tz+D6dXtH3mBunK4gCQ4av0oCgiR0YfGlVBk3CiQaw
MfeluC41lhJ5rJbTy5OjJd65BnqLcgPw21oe63Y2WyRF/ZiVYlBBkjDJlhfLTwjG
GvsjkfWTyFVPo9dIaoAvggM/48aQxl6fsx8O98S59al1Ov0kwGo+TriHRthjVk/L
+f4e2hBQu9LabywV1eC9kBtLXOqpNlB426TTf2Ax3PltzfCzv8cZHLPjFXrwmals
A9OBrFnVVlHEzV2MHIhDc7QEDRweJIpKUMLikvha1i8jKFm7ENUL9re0gJFPNcLm
9YqnQuCrLzrxa9fQI0lcKh8AbssoSlbeqqPmhuugv2kYwOAB0lZyxi83YrtkC9Rn
E1kC1ZVHhINGW1XAbnin4wZVPeJWoRTBF+oQwfBsx4kN7KU4IdnED3Mhd1VnGNOL
ZgLjd3GlhRSo3XJqAxT9n/H8U549BHERTdph40gIHy67uw78NGsf2GOcGFNACQIB
HHCOLpHkwV2tY9dlRbCiyrPaY7c2s+qBbMx2JBoyuA9GIsETryJQ/rmYjHx80jHe
WLwqH34M4RFhaqQuCXJ41RpFZ0Wc9p96LE947PaM1qqoCbFuMBcS/HBXYMTZgWMi
GI6br5OYI8FrVyDhBSe+dSi3KRx+9J7tiPQ+dqe8SEISL8ypS5vxhJQYoS81kHJQ
ylGcF/S2T9FgMCA39vHHCeVIpV6WRk2uhyoDlfz4zhF8zja/q4pn17q+GN8WrOtA
rexVDwxKxigla353KCedGIQAEiYZ5WSaa3a2z4NGAdPhQb8a2CUCaNHG+qKYOuno
uUJHB1R44F4rFovTEn3V/YUgBGdbLWmhbLeZxo5NciNONoLJig0Y1M8hrZSV2BLJ
gDF8leK0VI4IrF0aw9XWmg7TUvuwCYxTHTzlrpREIuuZX075LYjPMWaN/P5jRAWx
C3rLw6RQDhCcgq7UiURP3KzxTVyOnENwza8buhFwCOFzXhZY9Cn13t0id93wJPxC
LZ+2fRlpp/7yXPZk72r7Th/Dof3jdHWI62i1UvjY3KpKdwl+m1+3NywxAmYYt+oP
46N4Me5TRdXiXIRHeFVD128FaCxoZB5k+5TZ06vyi2jG2vv3PMqBRFvsLyPb2B4w
MCm/pOqNQu8jRRlqxOJkYN+pa3MhfL5rH+tGqdbjEf5WeUN8FxQAWU7E7t25oF53
94tFEpb8sWmLqizw27u+eag5Ml06NSW0AT8Zsr3FN4wWO/riuaojDAuXeaG0KpPx
sj8tR0o4O6teyEZO133K1hCsHLXqH7IwCyAzOAgJEUOBoqeSqBcTjdAmP6AG6fNm
C9VNlMJ6s7qyZ41fVq0f7YajGgVooJH01o4HMzrl1MrtfWutCDcsGvbfYinW0Y+1
bCMFyQGgNc8szBbAVppMUOtWQa5QKGHr9swSyQOweNrLelyqxJam/z4wyEBMmEiN
ZhdC/QX4GXttS9OFWsWh4dTuM+Yr0opt07l/go7PJMqE0IM4tY4jTGpH5uSbAbKv
zwL8Edpbn93Dt5OU3L7Dxy1BOxcTAAOTl5z2ZMj/5X/N2OwLYw8A/sBmIQu8Tr7g
5/7Um8XX9Xu/mopLK/O0gy4scWg2XqG8HcYZb5yTal6ey3IaYqMwjC+ICidpYcCF
7U3Sq7V3nqoD7BY2hdtqF+bogeN2TyCivnMLjkAxhcCo+tTtDAiqu+xfIkEh9+l7
85HY2FA/7OA8haCZsUBJMQVvqPZmJTzQ20qCwBHlwYAIlcPs/1bSfAErdEWH9H5t
8Z/f+eJbHso88mvwtyUq6W3eJIlAEkhIRD9dGIG89LPm0cOXHkGhq/oGINkgoYrD
rQrLl2ktZimTVJiAmhlryW9OtcyxX4h/9q3Du6nZyzh/iuc84gXSnP9WG7w198m6
Pyg9iMA16MSYRlunkdunaCcydrv0PTASBvrY8Qd/oMHpkfzMc5sSkP5ioaK0Br+0
GLrX/1hzd9ppbx93Ru4HnuVHz/YIEA1yj7phy+Qx/JcxW89UcNEmCpjKczDEu2Kb
U73ST4z8CbouXe0p8mkT3mcGf6crnCvNbiehV3jbMW6+EBcFYvi4ASBK/5krJ5Qi
3uo+020Vln96CdOkfWZvXdDs28ULyStv46vNOuKAqTKDdxZuTnsLI2gMVog9LOqD
zwxpP4KUN4rLTYspaPZwV7WroPIFzV6mfCI9JCW+yppofiBCW5xrYTdLvnzbh40c
+AwLixP2xQgDU7BTl1vP70pFDE6K0/MZe2dFqZ9P9mtuIgpe3Tp0RTbFBa8LdSOY
gLPOBfD7vwim38K8PC6D/sPSpAbtTzN7dSWZwv04Qq9c5I0ulPwwaJT40DyVHFkn
ongF61kYI89INFyNlb5lO50nDx/MnjSyTaq/N/CSl5pZCPRloTBk3fTCkNDVqrqI
NNWNqpzl9iMNo79BlSOR0u/Hy1wXSV7dCp2/HgVeJraTzc2S5oIKT0ECijV3/uFG
5GLAmc78pJu0oLNt58x0Ko0UTiVajMeBZk1T4wkLtczoCob5w6KyPqyC0fOOaf4l
kXp67bW9BybfCUBWFvGcW8tOt1H0s+yTcIfDSOal3EtYlgF1AkzIwqMgS2t+R6dx
Wk5gUfnyFDDKz1tvu3Dbo92hEAs4t2s/cCph4D8wIZK1XLszD+/p3toUTRC/jGEq
q/7L0KGxtDoRbzkKo680IY0UVLw5mx73j7FfyxABVLi/YCAKrL0w8kFZbrOoZgj7
W+nS07vZaNWve2SrO+i2VzcLVjdvN7zD9t5BK5c0O3nDkkxp94fV2GoT99cfTUXh
y51YIhjDhCaUnEqnhh3WRc9WsrtzwN0oJKuuJ/TEywEllgqvnUhoYBhPgu/sW5zS
QoZf3dJjmApin1c9qyTsGq/emCSksjYdG/o6Lgl22zDqXW87Ru67wJ9mam842GUZ
PE7FOGkRZPiH9D4ZKuL6EIAH+/tqOXFr1VfyfvBipiIr69KeRvfA2CkOBbCXjlxX
Clm5paxcS/mpH5nxfNlPfWD1MjU/pS2pqZ+PKaroxp993ANaUWykop+yU7kAs8MD
LFrOgR+9ZyKiqx5GrYhfxdQQ/VdS6VeqC4OAHTBWT/0A78+NAaXKyAypLr58sccL
Q+2L6eGk7XEXsNZFZirUuoc5NSeqwKNkHP2fHmyQFh9slg2/A0oWDlbMjMdslqAZ
V93aYUMOd7uNbjTQoBIcClWakgocTk77XEIgNqVwpwUEPgzv3IlS4CqFxPHQlsPw
hVTQ6Phn2FQw7ARrz2JKonuhZakX4jtuRB9L9L9Fu+I40K5rRl9UF55NREqrbKYT
hTUsesbPzT0gh1xBBFPbHrc0y83ahK41Kt8m5AWJF2Y2nH5Jp3nVuyAv5nNNRA1v
oS/zy8/krHF+NPLiRwfnT3G7aQQ5VaKhIxsSmi26UeBLcAuKVWV11J0wX0QUKDhU
QDwQ9qZwYl9uMcmvUjihKmpg8iD8ZDT0NDKB/AFR4f/08vsqVDJu5OK+SSbNv1Tc
2QE6W+i9qCAoajUxVO1eyg6jKSqftSaVIa3i8SElevLn0efEmAA3X1AYsG2NjPJd
Xcg/gs8KpPgapXt8t3gM3aX/Wsl87qS8yx2jwJmvTPglyjHbaSqBOVpZeiUYeaOi
D+exXiahMxhTvGrZgULl+e2fsNEFFrGJn64IJ+rQKrxEsk8IAbrvgT5c32VFqFXG
BxNeVo7IHBx/ekZTZO/1jy6nCGRWIEcji/wpsEdkwWaUjreORoExxK6dH17Kvo/f
x3a9c8VJKSBbede2cmOvnnYR7AK48yVXItei0VX+kHemk8XoVj0V2i0l5PdIvJwr
LAHpHKPCqr73fEi7x/VmCmkzSkU4Nxmxz9FISDyeJWeEd9v7Nf5NA6hLSMZSPQ4o
EI7IK9hOJVDxJ1oBagIyHqiz2WrEeKfCVkKlUDMb+OK33TEjL19S5RXr2MepiAqW
g2V4OSL97kBAqaxMOqg73QpfeSCgOy5pEN6kuOtubzCmcygQdsw6+1v4f8FRo7aJ
TAGduE+vt73L3w7AoiT+fEZ0B/5KxsCl7HBn0/cbDzK3R8b+xp3C5oNJliHGfN8b
M/XnVrtLhonyS7MUw7IAGg1fZS5T1lz72hIbH48HavZ1s0CVBxQ59dSWJFUG0R9Y
fLmAQB6F90gg5xG8QUFqoQHrE8exXbb8uQkG6bHwcgJmTSpnPoc2PWPxeJIm9CE3
hM+LPH8R50UzEOc8FuFqblOVn3fE3T43kuu7A1CPLcP6QIzWBnd+TRm32XY7wuvp
9w41M87MwD+zoKWMiRdgWoCrz4olQ1udechSs8bD2Y9NT6XGdcIQzxFxmoBMwcSq
xrD4aTfqd9HrXU89hFPUgel4D5uh/7HdbHXgzVcagYojPtiLQAApq5VaX8jS4AX3
z/muRRzDX5zKbqgF3yYut+7vNtdEasV8UeY0aox2+TUJ+IYdl+RKCzW+QqnbyKdF
FQqO1oOsKj0uVQlm2WnH1bQc5TvX8kpDcZWk7FFlynZqGCqUBLlPxNXKYmLKHuaO
BDBLf+JysRe6jHjITiSIOLY0wtvwp7GrTBDRtwsUoAiYcv9VoYayvnH3oMzW2o47
R8BT+g+HoNnqwYigKLM9yIgjl1IPxUGAdmWVos5wZJJpWqhHgTqb3TKGlKbmMNyY
3Aya7NO79LSgqsuAtmEjXplDVoLfnXoO8kHRQTmPrhqklfU56SXbA05JktjsnxtS
O+mxtnWgW8qNkkn+O0oJ0XQUDjuy8y7tUlXsfoEWUtq0uy0d0Ztgr1XTCepx/TGb
8DubqTbHQMe3q0xPM80PHpnzz3nCErVzXh3ds2yz0Or6blcYFW6WseAUbqf0pnyt
5vrjfDNXwmohegngBIDejXn2qSmBotcqkP/uu9PFhhrMFDd5tL8DcHbpgnwUjbun
DI442RXBH7+P2rzdZDMazflVd/wOQc5+PV/LplkDqimzxTzhTLyVPNOJKgfU78Gx
Hl5kBWUrqaxtSxsX7MskKiG8irdvUOJradsyR0wvWoGbztDQMugFCpgi+SJFQOpP
bsw1hPquGH8/+t3KRi0IN5v4we8E5T7xnsMLoRAXSReYh6+1hBdmpxt7fQaG4Pp8
PXbHX7FuyPtoiRtcN/I5tVCWWT6TEsbsWbjcd/dIA4WeuOWGR3ra3+l1596PEILj
jqxTPB94UfSCWQeVOIwZG1Hg4eL2pGE7FbixmS2mWEMDIL9rhwwfrsgP8trzRkRk
z4iuPq5wo2B77Jve0P/OyqXqO7BTRQC8j1FvzTCOvbrqv9ZOnZR0JIi/LCfbJmie
kFJtsP2Y8c7NBlBnkJbFIAxfr62xDU21eDCLVCW6Z4zvCw9YEIYSYa2y+lSgT40A
/hmtliDIjN1H1vnsWEuwFbTmzDsEkmaqoUz2SkH9ofdDFEokgr6ovO81Y2IfpBYa
4b0YcHIKK+8bAPhj04/4a3KMoC5UgMWs6P5CGv2YmnBLa5xV+Q16tOFbluw7glf0
83Vk968lRvB45PZhOXEidrUvUhVJTyoLG9Ls4j+alT4qjKgMPowUYpYygtYDw6PJ
B824wd1gPYWzI4AHbu558Bv+oS0nFrGHEk7Ud3gV1fyvMgUJf042c9DZ4rT3/oz7
entnM38++6r/0fB6qXcU2Ud/hyZCLvxYNk1rytw5hLToA8gPMZKhq5XlACZSCHgq
awlVBe1GPhkQIChUNlzUSz62p84lhgv9G/ta8pdwo6eS2HFnSAldtuEFo7ZHTwNH
CDIS6TzmU26AdiiIJeRovDzSoUEU8sTyXUpRWpH49SsC/06Z+5zxEN9ifXpdA43J
AqiHgOfcS8WCgwaAh7AD0eEZc8dmt+t0XXwEvH44h+eBoyzVxBQmeg42D+Dke655
9MfC59llti9vJSZQH5dEBu0XnfBKKLO6Teh2RzAF7fqZIj8AEpZOXFbS/CwL9SJZ
Ix17/As1pIlgFVkzg8XnB/U0NyY1nZSafUFjFPlTjCF1Sw8cSaTgKaY9nn/5YKPi
T5Hmfnh6Z+LC4yoHMTBrsCrA0Bip3dwfpuEwLLvAXNLcoZmt0iEoEyDMsoHp9/tN
PEKKKCoIULvfI4qdTkwGJJtuSIVsRpYj2JDnXRW0V2gibKPdalTS0sfj5yaP/D7Z
udgQyT3Tyfaoc+Pfyn10zqg6qRnVsG9/4QH/iEbCdI0vFmBg+sjUkM+nA1gOpIEA
x5kFYurAkgFCVMEmPEfXX8O6v18Nm+gHOjYU9pTo1MX6pdKhH/34wPf+iigNcpRu
TgWY7W34PSfQaxQBNsFQghK9q7andYjE1I2T4UYrko8zpMEktr+Ggg45e7SSzRI7
xaYTyg91btBhoeuzOV8qmTKNHAWndziZXZdLY8iPTOIEZ0/KMihmw59aeNmWoFOl
4bvJrGYyXdlmhCrMCLG7Jwp5yigTpIsOEXsuLrp+Ju6Ln8DA5YQXnvgH+piufBsV
YP1WnUtFMgth6Vlk3bvMUr7/VCV5AdsL/GEvOMzmGx1hRiD0metWdXzW/pYMSHfb
gh9wO1gdZ3m99DspjPXLOKpGZPskY4Izoz/X/CWC9e1ok4L9wgN9nlB4yY+w3ZEq
BLZmY8rXSzkBfOzR3vDfvv3NTRpZdCew3Fio8RztRly6kanufskxkVPNEkxIM+P3
9okhCw5XoBSQNm61zHSx65syvPhum679F4Bryy/+kG+LzbqZnogtVJsmrtaPpCd0
2fWawpZJDY9+Gfrbouq2opKZzta/6HSSAWXn/fTohbMVcUERNuj7/QfB225SWT+C
NMq/yBdZ/WjJCZr4MMB2AiRTxuA3OY8Zgz6nOLJHn1MWM1XYiS1APa42F8gPirf2
jEbr2vkh6KEu/a1WdO+rR/G5UXT9gL6L4Gfo4YMgar1lvcLOOD8LN+bg2aUGPpIu
dwPkqSHvR2mczukUvBZJBAl5FR6i1uH4lXNFD2DQi25vSsDIJCU1o4zDcsLAs76C
6sAE/0Mi8q9lXj3h7BSBfAvtaKLtOv0kbqbc3wG22veNS4hGATP3jfDsQHa5JXdQ
4V8X86ySiUqb5G6HAs+xrimBY5IG+rBuUsq+4DeKTv2GoBsEb41C79enHXRpfD4b
Ao9D0jXMSWzavKVI+lR8W2yMdsU0r/C7S382wtanKS88kgzGkQFcm2X0QNyntMd/
CQ3SIoHhnEn0ctNlqcIc0s/8szvVVR8qDFH7Fos7qgSxa91IN4EoWxJH/91YpSYx
WOwCUeaDQuXNz6wWv9d+uvG1O3rhqD5mDEA1uE3oq6M8Zoo+UA8lwKPpdbWcyAue
BduQH1+1Nwfu8E9upnONjPb40Bn4GN5zwye/BWHzwh96FnLIEjYApZRyePOyFgCl
pWtYMaltXgnRLjqS0NodkmP+zeFfiiSLGzcdTFEpC77DOsx6BX5KsFyPne/Yac4O
U9d39s4O26L78+7MhY/TqXk0CW4Vu7elrY5vB40hIvvbA8CMrkmEdJ5HlTKPOIFW
G63NFTH4Im16jnt0/LCMMOMZsyW3SCJsninqvVCBHbUUeOgngw74j0Tp02UB2H8N
MIDcNDGbK++Usj1jjZX2exQz/MFQgQYzGjVJWwNauL8GTmKkt/kQemTF7zVYsOz2
7z2o5PT/ezwFSDchOTChIG6njMrBfQ+lEaqL7ocl3P1K4cvyeLtnM5zMg8SJXoRv
qg0C75EdMnxUHFGZkmF36OMdzNB0y/V4FTU4D/rylP6y+d8Rxf4YkXdbNym3n/Qm
Jsiw/0djJLZHPnbooEFYRW3kCkcal6IWbwa6vKdODnefJVXJ/d34EIIRpZP8+jcR
sm8X0E3Ctl2fVPWmPwRdtO/fq7+1mK6rGy+bTFx9w5xEUtcc/o8c089rEdpgiYOh
UURnBodIEhOdnyc4SAqFxHDs2CQBu1+qWHveIS7Q/Id1keFBRa+8ZBkRJ0BJrDRH
299sFfwo0yOZH2H+WKGhfpZvC2OsJBjAvS/G1phMvaaRGD0HKIv9VtnUwOtWwGG3
56WVIxhhoaJ8TUD25ttXXNwsxteSxqq+2xlEWNK6R743pBoOdM0PZaLJh0xt6zvZ
IKf1pPgNaNqg4Kb+lznqmfuYMgnYSCeaURJb9VWDZmvsPC5ggwv9rQJ3PbacCwH9
mcbSXtSxc5B11ufKyHgms/EVJPpHrde4u4yMzeEAJe1mJduKUIzQt/lxAAurCHAa
PXU3CjLkm6G7qsoEr+TtBcmsxNMWAxlJHxgAM9ePYvpTRmqiqXb1QxCuKk6ijKWp
h2xEAZACrbikCyHKf2mQJcAT0bIZUXsJbYObyWtlO1FKz10nnmr6kFALFY96pL83
BTVzs1Xnu4YE6QC2zKhYASEyTYtfIJOG7zK6NZdL1RAX6ty92SHpj3GHp4PSyT+j
b8vJjuFF3hJqv3WuU4/6YCcWCVbga3AgxiUBasXaDGglr2VRdIOr9OXzPBQZHXuA
lPGn7ABeIscHRAqZGbg7Xfk/Gh0YyxfjVwVdUfpYr+zPyVYYIl84F+DU4AsG8V4+
+dw+W8d3RGQONzxS+sQZICN6C2bNy50lOUcF2p1r0DWGbmJzM5vjAVdsAugbXCxa
bDKYU6jCc/SHh9vo+tvJvmp0+cw2z5GF1qM9ZJp2bIYFKZmQQDKuNJ+6BYhpIW9H
fCmke/iQ22vH92XvKI7LEY7wUaMk+HTUeiUgrmcUXVoD8oVPL5ROMXtO7ewTWagM
vKnzkcMCpHx3pw1z+K0rMBayQ0XXBT+NpY1opwZGa7HWzUmF1ybN3AroDnc6riTN
70wmPC2jZc8zgcXj4HtWfYtR7FqH0fysD4JRGnosdX/ajTGELu2+0NndwonKUjvK
n5uF3pFNBmJ10lnzZBaFEMNaQ8rkAIEQQzD8fkxOPgwuxu/h+0YQ50MAzJ9njrRL
FkPop2SEeEm3rS8KKcniFBdmx2Y7A+kGsIcxcO1JRQi0Ss/cMyQ8XzucQLymlkhy
jXQEy77NDjvuGUGAukBDyu2xwTuULXNwsnK+m6fJovL4/wMLicBfu3szp5r33m6Z
TP6HfG8mUd9R4crKHkfPPr7mTPCjBpe1DU9aVioMEsHBHUgaImSaUE0OUzPHlZ+t
FPCvbPL36/CALN0T9lRPSlc838Nd+uhwq/3dHlJF5cvApRy8N2w6Ee1VNtJt+tvj
hNBx7X/dPTB+wtyikmEhslRhC+QuXiCsPMVkBkUR4rO1XcL26vXPDY0UFCh87Kq3
lmM8QGOGRquCiHsCgN7aaiERJ+PZvSmKUbr4R8LcrQPr/qHxeV9jv+ZGUUbRrWTT
ckZ81+f5QQ/RDXRlYhhZeQhtDVKhw9zoepzWX8mAQku9yYpnl6/8bOwp15No7eyw
I9t6EXxWrk0Q92nJIIrgxi7yHRFoltdl6EK+rEw6nEx+5QsjvyP8jAX2uqnIWS+4
8tpk23O+g0H1GJy7PjmgeUDEao6P3hB5HLqP9BnnkE1Z52lortNiONB98ljvRo9v
iJYrXzn0fhrmeMdgyxH5QaA8x1zlToqt95MEvhuLsIR2OuahoEdokmN/V6cuLb2O
YttTjPt5VBTT5xSXCpHN10OUt4iCdkPllvbGC3ZzCLbIc6APgCv+GTx5Y9h1wbbq
obEV/o1mmciP6IlK51mDmncWJwobglDNXcWP3TgGL1BQTbew///V4s3XrqJQopoi
kxJ4qZ7OFACzbRaYv6FvuzLOZmJZvedWueGiitXm0tBVwQ/7+eGe5PyZzMWaEhTz
W3ESabXNlKr0A+qRK9bzgcT7Zrk31aN2NwGlXCdB6Yzgvgy4B+ZXxrDPPnaMlHK6
tUrjq9EQd7ciputzmgjFlnxSaesXttqMMEnJOUXqs+DK6Y1OcqTH+y1MOiBlBFnt
j8nLEEKGTSpolMZnzRmCsgbZznuGm4gWr5PHBK2m9z1IidcS8A2Ogdb3RThZa3b5
AmD/HksTIUE2U2dPnqjAPxOUl0bxAAnvb9LqGausnNMZH/O9+3nmT1PcIh2xFKPa
NZSek70zNZAt/eGmfLx0eeS1VRrpu2jwaWHyIwa0AioR7DkdxkRJzgPIc9Nh4BAK
hqLc3GcWX/D/WCo7ca62d73pv9nMyPlt4w4TKV7tgkGn7L6PWDCBXbDNnqAgnH3L
AVF3w8ZR1oZccnO42DKP/6TQ5d5w62f+mUCZbw6lTW4jh0/0YYcXT93yRooG0oh+
lFWEXtsC7JbqdKYP13v/oJiH3Y6sc87qfvjjFY1wNsWqWrMR6iSa8CfgUANVfsKi
5le/Yo0CwA8cLhzAagdueiZn7laWll2fKDa9AC6FqI18JfwiZ92mMWhAAphV8nc+
k5HKfNh4tLuBpU1eOq7FU6s9+uSAOQz7NxbDDkdd1wYoLwCfIpZoySFuFuz22UBJ
zfjMuzWCGguMtFGR0lU5pxkv9jC3ziGW1Usw+7s2LOINkUJseIAhzsyQUk5D6lnD
BanSXrXT/jtEqqCRMNNAI/1q/1NdJ+jgUEPc4Xn0WrO9pvK70rAOrcr7tgHgH6I4
tQTPX0Y/0rTfABS6bKFuwzmtbOjRH7017wf6mHrYBpobAIGbOZfP1Pun0NfizCS7
pukHDyd/9UxMSdWn9i+4kMmO9wpmVONZjEvA+1/rqhBCa2A18tsXqJSU7JvIN3U8
5CcGZz+AK0Oe1ELNJ/krsm9CFbmniijKL3AZBJ/7oSE2E+8Lana5zwlDRnljlU9U
BOAnLns1uyYZocZYm9LTLvwGcx2y9VOz/KJmOFAAO54F6uOxIX69G4DPHZbSjgen
Km+c4QL+PU3TMwpGTKEZSSfIslcQKrfPXyoeSn2GfDMz+ifaJgYasHOippxTf1Fv
Rg0YQ7Fl1ot3vp4YKt5iBZZvxh+LwNHZOv5zQvb8WnJ1ezMF4akjLA+/r4wdc+Bd
NjqblgPY5e+cWkEMnE48dCh96pdDfSeF6NJ/pVPsfuJpqrmbqaZ/+LVUzPQbf1q6
4L5tELuauB5Wu/AXEk1gW/nxgyXOvu0ilVaw55pTaX0H7AOwrpSnPArdY8PlBAMs
JgJGfm6gs7fR30agfXBcgu+F5elPdV2MIQFYYk50WfiJWOKibVxdvPei3oVSNIan
HhvVLR9LDhl93OXPQB4RK9TgYGnNGbvd7MKulfbbeiGE3L9w8M/ae4bfIul+xVpE
bPZJUxiPCgZ7FKpBDutvyHj7zFwp6+kSzgGwIHv3JNttt2RnnfDHPR07umAHsEgn
Rl+aMDV9utBoDpPm68+q1+OZ3mXn8RZVki5khdzfHgLZ+Vn3g/J1UuNCvdYQIU+t
1yf+ztps8IdTikhs068dRMdONJTXY4fLPvqCUOZ3/kgKGTJoImghlrBGHr1QUUys
9M1fMUcMKc8E5Csl9aaU/dQXlA2H22bF1RxM8ZcmLx9XTzU4nFIjar2N8/W6yh8W
orJwFqbuUGVk/yJ0oIT9kd7IwL8Jx5hLUGPNEP4+j8K46I+zS3eqfkLQFdeaW3Z5
p8eNc81iouxCZMNyPNfF91OPBcl5QiDG/fWJIC2tD5IRwrr23lcCqSs34+PoGyrL
gscuJjGhjIfTfwb33BVyJJB366ndayDM4kRpRb7AMNB3S6P0p2/SIIW49B18T80q
C3IF6lZrBzQ2eduZw7ioW/TaxT6Uw9bl3hxvLYHLj8Fsed4QCzforCwOSN1+yCvq
cmHG4IclrJfJGnJYipyVKTIhVUIpM7CXWd9DBaANmlEPdYg+PjlliOohVIPzbM+U
hxjmJZ2QI2szCqUMvxvuMrYi4TnJ/Cqju3pdLdwVF6inrtptH2Ki7oeh1ERsg0y1
enJj0adFOgSCAUKwGoJbBXZSWwALJatzBZPNFNlfofd/cco2c4TyHj/wQY61pizB
fXPApu48XxOETr3rxACw/q7JKtVr6XIILeF0mslHDTFhaDdD6oeLCcfSRRLwpxBy
91ld4Nfm44LLrFNIyOnZnuL+4HFObvguUw26+5mxETk5Asd9FPgaBNA1uejgvksN
siBNrSpK6CGWdYAwBkA1zTMRq+y/4RkpPHrz7DzDvH5f8ZCqCI/CEzzJjWmrSwtW
irPY0tuyyMq9TN1kAPslU2Mp6I8XFSneENAhIbrzelc5sDBrfSRxKlKZ4XzgCZtL
5wsR9ESVpb3S3Wt2CeKJLv6Y9xDaLmVZjYZ1OEwwUdEfF/lEYj1ciY4v68+CnHzd
Ti0zitUaeS+3SVpAR23FZztze5/wjCrsSbKu29JJ5stpN9K4slFnqkVFViGGRI8J
Xo1isFxtHe3XjzFuVQOaZYzmH0zcs/PLWXAblFmI7Rs+Vv6M4zucxOBCnC8XG5v6
d7wXY7O4qJjCUh+5cPFvmi+i/jjXTrd25rQ+8J4Exeu8grupJX43XtW/iolfNN3S
RP5jsdvHnhz5a1SV4WQM5FawUf7YnomJEs1Iv7mM0beFLkAEFHwVMuJL3Znda6VZ
VrRh4P/YttSm4wLE0gB36krIChJuznDg/2xbf8RPAaL/hYw5CuUA2EYy/vdfQ1W2
2sP/2/DE1w6leFCIlx3tpVKT9T0V4JVVmbcJwNqfwovT97FRgGiGgDYs38AkudPL
9W6rYjb19WRm6+EE0JIjwVqNzom1kS9Dg4jxps0PhIhRUul2BGBj5X93mPyRVp0b
gZcEmcqyIjJxTgsj/gSyEFXcVY0OmMdAn7j8Hau4B9fl7oebxGyOFq/1yxFaL4h6
BvWjysX2WaUn9eK+JPc8O93GkM7WnzAH83s4Vajl/ajZ7ykC6TZdbX2EJTlBJNsp
1lVHz+h18f3zchR+3T0i10Oo2H8dlTWE48cTlr4QI9YMnkokJ8RgtxlGHFJoi7WL
/s54yvLamvJS7gJogBv8/wizt/QUN6uAlW8pzDgnrx/Qh8BuEGIH8/eQhB02jEbt
FpJ7BVK4qHgdvYqukL/sM/WAFUNUBsGk8RC8pv6uMvGqWIaZHSUuTfYEtGPTz1pM
W+cH+zufbHKB2hv6Vln5CJAMg0pYeSgssGlAynorQFOjvb5mhUYmbYb08Z4Wcf5J
gvltz/Vn8Br+edaj9G/lddUMdEuAWS++8uw/G9S1nCBniU+cP4GN60OqbkMv8C56
wXBClu7CTwRLOrrhF8Zzwh1FLhGZCiDiORpAwBKYN9mR5ny3De4QH+Uaq0G3mLtI
/6PFOOojWO170MDsbiNMJGyqkyjhDLpPdELdsuYXga/cs6sGs2s/vxuYCZmoCETl
7nQ1TJrrRaHTt/SoPD2WVRrI7Ef0kgfxPtpvT31ewz7TS0vzz+GwP2Uqbj3NK3np
zuPiQxI6kdvVgMFLVfq5zc4D6C7kLaZr5KB3K5G0wuSeBMDpeMpDWxUafXRpE6L5
pBWDqH4dJMGiX/bsO6Qmer5AL+SXfZd1qk4gHFZGSY9fyQvMWxfsT+Z5E/Urq/fx
w7uSzmvLArupJ1qGup8c2t365Zlo3fWAK57HJizuPRdfKp5Dn6ijHRTsaomMyRv9
UPrTmOBbZRbCTbT7iZcLO7MErUdMGdf9X6Ja8gh/+AliypZo5fJOW33NV6swTvnk
BDd99fQsNh/7FhvK77VE96z6xDtfpdYbSPBnDv9g7eBkds+WOlnMqzQPDhP80xsh
hAavSHfQamnWz2ZPq1IFSasIkqnCmxdQe9AEt1RVVlb75w7JMTnvTygh7AEbyO86
g4Pp0NQTqI5y6H6q7YIIURt25XGRECJmdMT7rAvI0eOVlbrnqYcS0JexmOb2fylY
vNdK+IuL/QOyehQeEC8lo09S+M7ziF5Xr0k/huPXL4B9/Dk8ILPFCtbvWHLryfKq
2YSnA5GKLBFSepG6x2tXzZVouPY9l2f/IbDVzdPQmgZMV7Jss30qGn3Uq+a37OfQ
SrEXG0i8GJFidZCpuOQl5BXVQ5GhbmYhWUDaiD0/rIGtW/U2M3Ynn+o/JW9fRkIX
n09zMHr69lTA3FgAdQLoeLueNSANcp0cm0ssDW+zpZhdN9gpQDbsx846yjbnWsqn
JQPC0mWZn6ANM429i8f8TljXAbeC90MUQR9MI3XG60dnH8MTvQ6CeZvTMMwDeyKF
ZxGxwBEEqAzs/HcNI7+yvGBIHHyWtL3/Bqp5Bx7nniV6nFV1452Jrc2ShKriBNKp
hdOVrq4wkCuWjKKCGoVB11dLiacNw16KPKfOlqIc/UP7dYAWifg2yXSQ2HwORaiS
UUgubO73LVOJhJ8LTCxg8hHE4gR7KTIF4tWl75KHKcSaookJxrV0nw7BUWff0zD/
/7pkN+GVD261ly15iqJeJJIH7fzWANrZi9gYAO5H7vQtRMstan7N1CnnFrwr31Bg
TP98zBO6AdCOuwfcqGWFCEa/YdZvI65MtcJQh9kWu/38+Kd2UKSTJuvQrxTCa+Ca
Ya2tEjjm/wkohNso5bne8TJ4IgIdcyrlqiisyLt1uijgHAMxZummrclk3acqWtiO
Z5/ZXCGWU4FEFWzfP/UZNNJKxVKrarRo4n9TceaUgl+Gk3TnlfzwPl8rDc/66+B+
iTOoYnNZEZxtKth/74URN36hGXKyIHLsxa/my1HEcCizrkCqmXmi6fRVIBgAQxQg
u2zoE8P53GAmlxIciDknJ7/WdgBRxmicks+wEUy3NLwyAW8q5zMIpFpj8hUlJbG0
r8TP7RgPNy3da5q7+23FqNXIWFJesGzFTYlharyqRCYCKswWEBwicNJYpAbKQ3/n
pWbvjiKnqwXOINqMFDGwlBhUkVkyWmcOzazXpCjRfMGkNwgOqhB9/2fdw2FzSYS7
VPsNoyBkFyNWFlzhRe8lEZIArnh1TDwKLRRRrd7MSFkScMQLsdoA1RL/oZkoANrh
hAQimuK43jBEClx56/rd/OnrFK7G0mEAEG4CkGGV4hkkm1sdfH+TygTalJ2KihT0
+U+S77CUz04hXjNdk14YHwQwwxPn5kfF5TX2TQUnEhMTU2LFdmYH4g4iijenjSoq
ZxujaK4eMGILgoMvLCgYwb9H/C/KZxPixFDkcogVni8FaDlIzzp1Ko4m4+kNHWD7
++qO+nwKR0HLEFZRm1YWgv7gAyR+JAyoTfao0xun6aPvw/wFcZxUQqBI3HWzkYbh
GJW1evQ73fHzuLPEJjHIxFLWi4wkwrPC5NQ8KA0r8L/ioJu4Wu6HkxKiXxR32Kny
VqOuUXQb0/eMrBQhirmEsjM1i0bmGoRWnOUooLkmSDM9uhn3MyeYbLFJZloCpwjf
CJP97I0g/uk5Y0ES5XrIdBqc2PmvajU6TU03SJdZAlsUCILfPn0KUtkhRRJttcfN
EHGMn9F736K9lFBRDIkFtkLLsBLIp80WmFhLN5kHNrM+6QLbholPkeE4Tb3wA+sB
3N4mhkpzSQmGfHOQQxf499MLfR7VuDfuw4XePg/Ah0W4+fibycAEonD+0/QSxIsv
TpbueQ+Ln7Z2mF5i+m+svE8CgASm3XRP6fDqp7u7AmcP6XRggnQTy0cxNQMCuujv
NIZM0vYPHxbdzJhCFs2h/cvIbkQRn7a2tS+sc2+Dsb4CPJzpWI1PY/p1qJxuBciX
CmbczZAcoGv2yf4pvgAs4vMBzPZXR9e4G5q45mH26YR9L+lra+HyCTNcZMbjXQtl
u2n1Gjjhmf5N19JxIJd2+QeS6nZ97Ek28nVKwI+s5JWNDPeBmnm7k+lUFDNbSUl4
c3hJ3BOJZGQqf1+hAsz937eY+ulNBKYLC9YXfCJohT4BfZYh9InFh3XCGVJTZ4Of
0MQl06Mj+XAhNbfxcGFpegBAIyndJm4fqYJAML+2laSDslsXY7es0jOEr1/Y68S0
Tcsy0nrNEuqv+0Zssutjce+odruXkYEN9WXdW8I6xiaKd3U/rMeXGobucbE5K4IZ
IcMoEz/safklMHx/bi7JDo5XO1QIt7ImzzPy0K5lpo8fERCinOevNlhqp99hU1Ms
dW7g/MZrKZ4bP2wunUov0WglieTyIJ26HZ/B1EahKVdOvFqiM9tLyQaWI1cTtpHd
cGGLKbU+CuadhScyphbY4Ur5y4ZuE3d9vzeGH9H2Vz0Xp8HIlW6D/3fIyyLrktsQ
wqRTJ41AJ90ftgzT0AQttmhUcldg/CTPHUOlfFw9u703Fa1YEYQ04LBXw0GzvG1V
aCNEfYs9NfRwoFA72Nowu+Mpb100+3SjsGle2XL7rmFKT21kXdLqvvsHT7f1UjiY
n3DEiaXvQMUs8MbAvtyjnwoF1nXu6LJaiXyy36V9m1F7JNojgn1SSRS91N+EqhaB
NlzudIG7kNBZ967aEB+4DB51R7I7htjwlzF2/9gqVPSXYpLvfh1CW+BF3lRKU85k
gLw+03ki7lakHbnsJYuHhn6DUqxS+G/dXxlDCDbEO7HHxk/PVB2bMcw2vL7ah/jx
kfjBqc5Qu/1rqMM2ZoiDdh9TrJEsTB3O3TAnnNw3o2IKel/HLPgw5xxXqQp7P3vk
Veu1uMimKeO3WbJnhINPynSHR02Bpu1HBPZ3fNrLp2laNbV4mSKZ6AwJtR6IGiqe
aGsrmGInIoUCzpE5eQ3t1aEKH/6YFtnsQOsdyeMd6lNK5pNg+uRNK70LlnDYEFBO
bavmwSlNV8/3PE8e+Kdvjr2q7AqDomveNdYQU7ojs1WlutNtoQ4qWaIFUOQ4D4OW
7cw1JNpABhOhw2wKrwSUR9adYoWcFDypZQzGn2vPU2q8r0ppqD2DMkz+3klo4DDe
eFjcrGPVXFc27UVXRBKsJe9O8UeiyPSmMarpTeeTM8JS3jf8QWp1R5/5uixGmYg/
ty3eButS09mbIElZDgw1lrsrJ4H9Dp+RTg8oLu9hIIEPfjfTLcrIQ779BTO3IQx+
9HiYYqK+vHjgJMyE6VeMLy4ojWtn2U+dtimlcRhsByo7DJ9KOFSxavC/AyfkWZQj
HWjeD9cjMyC8QPlFTxwyTqSTPw97ZMgKoXDhyOb530o4te2rfhIwt43CSWYMvYZ6
iROH0ImCAgh3QVUvRf1M1K/9mFjD4URJDeAJXj9iMLwyL8C5Z1MgXJpi2QqLX8z5
gKg9vDa1XQKWPmpzc29gIsQQq9IcxIQ3W3KTzvnwm40a/FceN9rm0On6SWKjQNq6
QZHvtwnsfWdq9expruMPJHPKKp/t/L45liwQlRonRqyek/cdcXz4VgPpkWeYMF1M
VlFPAq9N6+PBvlva4ltr4qeNBnhrhN3Br1K8ohLSAKV7LoNrSKtzPnz01O01Plki
uTLCImIh+fsXOOYFMe6OrBOlYEuDzhnH7bGX0TCFH27NqfPeFNRMAZNzZ7I0Pd8F
ZE6hdqk/Qb3v2TKC08SRAHKnn+roUoXkz/IVWbJghyfjrYYiD+4dxALUpRngZ99e
36GgcSf/AsSxsYqRXm2PWmyE2JtiE0q4ZQd3FQJ1dCkDTCAWwfDeL83XmMFSITKA
tJdaaMxdGj0epMoSh9etp4r7FGwwmJ4jkmpyxhJKAUWWOs4B4veGspAqPG/xm57d
dj/AEN9kFYXTRkqNLFrYA0Om+VdvpAVlKylLZ8cyTdyoT0lT+M9NM1BzomznD3lc
Ab6xAjNcxWymPqiQcqR1AAOUUddBCBG3Arj0Y/8MFDH3FmGaY/RWsL8WNlbqUR1i
1nQhTARsSeIi0drhsuqGr6vRqQhNE2p3XUexE1omFUSrlJMdSP1BTw+0D2mWtZD6
kgG7ES2ijkzj+sGn+z0BZjdQQjwoJPen2UETOUquzqFLC6lrSd0h1ouGrezlQQXq
5Wpc5oLxZUHGuQb0G/dQEj/tfUCX+Ltktav57d3QJyNVqaZTCpsMHC0GaZAz7O/z
JfIc6Cj2VTt4wYQmDxRKLkrK10OVThDZdUhzOkNhrGNP7/ohkdIRiRm3E+agEiow
aNxWJbZDAC4/8FbSRx5dpy24TjIN9wFz3W5JqycKB6ImiXWgvoATdFkrren82VFX
VhYcaP067sTJlNcb435HNJ6iVydWl6NOyXMDgb6f6R/U3XO/k7gOygjSUdOcS/mB
tUIfi/wqd4xuiJgEBXoBfyPhkfXIiw6QmPQPvrgSQEJq7VA2lrsnd/0S8VBfrsib
z2ZxrAp1/UWf/YbR/Vs8oNX84fa81yHg+r3FTZwkpriBf7JrB7PfG9zdRUf/5Bnh
c0FZzLluMtiDR0q3ZdQTCuw1UKBQ1UsP7ek6RhKvudCDOHEnowqbh+zEUJdu0WCJ
qEdDB3CcAdyWSrODvlEkuO+sErGpNr1+S/yCLfCejsRkJBFKIHJjpUu0k8YkUtEY
DmpHlYbqmVOBRzv2cbbGduetvoncPzSGVe5tftiHB9HIutcFzXYbPoI5wMLWIAC2
vAmjoZxNhdVaxs1JOlB+72LdiWgloHJf+rBxnh8WxQDK7bqhwy0sbphQXUjuyha2
tiS8Tp5uc1DfliOMOcnrkd4oTkVeTPygSEXeIMOgTMsT/UzMKiIbX+efsTysN13C
teXDh6pcb8YCuzsQqHL8tR+pILIpLYHAXEJHJiaUlhO0cOBHGiTqGLJkCKb8GbCB
yPjR2EYKzObs5EtSADiI70hSEALqnWMsENLQydfmsbSPYF04YaZr3VWZRkvYa4ws
xhW3w20cN0dncC7luuEqjf4TIlGc2I8OJy0bcIZlIKwj9jZ2+8YdAbihIg02Dc6j
jTR3dLy5k37eqCOVOZXTI2IOwFUrbZHv3mBZJLGEBW6fhQd4GktEvRoLFGNjA8jL
QUtAtFZLyuNb4nw3akgwnjk3k54U5fxqTiY5vlwYF/pmEqZhJYPPuNqFMTO2MehV
uy138PmOqL8lWHbaKpADzRPtuyIlI6lUx1noIVOQtgs9P7B+kSvYIJg7FaJMDZiP
nvUc9NnafuxG8J7t0+M4t0Qlz+WIZuw9cALcPtoTrwTILBTTIaY0dkyAGSTZhNvW
hG8kCx0+mp24P5F1wD4cYsnGRlz2w60g4K8XC39USEUOnQh+vkEc6GAvqyVTFxS5
SLnnLVIoNLTsAhm4QHGSz+1PjdiWrk0n4PtM+P7r50IO/LdW+ctqmwy723BX1NgS
B/03WRVEhYSrK0zogjh9t2PYtP4gqhJVo/E4x6c7iXk8C+I9kfkqqcyeeFQ4pQdv
j7PRGEvDLQLI4mErEEM6jKW+23kK++4Sau0UHyq65BdvOffT13qRzn/nHLZ9h3vt
9Pk2w6zdyyXH8PMIh2mWt2lvA4QE8P+LGA8V02+Tup3THTEc9saBwnbbV2cHNB4G
adOWs8krx2uDxMQekungbxp7qVuX2KFTUTdoSF4pH6U9YmQfV5r5nJJw+FkCV5pi
9JjP+fOo4D06fs25DSSVLFp5eXSUrmqrPQEgESg5PeH39xV6bija3GvMJKGPofCb
arsJxTpojkxvC6zrp9wjEp7AxXFTf1WFoMWli2yqwTZrwmn0hPe9g2kfQ1FIe70r
rCau6t8nZkM6lHwZiwcvShUdcAkVM7cGG1uDBUnBl36rJFxCOfWP4+ilr2yXvvRM
ix46UH4/chJIKXKCtGKB7kj98hsgArxaOJUKhafcbjEDvT+BzNlmFIYjakWLiM6K
SiyF8fVJzImEmYp4gU7D0kF1Ey6m7Hora+7LpKOJNgKQdscfdkigC6Fy81rVfWXs
8seUUzLSdGX/Aot+udugxKuDbz3bmcIRAV5kqBWuqPvX4IqQuirR+++7jBK7JfE0
7cy3Sm9JXD/apFqWkRmx4jyWRG3EL7Ipdoian5fFlMYSj9mx5e3ZsQmXwUwCZEZD
ZxOJQs9OxYzGjINS485z46kYsF7nvQDDtSaU1ZvCGk+cyLeBbU0E8XqNRUXl90cU
YsSXlrRWSo7qV4kxGGE7gvY4o25zt8b1KSm7TUVtlyb69XK4VxRfoWG28SzDzbvn
hBESJKgRQJIz8a2bQa90agHTj0bNRr4W9lTM6Z9OwHqdRZUYEKP3BAAXglb4udC+
/EAY4ejEZjHUflj/Lx4bGOKZZtNVMxoVNrKW7kG8Zxp6RL1FBqroxkVgDbjyzL+Y
bv6beJa1i6ybbQpzKTPf18T+EwA2MMO10qcB8eADnTI0UbVhp53N3hJrYa+CnWDK
ccRF1BDfku1DTtY++q3Jw5SD1hv9DJmE8WmDkW9PRQJZOe3X2LCxmVcuxPXMoWzD
3Kpvgikli3Njg5bPyf4KSJjVQSpoZAGSB31csYwnYWGUUTr/kZNuwnPfeXUvsBVd
/zax/SR23vu+MOf4e3+V3oupX+CULXupwvbrax4KMJIiLisp1cmc3GvAWh6HcMmu
BwyTjn87/3HPLHyLKm3Cznq9W086aennUMAEMow6KV4vG0X3DafzH3ScAQJxHK9R
tp7JyVhXu3ak5bJ4tIzaZl7bd4tV6YYE5eEhTkbRKpkyG2JXXizRTIBvmKSO8qY/
+DspDFauJ3PIyq0KQsCJ11ri1kqS+1cyxqEiXeDL5D8xcNAgIstXx4j9ssEQUS3V
RN/584GDKfnn4b2dg69v2Xj1p064j4pSokELGWGmMRUYahBaDEEGIPF4e4578PP1
c5jtN0cZ3eHTsAH8MaKWXoTGmt87pwgK8sLPg9PmFlYFyX55StbdnHqVzan2hqIf
bov0bM0MNkuLVppEd3biRVOak95wzFKifEcrLNdExTE7Tpnl57I3EZunT4TM6SJO
Hw1naBYq4j85m/2tRUheaGPb3djNQRKrfWCWmflJeSkOhn57La8TuV+Yqcw/oeoT
nskghQN614bLPGHvvgmnGQeJoK5NcxYyaLKOH1t2pgCNt8PQK1CRH1W0OZRIdRS1
KwvL/zd5r6BLP9Hxf0EO3PgrdYfE2MGwcvW3OdNci/p0RwTeus1/Pa6hqEVEgfDf
9BQzGdIegxxvfwfxBI9jCzDwDCzogdh0nfKEo37cFuV65fKRGSoq2ZMQtPkJFfPo
KDzEZE7XeJpeTsQQdN29ar0PqiyAs+gKs2LOO5gtaCn0yQEHM83o/+A12cMwYNoY
UvYjUyADyMlWcY0zG4xnvUqo7vnHfPgGpKdPi0bVs4oxhLp/qBv1boIL9Y+O/Ho+
Z6e5OD2ZrzNIiGajYTi/TdQ+MW28Q0HWEiEa9N7orsKxt3cXcApvd3JnY4JMI5AS
UI+Ei1/DjchTy0VV5FYQgX6oBgkXRFS0PFOz7zqWJ5+DS1jPyn6vRfhaFkaT1ME+
6b0EwNs4Q7Ba3Np9W+T5l5kKbd05hQ/SspBCO5ozLaf72bPnvgX0sK5pObyoRvki
T0eWfT5Q8/JtZ3kgcOkm/0kmBzOB+YSFXLf4sDWKNCM1zBsGeY6xabvGSfNTYpnz
r7zhTLodCyAdk8oEsOofYa+rUmNmhFQF1Do9z6t6pWI4IPVSTU7Xqi28xHds9kFi
uW7zCG3pCJIrC1Zmdw5kPG7h/gNrmi4Q2yEtg6SnHRrAogm/XgRW5Bfmr4G9jOmL
OSLpA1tMWEFgsuBQ70AZGdL0VNChYYz/eiXQHk+a9TE11qOM4dyRmZOjfUFmeOc+
Hnv/ihLgIIB9fhQwKHQNGqHjlRwnNsA+jeXMQ5m4+xnRmwrJrY9aO8w4p8DFRgTy
76r+jkrECv3hE61Fc5Xo3jsNESYsN9Kxsi/2GUq62xTVqZAEI/VRkomSFiMcAxf3
mwiG9fbcmlHdPum4SXQ+IUyBH7dINxwbpTGnMtLE2yRJ/WeCR8Hcz8rFn1JTh8ZS
R0jd0yBTPAGbrdcqMSlkVoS/GiOuewRjWwZAEe6JdOJ2JkfQm9JzUZcbokjsi7x4
s/EaNYIHvi9jR4+N3FcZztLehfKDtVGcIQtF8aTs/AQ3m1FCy4TqqnnzJX+MWiBW
V3iftlxNeNGrpGZpN3B6Zbt0qaD3+yalcFD8lzKLNBVMB+2lBqfkzBPk6COuHQQI
VBzZan/dicdYDvUU7dzpdDaceGE/OTAS/PB718anRkiZ8jxFRFPe2O3ryk9Q/DtV
e7BfG+FBPLVUSH6T9OYPF8AadB5IQvzK++1nQSxE+75T5KoRTv3ll1maSV09loxl
xy77NWDV+XIHRInz5fe6Y6vE0aAfW5acNDUaKuB8qPcO/tNdxBgJ35/WAqKYGa/X
pNYkcahl2mxSr0vFiZxT0FLN3wYN3fV7VEQPtV53UTVOIG80B6Cz8WuGeVeYBMUw
ZSB86UtwwjzBxQaw0SyZb71hGpTJPCvUYY/VVHzEvhHHsjtED+DhlJopmLda92cM
ixJwJUsASkjXNBmyAwS36TtjIFmtI65e14TPFjFDRORcgq8Nq7J0h0WQ6D+eSeeD
qh9ETTlS45bOzuqeZ4rZGM6YE7aRGxk01sI7fmD5AHEWHbWR01Jx76L7cMQziCiD
dh+ZwD1X3DXJUlszF5XF/QyJVTZbDcTa4gjjW1iAJCDZdNmQYyUmUA+PB8u0c9Wi
+VSNUOIEvGqi/kX3Z7rnGjpQleFgyaQu6036o9fK8ZE+8/fQJVlFW6fu9zWfWePF
sGBhbZ6v3pi0vktBn+hGMX0fCvIF8mgA+02wa3fcRJmhXSTjUHSzpW+oESl5Sfeb
NuwJMpdrKYxiBkputVCjlOM04mtUqFpikpQ4RGYmwc/hM4jOZClsOYCFObYS7XcK
LJrsfmoMK0c1NKXGK/iv+HURfMCn8irZa6RGYXCmFdG7n+2x2v2ufnc6E7YIhP1I
Fkh0l8ZB7J7HY3trl96T6CHDgaP/YUxQlCTlxyh7GGdgTicxjKTZ56qYO9PSbelM
jPNAqFjO6FbVoSSZstYnpa0sa6eTBzeWEDBC3mT6dwy7J55TAxFln+V+YRq4yXGo
e5d+YMd3gokhyBUOzwdmPKeDFDUuxgpKhoHS4VU71lvdyCkoPAvH/Z955yrDxmaH
T+hh7aMTEw+ZAEylvaw2pwrDZNBuRkcYJ6QEYjMlzoi/Jf3dw2N15JiBwusvUlwq
gRqPV/MkUKshKL4u3Iw9klj+fnZCr1XJK46hrQGWGY4QVZvxDk4gWLcbvDwfvGxJ
y7bX4ZErSxM19PwEonflfgg8ZlZdwTWtqaFFv7n9NYC/SyOKpYhyB78kOyVsq3/N
7ovGDXyYu9TvXy41Ll2Q4OSO8dk0i7/U8W7BoFRt+ynbD+dJonf2TWGO3pCOHQle
UpYNHDh5JuqXDn6AdMswsRhxlPM7Py+mrdGxaajKzVe8Bi0aY8SWgQZBeahlVzHo
TVu8hCda8zv0Ps9kzlhFE84EataqKmF/Slz69sh8YEZK30RUmOCgB2V/zAcUaTEI
un2zo2GEzXu5VgU9N7ApWv1y9ir0Gz7rs8fJXLyTuaS0D4m7dNy1W8XDy/kN3FPl
qXuKcM/J2MDG7HuDa9MMwrbdDwniIetAXpVjhg20Uux7lUk0cuVkDZBfsaRuMGbz
1vdQwpOPCcpNrhgyY5qAsrgA/cgQf16AlhQZJ9y0xmEfmQ/ma+QEZeoid1bGhG/G
V4EnvVpmYYmTXt23L7ZVs1uYscc+N4PunIyflw76nxAtPK0rHBxECP5FFlYFYJpg
kvM2TnaVMzuHyLtDVwLwKejrsM4zGiWSj2TR1twUJ+qy4SSz6Bo0enUDIT2NAP2Y
0uWyJdUtMfQcHsF9A2ADT49C5JH1rF8FQ7txW85/BhKmDM85ZD2zUsYVtgv7qbqg
3hbGC4O9q0v+2K9YG6nENNRkl06tmDNo8WivJQIYzmetLHAOkbr6qjnrMxt3a4i0
b6+sHbwXgKuWayD+2krWlk1mttW1YRmAdCl6V3vmvI2Wx8Cqmoij/GuP8DE837sa
85Zaw86pw6Gg0z/+rUaibGYhgx/vaQsLc95MVVJ6mDB1ihadOzF6OV3Bh7NSgKiY
dBDF5dQiw2Sunw1dzsCARzT4+T9aM46ImiOzUAgZagYZwWhdQH+h7DjkZtLj5aBK
NtiVdInzgdabM7d5ovR8hRTb7O030hY6HVxuZ1e0n0oEvPcxlBRfwIlqVPegF3XU
Ilh2b0foU9c8B9j1G/MR+R5g7Elk7K3Wd70GYbyR28vjjpIfA43Wp9I5ydidi5MX
gMoQf6wkDu+qHFqjp/VYM0R+tCj8y6Aw45NsGAI6tL2a3s+Y/pBghZe0jID88QHm
mhbQi9EI3kMMBRDlmb6B7hlXsEi52qV5NNU1bkgjqcR+VLW2quP0LObq0r8jEe/N
Nuby03hHD7K21fhnEIKI5pRj1pZF3bzZu8z94T6k1+R97hxxAHctu5yDpDMWxyl6
0Q3y9uAGMg2Otj38VFzvVAzDyQu8BBsWh1scySF/es7++8oRw76QSpSGM4SU5Zbd
q/6VwHgXzgufSnvirZPXU7dcJvT5lISW2luBKbSg+AZNdvPhSD+UstAIsClcukTn
VCkmWQ1n3w+feBgCluve6meeaxRxCDTJzoKYaJrThPZPhd4rtmsQ6K845NVM0GyU
Kf3YN6fNLPe1+pSf9oCGU429P2ANTt0oNjq4EJhzEt1Ihy7auNOH1uB+uHisdbHX
oHldkfKYPs73mwQdbIs9ZGjbgQqM7L9kwdTwSRQoGrfDvpqMOznv1cplgulpxxcK
Av7PknlaQbaDN0QiBfAe70I+TpOG1Nja85tvfKbITumFMf6jbzi+k05gyeXO/IUm
v7MsAYHzWsYtrEPwduuvHYhF+4BK20S7widWgApDHuVlFXRB4rX/wFkKHKKPJNHt
LE1/foWkkyQdRTqMgsZgsVnwCTsyYz+99m0ZhzU5LpWx9D8VXRM/5dhTAoo02x2j
DjISuKy7lJAGCf96mNuMYNGSsff+8uTr57SBoeNDQiXK6o9z6OHaN9ZUxGkNPBN1
ZoexVCRtB06qSZVP4W17dwgS9Ojq0pbZifyU25TmJs2wuXtM3vDq3Xmcexem1JxH
r6DMJrsOT0gAM4VqxfbNsYLNbBkFF37A4jZjTsnmJn787M0f3Pimok4i/Qu8UTAw
qQeqPTiyuiBgYFYwu1cYr5Gb/xG5F8dEQY21Uf6ucWtME3dlZWAFAiLFp1LX4UhE
W6rR3oiX+qAMCR58icWpdKFdUPo/j3+GFcyI/fdK8yreKBUVLoY4klm2XKlJxe+J
URJvmjL6QVS4h/E9FAX3HNrZOczXQGv+lzaCCwXO4CAm04UcW5KpCanl5bcv/s32
u6QJD4sLqaLnbM7C94H1YbyDDLJ8MlAedmyg3zEeiJn7emq1Dz8alE/ap//mjm7y
EihECypb9NiEu/nYuxfyahy4b/JJYNF9iIyJY8nTdSQXnEwPWidB1v24XEKG1crW
runqL+j+NUaRl4MTvUd+Nvg/gRA4hH7VW2KtmRM8Y8zpg+aUG3rOKlei/zkq8o/S
yO30F8mKMYEciq7GFkt7fZUZN+AgcIx8vef3LoK+/Znm+UKjc8I3N24uwK7z/ymG
kpal+G/gFuuSGqC/r9oQMxuIf4i2clvo6HfBkNkaCxMOdkuJ26XqvhCZpYnJJrUD
JTzTxcxse7QOSqnX17lI0/mVaoG2/M2mXZcb4pOaxcpD3wZBkviddabBxmu4hkdo
/rfgPDfHwHbJLisnLQjB3sShnRHDGx7cZvM8kZVF8GZBLtxaJzurBC5uqKXeC1Ut
DTPOSnV8+Bka8+jexxtOC0vNZM0cB1HNq4HfJ5lhZG6bsAlS4YLJ4FPvx1WlHSNG
5GJMXEGtS+PponWnx75kyGZT0buTCn7l6YDcfQtCRRUyIejCm7Uy4XnjcOT3q98M
fWsb/RRkodo1u5WX+5+tLwSp6pK+XPRxdoCHlxR8qdLmKzo4PVxIqG2onq+NrFO6
Ho4GYfUqz0p4kZjq+3sHI4jGoUnZrCPeOhXrzlBLyfsXp0+iqxN86GaUWE8f3Dfl
dOeZE7WtPjtcVr52lwoJTW15upFzKbQc/H14NUmIjmhCea8Iy2Q6syNQwFA3Wadr
SlttkJoH70T53GEJ2EbSyO4mxQsCOyiAfK4ktg0c06nZUF5AoThWY1AgBD6Rj7FJ
EAB/YlRVnQ4YEDVpRToAO7fN5rclGqjJzrWNwnJqAGzFgnHvm5agyX98va/IjniE
As8y29FbSK68co5CROd1/a/QJaptDXtRcykAHdvoCtM2KUtmC7d3YZOotrE8HDGj
MPQ5dLOjo/vHpTxVNeW4Syyq01LwIkfQGQidISId2Txr6CGhJ3oLpl+OEZnz6pXC
Tj4gHfHJ5HJkon54YeB0J6h0xApA6uX/ox5o5wfopb2v4SVsNEGq+1glOVRhmsAC
MifdnXDT3Wm/aLQgr0gtZkXz0+FDx3rbW57CqMqnmy8Vb1RSqmBMEaqjZZkvlQJV
qecu8L+afBXPFXRmOXf7ICv2WjrchvcPzm4Srr9keDSZkBarALhURuqwTcJPe4U6
Uq4sakUUpOPQz2Hp3JvtDeer6r7coCjZsHvWnDjZbyeRJRMcL2bwXgXeSpsCH9cT
7xY6F1QY9oQFeZA+HypaORZyvtewy4yzm5g0MIQ67Sx+hAE+6n+QmkhMWSNbha70
0Q35GoEOHGdJuNO1dPoF9GhFynjJVGlTonvWXaD8t9Dxiwr2Xy4qzsqPn5bNSIaV
h149hMObhcdtebIQH4zLAdwVJvccozt9p41kzbJf+Mlf075HMoeF7I962Kfki8RK
9L9YKbu7KKcdZkEEAtbbgnlaNBB5s1t2exM+05DVEc9M2MIO8KGIfm03DRcUbG74
QYu9pCPKUNXJTLQKSiPWa2lNBAlg9QdV/IVkxWcZWxP9Ka1lsQh4rvJSg4aYyowr
6bz6HjX1yAKUOYko68buM0OJadKTL1NYcAOZDzchzWZBc4tSIs3vzEktyYF8Lr13
Omwts/tIcCxBYrz6eU9SK+V3blhLdpC0UrtfjpBGGJni2nEyDwoqKa4WPaJJiYwf
1KrlJwegXJoChyRJMdW9VyBsLB/9od0/YU5qJTVN1cHLQMMBDNlGZYOtTWhQEegR
PUCfa1qbLKIdWKZnJ3aK+HFLXIrWLWpUoDPIP/QBJ3pGkDiaBIGjh0WCfCR0uldz
pOlZxzylY1EuwLAP+kALgKf094U00VUNhMjDxXV4VTIRYVoSsbiislmCcADwxg9O
PPWJTjwUrr0MF+s8zOTlT4GT4+26tp2vuC3Lk+6RVpEfI+cgOYPsZ+rwsuXpoKsm
ClUQdqeexnrsZYNgAg5kM35eXgB2GuGp99jfdrssHJJD5GYiYHW3DEG2wetJ+hQe
3nFjvpMoBlZo/vQZjhWqHPHDk/O0rK8whN8mrUPwhur9cPbmjfNxn92hjKlJgV30
vkDMsGdcfG0kOhArEqwQ221A6wBtNAkwsAt5xn1vN7pJZMsObGhoj+0TB6daEL2e
vryJ6jHMynI5RchP4ykoB6XAgVAqGUD+wORu4cGn1KvKSnuTqnrBlzb+lvXpVPaL
C7xnlmTowATBKtM/SoKtv5HfBGc8vPPNhgVefgw7LPsxYJd3T8HGVn/zTtJ859E3
UIE6362Hr6lpIgVI/xLgmak2gCI8desfFM8fO4wC91njS9XkXWSg2HCbLrrki97p
j6kCTVj3SYVHTyMSmi1jayqH+JpIAgoqqmnYdaL0DVPTM6U8fUZRafkeABsp3kWA
70OQcsvttLVwkVkPNYBjWhEJu/20D3VAq67220EGxQ99lJ56EvesJm1n+ZtcD+P6
hX2zZbYHg3NmRzKGYitTbajnma/rdKnwYgtTapbd4vnkCJaXPafPmS71mnxMdcLI
rq9isZOL2f5eQ6Jfx7vrnWblowDO24dXRUefwtRX0ev6fQXP1URBZkYYVIqBUgX4
o6LboCUyOyZXoX3htYihMH8+z2lS+EcDAze7a3UPkh9oOruMo3HiQM/TrIJDkG9u
AKYMKuJOxo+SIw7gW+i0MBqSpB3Ut2kmnLWc10S45EPhBqR6Klm74Mh0en1e+COm
F0dILW2R6hGspFZDF5SUyUZUGt5PQJQlMLpRsGdRrmE6v+7uG/dh6ytwzkTIlcWA
4LJu1CIhusTNPJ/+Ck8k4mx1HKk0WdfBD/pabVdpALeu11itg4ENjgOLGASgRFjw
nWQxRstugv34AMwt/agtUFgxn2MiMyYbccbUTl/8sBHgdpH3rH/xpe8ZHUVqiMTW
N6uEYVI9vSUrw1ys/ipz5srRujetNiH7mMz5NGA7gJ7UYPxK3JlQOp7z5snE+qSP
FgSz1brhTxt5NZo5Zl9CKU6qEgHC//4/QW7+pVcB6VI6fGBXsBJ9Dc0+Ea21VV+i
ccb5mE8pAVZ5z7NjlKT7GD/Fs+DxF+v3a6P97VoDeV7CgrLg0h7kXVNI5dBfdv1R
jTFWI1h/Ft78K6fB+torBCn1UJm/4B+RUWOcZZJf+wra9xih+oDOXF7Fxoirstty
g1te1RiZQhgjn2vPmDUyPbolU5KOmky0HvcSQ07sIPLHhB648E45nHng6lGBkCXF
FzfmtbhesB3JOMkLULExpAe1wrJjUXQvJT0pWXmJrbIkHJJwWxF1CNrrhtAbHWnX
j0ArqPohe+urSkBLIUJLd5fNJQEPbhYpTL7jB2rVeuv2UXKiRE6IfiRef5lG1tpH
DhftUKc7a8PerXVa4ertT+5jJ58WP2Rhz1/bAfzOhO4OQwGIJWq5F5zmuzSViKGd
AdHgJR05fqBC1ilFpjeNbfLS6RHZqtb09vTwI/IR8EpdqOLhquobuccHNBnmCagq
pQO6z4Sgkl2gqKfAt5YuvZb9KCgYOYTIxGgJfcJ4ShptTkYyNx+G5AUNTWv1txHs
mlC9ZZzUo9aRO7JVoezNkwgnKVjSUzjR1GSfmMRzpklO0067+Ilvw1lF9gm93I0R
QcZpfvlsyMw7AWwcfeEAvDuMk0DQAUCRckTqpDQN96RodyfRbf5r+ggtVMHVie6h
yFx74mZOQ2KrLHoWmdOWMfpnMY2JDeNB9OGnWYeb8FgDzuJ4KaEMwY4WukDReffb
9YWE+yU4omzEBLTxPqqSdz45063IPc05fYN811VlUFprLKdKCPJcYg7j5Z0LfBL0
fcJZstmY6YiFWFolQvsUHiFpLejSO8sCe7Y3k64BEZN4cpV/dVqLm8NKbuAz3+69
JLuqKSIozL4x9u4H/Je4SpvkNgya69pYInlYgQNHblEtc0eRDkiNAjLgqimNaPTq
HfXb2PFcZ59LuswKq+aFPsypZyeCPzKo8NMkW4RkWZpt3OdgO0oOCywusGOWjFi8
aRfZhvc8oyCJ6zpSUeVx18pEk48uBmqxyAyBbYxArJgEYEvicoZc893n2sYcf0RI
1w5BIuuJRjNxd0Lr+vLm07wQMUSMf2cdBlJIM6a5gj/9/w/VRdgEG9sLruSn3S57
40y4d//3EAKgbtwqzfDCP/sOMUqEzKlEP1hoQ6DkSLOnzvMd0gHCNQUsdacnUcvS
z1t8r+J8myaM3vjG86j+B9ZJ5x8nhzE19y9awvSsOcgLFRtp/nvXFmCaQ7RTgpzE
+5TPzeq8+WqpOUzDwKxMj7do2vjAHwE13Q7fM1nM5aSX7FosmYsdLu27xiRtGv5g
lWVmqCqUCla6qMnPrrKM8rFx6Tj1MnG3ZkqsnSmijDJBfxeFVQ6x/Io48YAdF0rL
4oCGeBS6voQFeT05J83I6Q8yrJQqSfsvmERerdZDgaMogLkWxGWU77XRUpFFrrsf
WVlWyNn965FGpalkf9PX/T2WRlKbWPl3Wal11kOUzv84xJgLycMYH7WCv+bnpNoV
fUi1sC15EqQTDR0dSfYDYinp4ozPtwIDebg/bUupFcsCo00SGVifhPwr+g7EyDSn
rtHnnS6jFmQn76PgU5J8O4fMDHT6GW1w8Hb0es+lN03AmDHN4NApPpaVq7cXHDk/
Nby1oizTgk+P98UFwPEZ5zbhM1glg/zFaUSiBxjyNMHwkNiUkgtEs1NpqRaEEW7W
4RWrnrTVHN/K7i1V68xOgXACoFkcBZpBRSo7e2RwPojhaH4ocLx4wek92gvdBOAu
doi9daEDzxREBZRGo8fw9Bsm+x1ZT0UMP+l1fQ2oWqIaU4A4Pl07zgh6vzEoxFLu
xCig5/pYq6pdv/Sy1xlMejKPYK8yu34MkWCpVO/7rD+QzOoJrWBCOaiptajAuLOe
zTmznHY+XmmQpfV6qp/zXSOYa8o3lTAwuWJ6u0GcfLbWXfu9yVqgS4Gm6tv8N7DA
hta26hDvSIKdKPQ+tPwhXwgPGvH/uyVtPq0MOFGHiNTKATjVmI1HK6Ua/FpzQIWJ
ZmaMitLGHva0t5ufm4S4ONnPjk/QjC9XCbZd6t1pr7Vm3Cb0mSiE+yAhxHmMUnXr
nTauys39kuPlPINzb+lf5T5vZ/ijEhtloZ8Dl+YgEPOetP1BPC/PsoW0miF3ZgG8
xN9C7xVhqyT2gIWT56T6h0APYMaGi84MIqd//dY1s2DtViEBbECKRkHNlVmmFbKv
C/V8whAmBkEz5bFPvoZBOH4TRUncVYL4lywYAuevbwR40zB3omm0fOp4pQ8xNFRj
XScOS+pCjdgikNJyib98fNTBU9eCPHQMoNdLkM+Ed/HZdPtfa2HhecXO0L7njOeO
oEZ8ffsEGhbnNJV54zj4X3CQ2fvLtTSeyJppuwdkUafkUWoK5d4P05bZ0rxKUU1L
sCM2DPHMEsX1o7F/R6QeD6UigmSwUhAWUYHB5urJB4wPyzz0UwXtHi3W1xrWDCxE
LbPaenK3JNOPb1JgSRqjQTxJJwEKqK1ABDXUJ6E1IiqGCfXWhHUpZhGwGy3UaW/I
5TEG4jKmE5EG9flfQqu8wKY8wSX/x9VKgE4hfVyM/qzRKvDjOUHH74Z0nfIPUuP/
R/HuC3j36QFi2THONKtg/Av6oBsK/KvkCIbVnyDVFr105Px5zwKoUOtcYySAEpr7
oPfpa4ZN+5a71+xDQ+svTVqPusK/roC5QUTpgtuSmQEm+rGffgzd92UF4ZbcT7F/
4uJ217Jn8QxkZXJu4jIsv0k6BTYY5bEm6OfwGHNIO9PLhyY99KyuB6HzxO7+7NCd
pJ+lZuZbrBhZPm9/doUv92oYiecS5pXP4qQQmEiG1UkI+mN5qNLnmiXMl+6daIIr
lS2eOCaW7tdjiylqYaJ4d81aECSTl1ZD2KfSLWWTcq1rXCECULuAykaE5liBPUTW
eY7/n2ln2B7kU8CTl6YNxQThFdolmOFMOwcOMIx9an91CqPc8S3WgEHcmjNupCtQ
Af4lEKazCyGBD6TND4SosLpezD+T7wXOBTePkj4wqf+qE5vwymYT+ccXXHOmtykP
Abo8y3KutFDK9HyD5VkLqoxvsOhI8vKptKTdK7iHL1CoXzAdUZoufMo5iunTn5L5
KvnJD4XQqY0QWrbagESXi70L3nfFjV+eeMoV/lSYoFVPfgzp9IUp+s55VECegAtH
tG4J6CLPaVq1Gwrknyem/bu6co+a71Aq5t2K/VwU0mNSpA/OEMb5QGx2cNmt71Rx
Aw4LceImZjjX48XB1c+xigt0Zi4i21gz4rm0dzSxauk+xGK4XNn6yFHKsmxE/U79
anakmo/TJFRPeku3Pb60Bsx+mF7/JHB1+rbVVWJIfiPVOE6T4tHFevhW8kuUPbJ+
/dVKtUQzeo1DMQbjNpWb1JMxxrUwFUWa72NgvqpSYqpu+7le/19bcw12jB3pDxKr
Gz6xIVG3mljAnOzYYYnhQg8IuujWv6wxUJ+kBTtgIxMy0rZ6cehlzAxWdMP0poe7
WG0wHf8xOUpDGM/bTMnaHTlul2KG1fh9Of6Vpra9Zvx7GxC3ryge4tku/9i4gaIU
QKh0XJgXsF5G4dNFEXOEJQkxq7tnjgNW4cDSDvKV3Y6IEqmGeVQiPKK7/H7mVcy3
AW41+Q/VDzOCwiXKSuSXbLV3RRh1eDYkggfZmBMnd5TbSXQ3Zbqh1LpEbdIh23jG
qZ9gA2ZapaE83bEmFOioHhE5gqKS4czmwcm2z6BEvQ/wjdvQZUyVImkheaB509GD
LNB/PZtJ+hh1XxTdsLlp3lMZGX4+B4RbOpIVvbwkgx5kJeSBfYsaWgGDgRTBMHQB
kSWdl5F8/2pE9168DNY6P9hTdO4epZ8yCAxgWjYmm41cS95oIZBi8bSa6A9gDQhc
TlomiGf4XHovPLsUX33eGUvahZJPf4SNpk7WnLoZa2+pxaqYNVAzbg4EsDiWQBjN
uPFqhlLCcBJa/p/ER2yXCbOO0CN5EDb6ANavEcK5tXhdvtOGYfSt71be8NG0/P1i
nyjdOo9OyOvPvR8mp35IBDK+7YOA/62/NRPJx+yf6EmOA6IL/fs8FbreY1uoXyZ/
CMa5Vb3jMm2hzI4sljFDLrrHtEFtcHrKmQGncL9HUKp6eUjs/hijNtaFs1SnKSfK
R7RTwqFAietrN2tsynoybF2h++czNoeBSnsRLFefu9+k17OCs7ZnTR8aZioLEWoB
lEP86mIOOklsMT3zZ8+1t0eLcEKvb/3ejw7LAVTWX2DIUIsCynO47ig2IlXEuEXK
IfTWCKzzuB0kQg2e/PfMaPSnPVlAotU0A72U0fBn0gUMxwTMp5nOZOn2QcMQYJHj
6QBBiGorZL1Sakb0kvn4Wg8PvKuwGLbYZ4L+UcOvDQ+1qwuUkArAqE6JgG0c774q
6k9A1n0kCdZeCB8jDY0hfuY8IKuoHIINd+6+HXNSFM3OIln91V9I19tD1M8eRsOL
CSB0m0rZ3hEATNESyuV1qi5rm0cbaufWIKtL5fxPcsVGzoBunKhKif6RLnAN1cMm
JbrccDck9/De5+cmdE5qSkHt3UsPgN/lUnzbyX5+IycTBCiiig0bGYpPZU19kCK9
5wGdkMlIuMdrlhmk+FfZxOVop89OGmr1ewvFDz43fBDP36PKD+gbCDFfAJTSr5sR
Sl2l4SRF9EwW8UzCf62lhxO/fsi8weoFBsd160aS2MMxAF9n1sU0Xjz9bc6CEylM
ceg+FWRdKQAcB9mCpY86gjFs3fLdnyELzxjN3/L+poTpuh62k/GMobny3C9lHdtD
kMwNSLcVymsqlugAA5YK+GTIjYIwev/9LNFfQSiNpYM/hPNqPmSikFKGSks8spJm
q5K6Foh6UCmLm5DBOWvKOWe0M+BbBeZojjqEn7xn40YheZm5N3iyWhUof/o3wnDz
4G+HwdQS+L2Yhkijn7YokuQyvVfGdAP0oWeVl3rVCywsXEkmp1BFEwQdO9fXA5Il
0nYcPleom7qORbIwGqx6H1wTB17N4gigEj/OURWRj5dvRTbGWOxakvqEXbJeOvhq
p5javQJrPUQ1NW/shf3YQZTEe+zhnaxJyMpd44Dcd5LlyhsP9uYHQKgrrL7JNTJr
rmHMjLONfdtx8kVsEef/CN2t4KP9JePGyz9/77HoaiutU7OVHd30cW7cctBuuwON
9C8CexlkD1Sd8TNuZWwZyTl2CK9XeBGqluJwkNjq9bXMR0nV80iUq3pdeIASRnnH
8fa7yrgTNhgRflgb0LdZvjZHp6rwzJuaMm1CgzmTXMrtJHl+omkUTVMnYywnWBkG
lxnXyqnGUBdB6Z5IAn8IFcRCvfRwUTZ1PN50e8h+jIiXSlOtfnDVA0KJW4jfkRyk
10OxdeVpfUhwg4jSmQE+yTquhG6gEy/pqU6pBGxd42vTPwhyd0+ORqZ8dCDbgdou
ORNxbGNY903iUtU50eNI/ONWiBq0YcdeDuGjyKecrsQJfGUEc6pP9CSUc/sYAiZk
XN/ScJC3XwDSM1YpjEscnLjEu4Bc5osb+EmTFmIUJa7sE0ju9Maf5FWqoC7K6M5I
HVsNBuc69CiyJBTNVKH1otZjZl+0eCs7ZlmmMT5NHTrg9aOkjdXM3Q6lC2MRlbZz
h/rNxT9FIh94NE5J1tyDJSHUAg3afgkg8RHD9BHI2ta9XWoB1RKrAMfVuHh37OBG
gmK+EJQSGvw+Fm3O+ti9mrRu0CBtTy1Ps9weszQcfjrJjyavFi1SbnPUr+Ku7N4X
EII20PgQl09kRqhb+w2pBmqdRJD9FxPI6cLNlhBOYCJuPNi9Zp+ajh6jsNxbX1E+
DkXv8gcbewcid8vMu7W8DwKN1w14vC55ksdpmbPeb4L4lMZbJehcDHBGsJJCxVKT
Gou9Kc4FHwB0Qs4z6lf/60S7DgB4wV4URBwPIP1IbNfUKSvgA6m8VsTlFGa/BAkU
EQ4eWE+UwdGltwE1ah1J5wWSNaaFhI1XBZAnFAV0zIc7IzwdX4iDJs1ff6PnIN89
PbCWGtaIztP3b/rd5rOY610YDxeUVN47pwTKQ26JUaKEniCCZnjhjg8OWy7QXwrF
80u3IBf++U5p9qe6vLFfgattod96t3xoMHTNQgRctZ1CZ7rMCroPHxoi5BF3dk56
RaLlROTqkVJZ+zm6/DbB4pZSjH1SWLX8ZduJOCwv2YG4erHNOA8FLyu4rgg1tAQw
yshwTFdHlBDHq2LKmpJwJN+L9KeUK/NKWEJA1MHyhDPco69OQ9dSxyc78MOFIfz4
K/BbmQGJ15Y922jGm0KKdlN88dNfD6+oq4DvaIxO6w8nOrPOY2OMX2iqK2NmmDeY
5LBLBvPp7w3P+iRfAH8d7pwOFTJwmqjSP8JCTSQdmLLUfGaqXfHJ0YY1oxQQ+YXk
mXHhhOw0Vh4ExM24cTpeotF+dNhYj39VEXjdXyQVmgNfBC9l2KvIejT29/4Qc3t9
aWFTdVu0AmG4PWqBUFCyMeekuZVOQFVKJYfbIOu2cP+j7Uh2F2OQN20m2n+r80hP
KYEt41VV33HJMl2CGYghCArbPqmXx5kI34L3LihSNb6SZ1IIkAg7o7QlW9KmtZRC
2l8To2MWgTuXUGNMcP9n/5qh98wnGrA+9x7QgFgxgZzp9m8THRUT7C4KxCuhmcsx
8vKl2i84vrj2AzTon0QBcacZPAoNoEi6DgE9Jb4b2Sb0kwh/wJ6SuWt936KvzfLN
GNipBlRwVIx2exg8pp38E35rNIJRdCObwyMDyD2SbMvkfxSQRQ4uZvfEj4CXN+um
wlDQC+mSmvikMqcpYBxnzK76Qhqg0XSc4dGRbysC/22KIhw1c8ZuY1tUx3qL6TC6
MB3fMkWdssaGxG2KSPLNr4dO0X1z0KEtKXImkEoOzIWN73uEQbmkWgHCzB1fFRA6
kYykLvgflbMN6SE8gk5sGe5WKa28S5yA5kI5863DFmfUqMpJsZKMX95WiSG6Bm19
K5ZwCku1Q0GHB+iTES1tVum+eRyN5goTHMkTke3BoKgruPaDCUWEha6sxrFhaBB1
A9dTZ9K9pnFzBQyfF/HSB/SI97hxaP0IwbsuFFv1QjRLd02iybNaJdCAqby12KlD
HCRotGYDIdb5OwnbVKXZjUBVd2l7CPGrvEYPEpNP9gyXTm445BwfBEtW3tZE95GA
S1c3aa45CzX8XY/bRqJEgsqytjXpQeIfgDKxa/DAp+EEEoCYvyUvEkI874yHThuD
41/t5X9AV3S3W7oHR59xaOM/sWccBCzS6pDv8B4pkg/ao4NvVkALDbfzgwzzGKey
X5nQZWdj1n83OdbqFNQm9966uGLDWLG9BdWWXHBh4c4B7EvgyjPYQhC0fKhnDSjQ
rCYNfPv0x/l+EklI71Lvk2UupthCKJdZepaoTst2DObUdB2M/hhh5eRXQ/i7g5XR
ohGrUZpWBmm/Qw+kwVXInZqiJxgaTiUkMHlf0c0lszgPDb9lfYCrMl0IlPHNKajW
c+otCoLl6o5jU7o5JkGjwYBtVdNSLlpslFwVCZrZGiUxgxg0khbWsDrNLpyztjjZ
DwUiFaxjetGTdO0Q/0VjtfbY8tnrADVNYBJeHhg+kY1ljaVpeo3HAqpIZrRLbNhW
Kvw2dABiCSvXGmXRYpABRg0DySa4a5EGlwnD7G9vNgNE40U1piBqvgm/qzpImu+y
sdQjUqOuGDjhepZpfNL/y5vB5A8TPyMw1IER148k5Xq9qfR4D3+UuHrgPgKx7MCS
fp8l3JUDa3fcrHJw4KWWUQUMwUychVjhakl1yCIryttRtaCoPkCygvBk0cCdas9E
lg8k5SG+/V8x/tXH0XNjGjK0s9kw+1qyPI720tjeep3NR/hfingPSshfRaegAeE9
3mY5qDKccX0McbaKm5xrZmyxMjEaZICXbk1hDZ+MUARDlkNUcdE1drh0bxG0LtJv
sISMm8GqUoeong/zabnCc6mMT4WKxvGUrJ46zAP18GmXOC5wy3x8nWuhq5V0ussG
lilNyK3fY+DH5FaGGGBmlnNRiSJUXorJYH8V21rX5UPXbbvWxMXEJsP6tnBySgll
2Cz7cfZJ4ybyxnt1GsEdugVa3kFdYivdG5kQsJXHOdbPdVDue3DeplZAz72CGpV/
Cnb558VkNvSztzIPl6LVAL1o1GqH+uEsaik9w/js8kwfEkG/hyfcHl9GXuvgo9cD
dTV+ziuaf/UKUTaJzDyx00SljTUBA3iuoXJDeluVCMX2wIb0sRXnqLTxZOvLHS29
1Vd7WwFuUPhh2VblylnFcw4q0vrKRGQn0gqmkDNb77L+6vWSibVY6YP0ZzTubfGZ
t30lgXmg0OtxDfmDOJ56lfGMwM73UXS1o1uawtPKbPsuvvHJ1AeNFpYhNbS+z1Pt
/udZ79pKm7ez48tGjA8UO0dVty8aZMwdw1k9+7J5Yl/Ilhl8qK497fKBUq5/EPGe
tSvE7SrzDlGvJIAhb5ZIyrdtUPusQXsgqjZOmt5lcp6NGwjhT84yP4Rk4aubFpHA
vmPlOs1KJMI44BaRKFLWA2/653KfrKRv5eoxFgLPA65Kmu+PphpZpO/ERV2lgeXT
tRO/XwRTbpHcsF8mH7UUQYQPGw93eSMI8WJf6FvJpSd3/0/MxyYqmx+iO43wm3Bc
tFhf2EIcrDmo3D9kzAFoBmtdxQfQ9G/sgOfzf/SWw8UcAtHQjE4D4kB/36DSWKUh
MjbkjSl7GLir5MCwfvpKQmNKXGjMCh+yjIPN2c7cqsfeYgvWWiMbO7aa+lVpy77C
HGI1K+NJv87HyyFzMTJw/Jxr3FfVEWMtTanrQUPaPzBnff2QdJy1O/X/j9GKJu4O
mhwq5oHa9nUrG60UeXTZ7rU5qK+Zc3/CrlLrGFpSX3TYxYFv5+kCH7KTK4hZgsd5
cb8Ju/5U85kRMY7v8hlcBGO17+zxtBiF1l4K7VYCykIFO43rIeO8CudKr4q6zfoe
8FvIbj+LiT68D3cRLj3+t+qF5M5ipVWA47tqtZs6dzof4/fL3xqmiGvxFjzcHZDO
mKa6pL9ftSu5rIiYJfkrkwYXIihp3pv9A952X5+I3qCOy/XiDcaupaX0g6VMnztR
OsitNFqli85dy4iVHZ+C5WfmWWpAmCVxZHy4YY8LBtIWSBhaiIA88pbLA9SvZafI
Y29bOGcyE1CCWijGqxVYHscCfVTGzEOS8F11nMXJIrxsY+cAjK1P8tNB7jeUzSq+
YoA+CBKW3OquE/tNH4CdXhACyylHKUOxxr6E5qYgwZspC+s8gMSqyYW6GBBe/YzC
72IZHqEhj5Qczm7ZFoAC3/QzJUoZXVxZOuzQ7dlJUDZsSRs7MOUbIHA6PiAt6+Jv
UvlvcVI4cJr6Ebu2IDec0dPNPS4LpFK/s8hSbSkhKQkxn5qgzkXdZDgUKWByHnyn
iaz9oMb2ntx4cuIeKymGgAu6l37BhmoTpQToKdBTAnIZ/KNsWcnVLrk8oyXz0dTT
a4LkSbmKZVMPEF600j7uQwr+V89TDXSSEBG9t6wdcDfO4CdJ3/MWn/Pfk5eu8lo9
Xok9/EmYGuR8MzqG07UOLjeBkK3JM/zv1ERiPuhm5q/gOpkO7Fx5mX9PSJnZgQuR
G94eyYfaiMPRtAwCtABvR5yHF6sIK1j+EXb8qj+FelpHTZ6r8mYP0XVtLoyFyrTL
EsuPozExmr47mz47QRqflCcczRaH7/33/y2WePrXxqjT9tyQeoV6Mp26sRAO0WVi
IfL0tCIn3ywCkJmlY5CADWVnC6PCOaSBPaIjYpvYwib7LK83BHTNvCnZvnFewt5Y
AgmTdjlWkeT4+Dv9Wcxf3IBfB+w3wBw66cdc23rk1GDd2jaGG+780tvkMu3mr0NL
Zaa30kyXieKSMuQWKxevivR0jvL7vYJwqKMg8I92L8BraO8GNs6X5snjtFo3FakR
TNUvw7cEYwAwfw+Sphl3wGyQ0JQj3VPebLTzD6aLZOri2VYtPUx4KcpLx08o9PBG
f1Sx/1rJOXlM281NIDcV6dH3HSIOWE6rr8IuMWodNpLG0JvY6DlmCvNXGBSTZokE
id0DTkddP+uDcBx6VRNtL2qyGNIqjlrXNiBjPqSAMGJ1fbUHGiyt2SogOehVtXrb
sdQT+w2iVYlS0fyfLxHWbHfKabdY2pCGKQhBdqU9H2cBtu1EBttB+LOVF5rirP+5
2JgZ871NAiyJPrtOYLQsg+ZsXYzAW1U9DxBweQj4ts4dMTPIINK42wmxZfYabQgg
roZ+xZfuzUmmFjVUvMit+0FiTk82FhfSWyL2bS+gfk/i5RiysSk61fo2yLm2nYAx
4gnirL0Wo+s25g2aHVCu46MfXRSmhCMFs3x1rybAklp5ZGJSRqFwWxHz/DH0hS0M
X+NWIuRjOImqaes5nfhQFo/3MeSg+xDBjuSoRQ1SDE5CiTdmFiy7x+8xM2WinV8s
VKGviZwDgW+VJqvmx13CWTUxvmRmEVBx0CbQvCM7PXaeUOPd/BEWDws0FS/Ne7fu
HSBUdZEd59IgeEHPqzof5rH2kKYKaocGzjD4LafjYzpLQyEK70af6frb/EbtYUkW
NC6lVo9ETtYVzlzunfVzZ+5mnkMecN1P3KMVogiW1BngFUYwtJyHmXbbMA2hAC/5
b+8McQ+D7uU66v1k8B/UF8JzNh4HZsqHgsBOzetCAOtlKBt/cWIGZbzvLUus+zFl
CvIuMbjZOQkslpb/4ci6qjVzrr7L4fUTPxcXaKvgSuyN72dsEQ2uYqPmcfoc+py2
b6Xw2risCIJvO8j755plZhnLw8FNmkmA9sXy8IOrTfJqkCdOhuZKlX/JXs9beSan
xw8904mfzM2Rr3uUa9sCARLDd3RWkxnP7d7Se9Y87vilDzfuH9shFFPrwzkzpKpT
QKKoogAxaeJbWqnxWaulEH8aCb8+0NYjDibvgmD+rE9zQkyax+sqtCA2trPgbx3q
HI/K+4ySwvOjaZj5QEk4GvbthIDJZEheeYg1O3sDUaWLI22S94NBNhkhovCVIhi8
vSlSXdi9O100KACe1KLfLgDBsOaRscCi3hoCWVAjPAwyB56VXs+SzZ8RNCN41FaF
XDA0dadByzyHWnn4cJJzDnMCDXlXV0HrwwSEv4kk/EuQdfbzCle8K7fmZA9++Fvy
dTHl1G25ij/b9PEsE4aePLbdW7QAiACslI0db7bo2B4IynWTr2tRK3d9nG7acmzP
UC1dOGueAzrBulbsqI9P6lCrQ5fsuVtmJPb9h1g8cxh70HYZfLqFAvh7rKb+nFIi
wcXaa5hm1a/Jct74IeBik0bDQtqLBp80G+s2j/87IFAsxGsPrdHEdCXiw+fO5Lly
Hg5uOoA9aAbvVQbQ9fzMoCbTVZ7fLZqficem0trEyEvnNHtfEbuyOj8F8a9eD8p4
/C7UTh7ilrFEsUKi8PR7kEuwDx/gnCdVP0x8Tr/Yb1uou1S7ByXZxDvc/WFszgQG
fMNIHCZz00+ZgSh4CDM+ZtAKA0DfsVjpGODCa/4qF3CHHqPtjPg4iJXMUntZAuYS
Mi0oq3FjSvx90duG6ZeuxcBGB2yX1PIWxZaYMNMc6n02xGrOG5zYHWtTtK1RYW1h
WQKc6iHke7qH1GsoL6ugR08n1UtmT55LRRhepYoguEIb+bb86DpuIEsyFyKYSVTJ
C7xq8r4hbL1orfLBiy8oYaSEqmlZ6HhKl2MkpOY5ZjVi/eJ+IFUTiT0CoChRxpoy
NT0I7SNwSbAQrIsg0BxII5+QD96mF5gq9hs6nOSxq+KyKL+mHP06IyXmWjaP48Sm
oWOGdm/wCkROCURwJQcRlJwgOUtvYygyWWZRRy4riZ3NTmh+CWimt9aTPUgrBkM7
OAErDjQmzPCEFYDKlt26Tuy1DnbegXzqLXvOZvhzmrRnOT/XdNfxSzFD1Nb1BWSF
jvpnL92arhk1nCrEwjPDzNTdn5NzhNgvpuZw/yzL7Gpr/zTjVGC6cPVUu0EAPXrW
hXeR1gVc1F4ezmw0ZY2lXTpn3feHdV3WQSDzVsBxuCZiYvt4Cv7XlxUhjkGR1h77
qGZKicwxv4bn+hJNRWEJ5q0B2eIcbsCPYATRogY00QsYHPsnwglP9/TQbk0yDNYM
qvQk3ZKCZ28h/ztvUlMW1C5ezOSnRbCJI4Vg7dwoM4Up5g/8U42ZL+Gx4QBy8T/z
hsunfWw7c3Up1ZhGgR0Ipby8AZQxN6RCtPQvpGgcmdh+3F/uKIXM1FdVL/5Hj9nn
GtSKK07nZ0VGnMxSzjTh6QuXF6WXSqE1fY1dB0jvkbWzKzVQrUYutaMOmECzZ1Ar
p8P9L4XPmNpuFUqfZo9IE3/RLzuTgTjJCpuEQp3DaAsTcXgghNF7DkolfZL+6hws
5utCJLMixlqTpJg9ml0Nkob1RncWDINdrA8V5fmE1CRDNtVhwtl1PfEG8MpfMq2A
E6vzCD19h/mnk0WD2932UclCMNNEnr9nAUKvCIf3Lx5wzuuqYiNQ8UGGVmjKu1Tn
/usSBXoqegyni/US1SanC/5TsIJU20xirLkT/mm9aVvAQ03gAr6aaoULGtqND+IW
/BqSS+C9TJFkqHv+b4bouykCLzaZKN98i8nvFY7rdtGE/czJvjzA5u+2QwSfjmPe
Yj4K6PagJewpSTcd9mVQ9mtNCADRH9RlRr9Tktpvn+k6zJER9OU4NNMapH9CaPdh
DIqoSeX3P2fCw21wtxOssDHfIQPWunbEw/xgDjGY2C2Ka70R2pWk6HXdTk91TRSn
p1I0YIancCte3QzqaolLXaZ7l7zfZOf54YQza9HKadyDuZS6H2XNO6xmbbUj5fnI
bxaEVk5R0B57IYDuKCwGpGzepVLdzzaM+Dz+bO6EBnFPAfDVj63MKvdz5C4zq7UB
oOxyRiPp2zwPaiqZXWIdohwMSvu/UAcGMmrflLEDzVd102JVIfhYDfoFqkP74oTC
XhLkf+mpUttgVyqmR0XaRrfdYhggWbrElGK/ZfChGz2CgAy/e/eCG4sa79A0JQdt
wK6N36n45+ZoUYUEjSwgNOV+L7V1tASpLm9oFdE/miDccPczUvkl3Qh2ZQxSnU4Z
qwHBEzr2lyr11ZFgF9rvAQ4SDxsrUIBO/bcwUFM9VUyeCVsBjSR+ib/09kkFiuQ8
l9cjSC7RKi8gsuOQfKhYd1NI1654zSVU/kyV6kctIdxd57FtMiUgRdfp4bOL6mbx
aJ/UfPWtvZGZcKqwsM0o9sJsRlqGULJxVTrGIoto4GV8TXv1oyBCnRMbdyiNtqRY
Ofr1bQBidHsaZOsALkgaPHUuNkuDpPMcRa9Q4OnhokqHbbWEQnTSJrmasBE2+sH7
HbKMh/R/tlA5KuYYW1dZDappZtE5OqbkP+C9Rv9nW0p1BRk7CRYM+Jd/1dd/iYYG
bJbqrgkpuvy3G4gLwe6NMak6Ms763mz/tY0yZfd7AtHK7ko+09iAjGLz8VlQgTfr
iFpi2+853RtJugqC7VnIJZpXhGTJZ+FJtAyOaqyn9HkKsLBYw5j4qkXTgPerc8qB
eVKk1KQOJ9IQbCNSvquQlnWwRf6a0y8/QDqNKbVzEz5MchMjWY9PGJ5wmtms4aYk
huf67YVCJ/ISvdtCgWu6g9kzumikXSjlDwzvmL22odmEm+DiUk7cHusX9GUWlJiD
DFoOz8jvC2k72goY4Caf0nopdVqz3f9ZgmloX0ccuzFitxrdXEieT8JJdYCMEIwB
m8hjdGW2kzNaCH56ckYJEUYc8UsT6ueytnIBLV70+lEzU2f2tYmfUB2l5mpB7P3X
XWafXfteUydZl+taCtnC5BuwvvTnH+vZTKhjkI5/+jvbMhUTHBmMAzrjfA8ov4ul
0QXmSMpV9ZStfBcEjZ5CxSlXlUlleH6rD3cJz7VwR2twCheuzmxhNRjSudlIrQia
ggB+s0cEBERRw89L2yyfw0RuSYq1/5v4Rcd+3RsQyQZU0dhew8iDaYl+4I4/USk9
OX5uuM7w+0SP6lL+4mwXWAg2K9hzRP4OagBBKs8UvuruBuCzVPb0GxfnZFk/TGEZ
Oq+xe/YpcwrQi9iKVvo5/JeiFAVl7Zalmr1xidzqrAuCsT0RcpjRHHk9Bi43rj1P
ntUK6xLwUaaNGKAs7KYVvszHDO9cY7mly0EUHlUxWShyYWuNoxLQFiLiiypmBIrm
/MFrRtp/9Ky3AbEN5NLbhgWtYldS5n+UO4eZuqoC/jIkxXg8x7w3GosiECXSpFYG
RjCTi7lvj5hfLs23zhCQHmGvWF+xfHXmNQk12GL4fT2OuYxOwDivuaV5/V9lTRZc
40d4NCEWEBvViQfdJsFiEr2lVfK/IHC3ryPCr9Rn4AmPKhRjDjhP70ysw5qFj/3p
uq7WvLY8ex5QOZuTADygXzhOL0nSypJNMnaADNe+oLmtmKU23SMJOuDlflujOphY
o8KJh3uMlOuNkDBrQvOVVlmo8KQkQXbmE9LMR50OFFio+7bzhsUGRiV0nyLfohMp
Ur6BrmijM3FDzi9PxKCovg/dl2ldHa6x2ao3LMtGyjVlTO1tiFu25OAHmNrwcxBP
PxrMgO2Ya5wLFhTB/szf8ZkEIhfFD7MdGDcax/Sup4dy2dchdVjU5jJHdjQc8uIC
drcKztOSRmnwQBXrqDMEWrqobMMVuq7ttBCT37d+sjFScKPyPUaFAeckAUTBccnj
4KX8gKZGw29sVF1gCqHrV5LYXRjzL1jJxYHYOCLgBxdjmtYvRabBxV2Bk4PJSA4n
8TDWo7f6JTI+ZIPa+KMR+fssuGmCWGzTqlFIvKgPIoxZN9+9mF1IBpmI7n4G3qt2
93Jn8R56IFFui2oG21m5b503DfH/p4DNEZ3AAS1ZDbAmxrK7v6kUosbkYbn4OXlq
E6cuy+SO3X5znNvGQtZVRtoYRBT4g7O9vcaA6a2v2E+rO7OK0esnRzHkWVMhUGH2
PsaV2lS3BODTCr1f/UOKoEAsVnWeq8C6vv61Q9ObyaUVrh7GJClumT/+Ckr4sIgJ
9LXn24tHID6s7Lo+H2DDiSJSBSS3QaFWhk4i00/zaLVTn5hE+GrbIF2zqhlI1jWh
3ButpvqWpr4r6uSe3yVaIb4MvNYCeKUncWrtGeexPRkCf1/jmgNaSedLX1KomgIF
ttu8TNE91wWUXrVDPpqoEX3n8VZ8EnZQ9Y64wmuCnyaHkR8fB2meWq61B9/2zrrg
Ctlj3AmOnDe6qf2f2rC85W8ILFRKT5fD0qlK30muUwLvd1Yh101qlAopX+IbRtfL
C3ofGx4s2APTjkX/tbsMq13uL2zwA1kCpmAEYw+SkhHJmCAV8cTryxNiDMB1xkqR
838lpKAIZc0CCCJBerwyDdUKaB2WM5bsjjtoZ/fBd418p3O/06Pnch3gnJNTouFs
LaS1EnHGqLL86fJmkMCBgZgc/p7TJYvUp20vGmLP2isSKuxHvjcJhIjT7Bpo6hKv
odBCF7wbOEZ30czEPUFYfHFv5AQ3osvHlAF7X/rTmwFS5wknzS7fry7kb1i7Va35
JnZoWsZGeCKcKKWJD7mLAbcE+F859l65gV1Jz/8zhpsZTs1rGqn9z9H6uqUmZCQJ
UXksqVhaEM/98bx3++yAlXg7keQNNmpIwRYsEFveitXhxkBqnDZZwBIToJWsvNXw
t8gU56XJSwy1xcvOVixUPFrVzzs1HaZOK6vAP+dxK1441TwdSAaOlnxbu3LC/bYK
HU3Pv2Wv59taTnV1/hIhDTLZF0YOe+k2BeR9xr4FqO6Om1jOZsL0JYgjakaUF847
PgfYxm88BCnky7WNtwWzsYOB7WiVWb9uT+UX4QIciGsSQIS+RrM32UwmtQry7rh7
FttYnzD2/fU2AuSP/gKLGoDucqpKGNFVMLQIwmYBdYwpaGh6UJFzdbZGJunpdMqP
7znvzBLrLopJOFWBUkxdENC/w7N0u9OFYMKvSpU/nzXA4+VrPGi7tHfrUGQNd+9G
2sWVr3IacHz4Vd5veBqwjfmjKxJmTNIVmT/yYpqY+bbIfdIXY7JxC4u+hk9uVg91
ae4Th7qIYM6RSwH8ur/uW2X2xaGGWq4iDeZQQ9l9UUebmW06seQVrMJ/z/Gkm/P1
dulagg8MrC3Nld6RkPIqWpdaYBm9RDWZAZYJ4sLcNkpauJxpCYxGuKrz85sXuRH+
rKWSLQJZ4zjWv/DC3AICrYBbN9rPnwwRfXE/0/MHMH4ZGKzk3oDID5UVsLYzHdOh
0OYpoaoLx4716NFV1bp6EzBTwWnRu8KA+TOFIGxM4i8lQZaEghwT17ydUFksOIIs
QNujrE9VCbnDFsSA81qn2wup6pVcDVf0JeFCoVlsB/ImxbPZTEO9kyy2uNCnUiLL
jL4c6wJVnZFm83yz1ZNZrQwwqVlx2it3XTpVp7PrLyG/6SDLTMFdjcNohCMtFIIQ
o4s8MVL20odQAqfld8n+gqCftG6/qt/wJpbMLb3KF7QoLkRuvBw/05LEeHdx961J
bbUjUlJqV5GN8PCKhb5RZZpeL7szM/Iw1dVGyXRUhW9gCwOmIKLM18BqKW+vtPBS
6+gk/x/4s8FePYyt0JToUTEDfZgzmM/5OfOpzYrv7FxgEVIUHVkxqvNuo8YXnRfw
9rxoPfP3lpuqEQHTl459PGRJcX5QY57yF1ACrk+rHMAZZ+i0LnB9m8+NiaQjqzPH
G4uIA9QDF+e8N+z85pgoBdEFwlsfFd3+YFUcTg/03dYeAn1E65WmXFfJCO12qF8Z
KjjcvdvmmxMAW+jSme8SZntNAyGYxSVG3xpI/Y1lrtNiLX7wtHcF9POVAOAt4L4H
NJPbuU5tw/PGgqdtV/q18FoT9E000FrpZYRd/lYh3fAjZ52WrGCbNGz5SxLBQBQY
SUKz+DXdhcDNMXF0FFihri+OYnhUeZktCDJ8qMz5O2nvbJXQHSsIZFrgvxriFhYI
VEX4M4M11AKCli88fL88WVP8BfynulW7/JxQGysV4bLqtRv+hYE//hv3YblCG9P2
gHfGSluJ0LTVGJBCBpXFZzPHZnxQNrnl7W0thooeVkGcvot3rzmxKpQ8VYJdTzT9
s9dcy/VzSZaGE8v6/onr5B5PYDhtp3ly8WUK5HAPDDlpQ1t6F/5cDxpXlbcgdMcY
Dcn2qOKWVPhkU2Ujmk1/0vME8B+fkQa+gjiNv9yHryNxqKMsgfiYieeACVPh2Gn4
Ut0u2Iyfct8pE2LRz27LplF//ja1PKFKNvil+BP3LB3dptzo6IeQDkhCgzZhtz74
rLRWm2tUei81/fet3CkKwlBcUOBGi5FfFUBY7V3hRv4bWrJz9QTQDrcAyP3JpV8+
IEQg5MrLK4kDBC9RM7z/ZX4VqRdTeRu8ZJ/KXspu6+h3UYXa3d7BL1UAXH5UUyDb
iQAK4vn7Y+qU0jDLPUyDo1bc4ukQaV3X/gHHJjgZbIvdCAS+dnw3aZO2/OBYPVjb
FgzRUmk1h87S/XL4kgiKdKGoZB6iYpUsQdW58RtC600thdpVJYqBHhTkG0wWA/i7
Wr2/yb8qZR2wpM+K4DyccsMl1/o0ByPyvoMCADqri4XBPmfFQjI6PDFFL1hJ14Vj
MMCJD1n/4cZ6tRywN5FCjGiHAy5AQQMXm879G7HTjYdUwc+Fz88YeA5y6tRio/9s
vkojiPqJXGA4+ikHL0uzz3Z1rUWRJEBVOcf1X/eEZjJAw5xV2cKGA+9I823gAIZ/
82GxOJhTL6bq/FxaUY+/Wr9dAicnFsFqsn4Eh2d0vlD6c+7dPutbCowCT5ocjJ/m
rJ/3Kt+dGXZZCllxXYjppHIS0M+8RMYMDnI9BEyFQ5t1vEh7ddAgllqThbVm62d/
5MNTSzf+R/2gzy9caNcjp+Ki1SXhCE6aoeKAJ+/vJitREE3Oanzo8TdorYWZO4i/
GTRUrIY1BZOKvWx8maqbiv9bsuwqcdlioCb7CY3UgYK9QPAilKthW6pT3Bz5qXFz
lmZPiVOs/AFPK2mZWxa/9BMzKRPr5paA9lUMedPE58mGNiw3mwC2rTRSDknOJAYa
iCf4K5Nixw8G7IudGNcg+GabbshyJH6NRf5tq3o82gni34imhFFf4LgXwP6v+hlr
s1sKKVuLaDXFg+WlTuLLgSzwG5p+BSGrgEvtUmV+szC62/O6uFxGs/CUufUlltH0
oi/KplYkVItKMBBpmQMXpZAoqHfbiRA6/1uSldP2zuY6pMt7zJGBjyIlH/myEHcl
mLnKSOvEs8Q+4En+napNUUzTCMfRpe/rvSkFkN5pDp1/F65GNbXr10cYSJzerQo9
3GSa0QPOR6ydaBblWXVeFoJ3Xxs4VYKfsKzgNa9uDAOp7zLKv5FAZBkskjhP1lYt
17Jr3TYUjplqweM85LoqhdiiUm/8mB080a5WtvEbCcPP2TkmF+ROrdqWRRVokfng
DO+/F7ClWkTrNvCSXuL00MQUAvVd5C9c7zcXAgkRekVk3NhknkvnfJUL7Dlinx+H
8W1RQO6hTV4o/45fCxt9xqALNFjNJtQzrq3L2ROKXa5OBk5BEDQpCh6t1V44VJrL
qvfNK8GZSz1ovpNGBqtL2HJNzqfKhQj3sggCrX//Cyu6lmrJgvR9iN/mCagZIs2I
e9YbUANN/A3bJjeou0I7WY9nzWaXNpcJWCQ6FWhyV02L+Pdn+JVzkwoyVXslwP9K
PGlSQdM2TUIl6SywPewWLWKIPaQUimosAVLd5HXmwBCDNCRCB2xaFgiaa9S3NnjD
WcNOTFDO48EXq2pE6LUSzwiW6wMifJOVf5rejKNtUFwM6PlB5qp4nAElSiYOa84h
V0kDDEr7NZDFqrmIoGI7AoIyGKNtx79lFqg7FGxrNNt4TIxrsvyhWcjcDBo07hO3
rlXpBsDDiGD1M6ralQU9hU+PL4a+tf0z2hnYnc9pCMBo1hfGyV8xMmz8Zd45vGtH
8/p2hlFw60TTOptOutwZ7uTDAND/ANSWMXNXNG6zRQwzCFMgS750a8CdjwDDaBsV
oMFUtuSdvlcrdTuraNUtcTPvBBjQIGcYGa6W3sCsURo3AGZQfflryWiawRuqz+Ww
oUwT88avSaaHABB1lUZwyKKuIyvYaHbAJaZ0zRsMGZPBgWlEU0QtBsYn4PVuYbkR
xfNlpbl71slvEEFjNC0mk+x3LWk7UZgS6E/XUUTvYJIEP4BLStEL4Q/VtF5H7iNU
2T/TnadP6TW+39INszb3WYI3D38NAUZFuKbRqR2ksMLwzmOzbBoFGv/Yiso4TQ3d
8H/SICvEb6oL052JoOV7bMhMIIjKxODA4ynGMoLdXeEFtEWXsk1HhECnl/Ir0Jml
zqFjxCX5rjuNNtaTEn9FZjBBfv0iZ3rl7MSLspX/yM9uPCy49quvmajtdFYU6MVj
cmAGAhxrq1UazLdOfdl3X8q2ziUhVJCsBXSKk5PxSt+bYSyuDVxQ4qZKGXN6dzzo
KYmsHiT9aC6LI65c1zep+Udm7No/wyicTcRwosf/hl7zkXAXrAVgmVczCQ714zgJ
tVdDa5N0wmVmC6g18jhg2jajzRs4R9eb38jQQGlRnEy9Iv3oMmkRhEEcDBRc/mch
TP4WMUyQOfwUK7AlQgSzsR/TBlu/TXEo3nigYi3c0bvewGRmvJJsz7yG6adcHFvt
omNJJYjxgtDVJ6te6kboybyQsEB/BGOKBDywQm/B9jkA9kHFvAgSVsn4fYpBZgQZ
sqzGltJ40rZKAhgpH3+uAr0uqnmPl0LXAZX2NNhl3/aJ4BNlvQDYOFA2HG4lxaeW
aWl+1mQlRgQJDm5ehbV0spIa7qkg45uMRbE4DcIxTHVN6loevJ/8b7D1HcgYCd2I
cRkHf0uIJDpXixlDp1lvuNYBLTLcpopnVTFZJYOmhrltXxbfSZBt4vlSEQj7q8du
ry3ROGXxrYz1gak+bXzcdTC4g4I1CqgrOFdJB70HiU+zX1DWkcN0nYFn6q088vc4
ZxAGxGj1s04JHUI+2GadZ4rYfcxYdWE66DFXHlT+ZlKt61ydYLpvNt+07/ytb6Pw
3YityU5mTomZmofEbM3UjRTGTS6MjZXsfB9/U247fmf6jyxa+2uZZul62Wlwl5Ar
nDK+KxJyRyTxWq3n+83hIeJUOb3NE6y5K24XINZfIVobD+x6683DPaSJIFIsWIHf
/P6Cyd/yv9/spjQ5KRJLXkpiy+fYwlQWCXx1J3Ihntx5/JLuhAlkl4ZQxUOEl8GU
sNw10LGM/qrC95KP0oK+2IPbMATH2yrzeYUTKlov3LO4MNZxZpCrwcvtAZ1kJNCg
K8Mjppv549JcCCijgCxxWGO3k+GaD/QYoaPl5T7FYBg9uJAh5NOaG+WEmgqOmEVp
C08IKptpen2Zhxmck4Pi5rxrdrZ6ZAJRwvwik6IZAQqzuK8hAn9riwkXFEedtpaz
+TFe23498tRxfnJ/DKrhPwxFNvurdKod8Ue9bQ2HSc0WU+QkyhPqFl7E7Ef07XOP
vfWVbX4pNbYaK5iLGifqYoyzYvj6ToZvlv7eiLgO97Jj9QslbzzbsygSKA3/L553
h2BF4ZQSE2ijkgo784zZFRHNOo2yShuUVrvE/slFwinVq2R0F61k9JrYxL9VWha8
UJMync6UI34j9uT1X8715qTLtEzEcFaNdgQDjbSzSSNUSS9w+Qz0y+4AQog3ckCk
jSw2938/DGEoD7L0zlFC0gU1G7pIZKOjpVNutoXQnIlAb+yeXWBDuZ5OcHAnqCZt
hniiKMb/pBx5+96AacfTJ7Obr121FvXKiTe+jwmCdBfaZNDHFKa02HSTwUSxOL7f
BqGQVV8WR9yXdRVdOa/zqfgrBVI+N1NhR36pqJTnuB2HH88n6xCFTiYJUSPcXxLB
rPMmV+516zJifGckA7z14haylsvHrbdv6V2sf0Hjxhi/iXi8xdb3K1ogfJGA/nVh
6Xpd5UYrkMHCwGlcYA+N6SnjL8t8fqNGI5C8ZVf0LNNn+BEqfKZyYjRz13+zY9b4
gvP2NYlGzvsBLdg/xYrwIh1xl1YiQlp5G2J3cuPH7GaMqIoSrkbL5VhFRg148P+e
zcETeQrZkZ8Le8MeVSnp5ZJ6V2rJvpcVGBiBJjCTSxEYHg7H9JSCkGxT/5GTPun+
yVZ1Csx9m1eY76x5Qy/vZBL1SMmNzM2rPfMccrFR3KBEByahBzTS3f42VblYyK9K
9bdSjG/AeNJt+9HrBF8LasbzQFXhwc0qBqzLofg/8R5h/tDLp2BHilRKu84mkVRu
cQaSKzACvJoX8V2695ke2F47MxZwOjDQ2Weh1iuJ9VmWO9AXrH2KfR/tqX3djb4J
wKxUm2vKK00Nfe7mULupzZKMZIUBhpFxDZpDr2lGteoBZuEdZim+QvMFC/AQVMp/
EZoc9vVfY2H0r4bYdCQHlKkTCknqXyihy/n/kqRLyrsrE1TSLNvpSSNch54RYvhM
IF+fO801Lt9aBJUGnjDTWdInHVX9Z067uIVpqMvcRd9Jmjr1Isp6dx9DFwA2BmqE
0RDbvPcVBSZIbJcq0wwrudX6GKGMilQ+1hZo7eVn5Hum51htBA3tnk9+a1OS23Fj
4qQrN3o7ja1T5nGVx3KtK2GpSYalgiAeReEiSsFt1aL/uPO+fi8qairejSXl6uI3
pn2PVlwt5HL67/dcOyDE9nCAyYhSwHRidaJLojz/MR8M91gJedQAnAp77ftUQAot
YpO+Qy4OkHLu5Ek63jzGyJsXnz8P1kMn5SUBmGSD5r+8wy1H8AMeFp3Y7HIdFXXe
CRdilyeUQ+A+brYyNAO5l2EMqkMotF+dk4QPHVd65byyJGfzyHPZbKNviQuRLcrd
zUX2MfFjT45HslI/cejwlCyegql5wI/Zbi/KnPN7AXbyxg8YDlUH1UUmv6ZQaD/X
ETgwFaapSw0HR4GXns7Uf41OghCVTnFhAUpMy/JaPTD/z+kfVT9/HtIa6AYqop+U
rOkQ3qwkKQN5L+yR1iBLDt5gCCVB89aRwJSFztEvGtHQ+w1O1UZ9x+Mw5n4kvUCB
uzKiD3G05XPqeCCi8YXAY7k1y+NXlAKtnxSDPWqfAYiAGv9p/qRRipEVzvGobuPl
fG6T2YJT32TUz0EYxwIehMpDMjr6kWKEZm+viAgN2HzRBAQ/Sr0ktq3xcUlQ3bsj
5PRg7+W/8tUrPj8RG6HBQ5mipNUEdfSLUyh18fURh128tGIh9aualGUBBLRQ1RBZ
qIendn8PsObx8UW28kB6zqr9LJiUw9oPy+KzdUpS/+8Y5qb9r0mt4ODtNLu82zd/
VPpp0ukxFGzh71bc5wzNHJxS3ueEzYAZ4u/WX9dgCUkrmrDSHFtjqAxC7c6C1zkr
01/bPmvq07SQ9QmUp5rWk+JNBNTbFgFCEFaDoWr54/yIHoplxPKuFl5tJbjZcMUc
iIxCMA+hjCfI7cXvTOUMBvSOQmZT7r/KQCdjHxe2DlnQolk7RubJpVrZlbxTG074
5keBIRZIEcIlt+FXv1Tbo06xWEA47KKC97iMicxUKOggJlVAYjfxVVIgNWGh9hgE
oKG+w1bHK+uaJa+aZKiuxaWnNnHxrcHLORs5OpSMtgQjeQhkiRSQTGNyEyvQj5oz
AaORtLYfyTieB77ElCGILMdxbPBHQJWfVxzwdheYaCoSYxRRghPtwVwyiKfzHUHV
HrrGYx9PxrCDnKfMJydPo2vqo320xc3wICjFFhvQgSjNayK9THQRO0M5ncXc1Dgw
FjTNd6radfdk3uhPLeGABCAddJo6Jrh9V3iBwnHJ6agdTy16cNlhJC4IoApf7IYx
NP/r9XQ9tJF0pnQEVub1o0SP3Uw9EopAxhBactFQ6//e2i2sFdZ17U9mcdHy70cu
tf3dQOREfr4ERMDils3ghxKwdjduHmJPkwih+QXeMQsU+qa+Eg6FzBKdosjJaypN
/+hhS1MHP4MVqwn/8u6x1AALnqcMcOzuLrIUVL3df+LyjLRNrdcD8gbKGeRF9e7F
MjP3j9GyoWqtE+T+qHf2DRvcWOWHZxpi8i7vE97bNNT2FSPw8sjds0srU1SWHr+O
SR2kWUI2f3oAlKvWuso/2/gwf/vLAyQrvXZpQaXFYpWWLTB6lUcEkWUBCjDpEWd7
ndsYFaGZE/8KE0rToEhaRpYhkkw8TJmaXLEn4XzCvoHyht71/mIEBUWcTNjdXRWE
96ZEYdSE8ylG9nzhTqpDHYcNHdek417ZzBka7aR1DHLntC9N/rHMjJymCeiVo5hz
ocTdtHVEjFsG9TlYg86sg5SNXKXVdQIY7Nn5bd5dlsmLdjU4tPPwaJBt+NNfuCIt
rFnrq5Ocdra6IELYTqTkYR9EOVE7+JqJePdu7xQvZrLrcZtu9EVWvMkmozA1Yw1B
jMXejjZ+2HObc56lxokwNy3v0bpvvfaafh3FDs0MojtJDY0ZQp0mKSKyF3lCXtE6
+3Ks9HU6K6qOkBhIEpR33+9z3ZwpZUdDDRR5evjCHxDFptAu8xxc3KFFIvt6ufBO
3BjJMKaC1omBWjrgkYZDSdUumpJAKzOjU/gAMqriP3VN7KpJlAkgOfD7TeWQFKoN
IG9GKoLxeT4kKUBEGMWo8FxF715ZRZxegEpSrzkmzhTR9w6M6zomPwJUZe7nqlwA
FLUtQG1ET1TkYNBy8iwbHKD0ihzr1e8lZ9byxfz2bl7QumgF7I/fav6LT1WhJKe4
5hffGQGg66FkjOWJtl13hUSSf+Btnc53RqWqLavoGq7zBLq6Qex7lcGb1mlKYhkJ
EiY65xwEAxaiIxgfJIjGvMXnTDyipO7SBocHSZ7a1EioTVvXexKT9GResN+vXFHR
X/lbu8FseYm1EEto0qBZ6QWxIevLIO40u/ihPMR/7bqhzkq89mrMeYPzjfdq8M7C
/FwHumkODkhS70PHK6vkcBE3nXIKsaEtYt2GKcBf7ECUEgZHc5c4h+w9sYKim3su
xf2e86lzM+vELEk4/lgx6jXnJtYbhFl88DE3x1BYU0B8cqL3WvvK5gJTsKToSDPI
UqE/HVRJTR1Tk3p9NuWf2jXexe5zWFGCK08PrUcKH0HQ6eaqtiVMAqRxiWcu3sjM
JirFaTbQTTdZxNUrRdzIuOcjJ4BAwt5aba1L7wtNnd8uFGTQVWLp9E0bwZ99v+TK
CPm+ClZJgyb+MjHJLzlLWArZdNELCOEuA4XWDiWxaVXOR0zyckEhk1K56p5nyzOZ
bcpv8KKFJ+g7Oqwa79W5owcZlpoge/Cww0HsbkkRvWMLm56G5Q2fJJs5wlVTK9xM
aeyG/Aujxs9O+LO4J7d6tRL030oxfnZAUllcH+i5YXEz7qvNCTCT+Lx5jGnAro1S
minGuMDFwtqTfE7bAD8pK/GXTC18zFypTqrPBLeR84tNamVjg0nrtQ3OByFC5Afa
VMPc3XKYTLqjAFIhtPk7SRrzopcS9aPbP3Z68pk844SYFH/l6mOnAuNIrhFtl7+8
zPHKlpgYYmnaGJA5FppDP55e5OFlXAu3vX88txYnwtKCezZjJ1XjKyuIZ/ljBCaN
MiCj4B5E8uzij3kx2Scr4AoHRje7nqjiCj01hcz2MkMKr6s5nAHNC8ttgZG17/NG
econziwGnkfsYa6CesZovag0FtKwIJszisa074u5wL7cqIib3Eodi7O3wEkGGdCL
u4667ahsNrujKLnPGeoTzzevj5Kw/WLuIl2i4AncnsKGjOFn56/soFZNOepP4ULr
hY65CjbGerGCFxCmFIzS9zDeUNJ9+hpSeu4LG3raKVamO7/F4PP3sN4S3apmpt1n
hQOxQ/NuZq2hf2hobPumO4kxlMIpv/evouY0RPgfCtFeTHM1y30pD6DAUT8JXTKj
7ct+Hsw0/yRLRaE/oTHHyxUH9NZL1I+qPwnmgR3tZCh+PBblQAyT+tQvpGqO5AVi
hLnJlrqz3uFNOoJPh7wi8Sn0k9KuC4CmpFnesGE0rZ/ccXTJYv47OO7YNeoy3aU9
+uWNuoGG0eHhPS1E9Lj/JcP2I1gegkr/V3Gwo0XtwjBk3YGyEyF2anY/6mP1RnR2
hU1q0Y6X8eJFXy7nHgJ8ovEQSodB2aC3gIYR+jAA+UOMtdgYylA6dQREExNkb4A2
r9qigL7BtZpurcmwM7O2LwueZ2YBEG7cHE7IWzorQj7KuyzafWC5P4o5EZBgly9n
FkFez0EFTx3eXBsgE6R8VvoG0MhvhaDdxJN2+X3WOsu1o++mz49I44mXc+13loDS
KhhH+y2MvhpzIz36zbaSdymISYrl+5w8cZk0F4s3rmDOmIY0+M7YIa6nPkzEZ/Mm
2QjIv6uACoFQHvZNvCrfSJh1rFY7EVsBotmiYJoFj807PhV1NDjE7IIvVBNHvglH
/Nje84osB45lTbnZY7WqnBQQl2owuRuD9ooFLMd96bSCvxBrmr83xriXCdqNwo19
JOVj354aVQsMm+YewyCsafbo8Q1N9TYoEGp8f+YaIzFx0Ll8TsUAqlC3CQ695fHx
iImthn07O49l0fUbS/4Q6z/SKMqL7X83Zz0JfdgyHnGBlOEP5emtGBKGee5qh0l3
hI41ZEAaOVfcfSaKL5fuNqmD7gdMnS7weKDw/TqHXIsGxtbzTVA9a5+c3zJhYlwQ
mkOe+diSo6elDT9+pVbdaMdEN2Y/mtQa8tj0ZOOPuLWGLj8o8iGwdJ+ctwfDqXz/
hvXnS93lsA6CrbjhLLjLyvJvMAKIZqbXnSlfOHkSC6ikprENvSDTqv+iJZOcT7B7
G6dwExArpbbflC1ztBu4StNEddTubMMBVXtdqd1wD6721vwWAXLQdSxpn1eLL62u
mT1wbWoLePCR03dz7jG3VTpDy3oqVmZWEPjKGy9UdhoJwPlNHYaV+XDBGv+N4MIz
HQD98TF2+eOuIGxXiRfSk19pgbqRucMEUZsVbx8eJ6uk9LJMqJXdSFMMA3+fIq1s
`protect END_PROTECTED
