`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
45t1tZcLRVjMzxhOHcRyhbr7xtOrUwNSsUsj2blL+PucE/c1B+fR9oovVg1ee3IF
YhQPMzMJ7aO5IXmdkOLzUusTP1FplyLSYs4kIAItbmGgiDQH57R2c1hNnY7Z+eH0
5TJt4z+MDp+cYd1AtJjd/rUQxh5VFYQB8NL5OUPnik4HxKPnFd15KoltNFACFFZ2
fEDTDzdWqcHRF4AOHKIuJfevNXBoVJS5B0od0hbRkiUH88Gs9R+05vZ8KHPsymcj
0FxfBdhy8ahvqECzPh9P2JaT3/J4yF1/G16MHygsrTKRwOZxj6Hh53YxkswO5dPi
JJX9azyKJctQYSSowsdrA7TqxNPcZuQEi1LtqNS70U99fivcHMWFNmT1SlmHeds9
7IPUubxku5srhJHrIaC+PQVf+hUNatDJOqN9nlL2+dZM967Gg13DS8OBc4F9KVyC
iy4uMPGXgedKgTbztIublfQdq6Oqme8bwl4yQ30n/Q4CCK3lixQt2hTp1KsmYNYF
Lx+eF1q7mbTGLEYObvOO4wfWruo+jvKR+RSpQejSNkRuHeosMFVscZczQDvOoMuT
pEol1D9QWyEHThejCuarr4wrWX15ZOCOif3s4LrgZ+z4WEQeiYZyKcKfSFZ4s03q
B/x6awpbhESIW2SURTGS6PxsF7QGFGN6jv+v98eMOE66nNPk3Bu7pJLDwjd4zxKj
26jsfVjGdlUwLM/7S4KHSCqmOhwNA8KohgR8a2Foyn2Ncpbc9Z7WKURn2CMKNMA6
Hzjho+JVxVtl39K00swcUcTiTBwRftYQ3esePEjjTmdTCm/JGQLpinUAaekUB+MZ
Q40J8SJ+3fxnLvtFJE5b5V4thyZ2Zumj1F0jYDX9DO0OuoTWzVDsibAFdBErOuY0
FSg2xMSijcawGkuBeyRzErhXOyF4uK/2zWjxxG1iib2c4E1HXoJcf33PKyWiUpJT
ez7O7zGwRH6Njt/BWup5IKFUw0NzrF77unTk1lHhSbEgxjyQv4WiGtIH9JT5jvOW
ZNaJNmsTfnZVbWRUpGcMS0OJlbm8q84O86OY+vfrylXEybRx5S+5n9UY/1yMkObr
E70Z+rfsx/QN27RZqvfb+fvcoPs/aU+qyn9dUouDX3MfqFLcAvr2RR2wpd399qfU
KRKYG+TxgXMn1+pfs3MVQL4mLNwokkg/nzhbwZrgqIbFz5kpRyPQsxbJZkYMv34a
+R72kxJKnRMwx0UneXxnwVgjChuAbp1LLuYDrJ5d/OjOeCrlutXcZMaIF4NwGIYt
KhS4bmpFCoNckDki/7Kclsl6lTW1baTwihFmQ8le8S3tRwCacR3BUyAXOQAMzT0W
9NGiqGNIWskbePO39UloA1q2qEQA/bRWmvjBBTXpdOYcib+t++doZEtFaB4SAD0e
k3VdRnEJZ2agJgPPuvM/3X2WR6gZgtOegW133ZCKe+MUVjjJ5cLOSuSh/xcG0zfL
ydNukglcWivO0bIJeImXkqgY4GQR9/CE4kPIsAkvaoAX2zyGL8JaN0HzdlCiMB93
FnBQhOK791CJ4mIDDgji7l7/k3/aH/8xLiYY4Fja2SY=
`protect END_PROTECTED
