`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NfOoaKBg0/apQQeQIAFQgdXn6ydubBZVjk2U/hlJlSJ9LSx2m1Ue1vyXE0vGeLyr
VkKeca55qOxUjiOUZBPGYIXLuDA3wtavf2hudyAMKIPz0XNJ5x2tGphh/UZBEH65
V1QQ8/t78IniLd5qph27JNjbVyu+G2gdZ89hEAmUhD3iSXfrsS+6g8tgUFfBeGY/
Hy6oNS+WtqpssUshKimUzm4YRZgtdUGVt4Zbj1/zuw8kHn+uuF37khHuH/NqWZFU
EAD9IlkXGVqQNUkbaJTMRTaLKYBP1J+qx0uUbBBpBSxATk8iZ+Th6426WnL3Y7EO
UnezgSfPkDmzWGJ2m8q+MdinFCyohFi1zeDv4aY/J+TQChZn5ydJFCAkTH5CgLnG
ySyH3dGEcs87QadCRDsyWIUpRkncGpetR8KC8D44Ios=
`protect END_PROTECTED
