`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vkBntRiNLJcQekpJ3SdbPnoK7huSepxzNrk3ykfM8z3s6PZ2Ra3WSZpDWfDUvykh
MmoKAEsWwO/C+ZhLvJJvSsMszqClG3Prubb5gMnLq2DdkNlSPa1O8xsTvakQyr/W
7yffYliK3VcTScGU/lMO2dn1oTRJq2PRxWIxD6i9UmehYDbCsg6EoFdIrAyuTV5P
IVOSi7ZI8kV/QbZ7SFGtEzPTaMJm/mZGi40MkmTMwUbfTp71dMEtoui8bLar36wY
N4JxRjOMrqkNp1d/kdpo2vB8quGFx6z46MI7ulnrPZI+4QYLx7GjNftqGOXqQ7mz
qLt2rBv1BiCAeN5Zw0ml3vaQo5sJQuP84D5YzCIjBEtFSiAwovv5b/wPPEWbtHGF
KXgthSodZ9TjoAESm80CHOOfQnUEhcp42tQGUm6YlZT2n2trCS/1TE8O4pDq4a3i
1fZJ8sxxpyD+2NbxyiTErh+w2jebalDi1g6sdYMd5z6bd0540Kl+lmSvnHrTOvrq
C1ikf9uvn1tovL+vrIO3cXyxfVy6+81oeTc3+uA9RZRsFtk1F+U95M9M2hgqijpt
Pxp6UYeR0ztN3j8O/wlhY5bGtXDwXcWucWMjYpfqod1v3b0KH+Is0XQI2ssGEsT8
kX9LLtRZPIX5mddJ8mmhDymmbFV1mTmPFknL5HhTdN4Xw5AmTM/V022KuT2e3Bog
tuYCFZTIaXtwjvyALy1wUCqxp02GaN74VO7m+g5izSv/McihwuDHLkwUDgphz9xV
iwp4Os/45vmgBNNu/j1+5+o+IbR5zDtuKI1PvbP5KsPUc6EsJ4YDW5mOD2ZXIhGJ
myUsoblM5eyJn2eyNdU34r1ChQBvNkcyFH1GtPdCmsq+U/jGcNN3fI1tydyXu2/s
O7cW6xm5uCKoMd0bUpWJIG9xeMIVVtjRk50ib7MJufyMRgUt2K9mcMc0j2Rsu6Xu
iS0PJs+ZoGnpeM8PzRWbyXVsKyZMo016eLeaZxGfY0VoKMMg7nHCRMNlwOVBpPGK
OeYipQtWTLYMy/EDMsBQk3RKztJ7fyddgXC75rTFo4R3bybssN4wM2k3DpfJUjgG
iNmt91ylZPtf6Zz/YPMFCxMIE/yKQYRfsp/p5+T6xqyGP3Bildis1cW6OHt2ryqg
eqZ5F8OQwoXDn4WUtAaLPnktCBx7xKaaOiQb12Z1faRo4PNcQXW70wwKPfBAEQkh
JCv9M1dWNG8iJgjQRYjmZfkl7m12vfXG3Zw0hY1xquZ1UbtLzL5CgUhyoBr2Cxz4
gUkPU5yrM0qvAhfw7tgu/oSwkCHJLYUy1rbdRCAmUa7mUsvzx/OaNJ423K4GBt7s
09ToBg4ok3fbOCgh9cJe+tFkVnj3d5/pEqF/LPI2Qr+8oazXxH/BxFnCJ+FxEXO7
Slo6jsJP1lOeGBBs+OBYth6E0G6V+l5uqqfddsGQmrAKdju87h0jOlSNmxdfINSc
/zQngXjlavirtCVChWC9ocemVG5OkrfVSSvtT3SibiJipSOz6fnPmP7WNbBITvMP
pn+zqkcy4ltivYnrrFXVRWRvGuN4QewD2f6SNy1Baf4dXkkA8Ym9ZInsreXEDKKM
JvmqTqKGjnHLDl11rOH8/bbi6rq/wG8mSYnEZEgq3S+R866HoLnsq2NfM2mO8Y1s
bUTVELtWU9jmi2sIta+pQF5/RqIt5W2PHdeTlXYLoQNTyPc3aDlM56fckW4Flk/z
LD3FBKKG1bpObwKjOsmRAg9VCtJojyAflDx0wKCRXTq6rEi9sCwINEp0p6QV8zd8
GjzWU1y29SXSl6Z2ASvWFCvF6IsPKprxwEH8QvrGzqzYOKS/3Si49CQSUBBGkMd/
p7fcWxGjxYkcoSAJf0KdkBNbCjklo/niwXASFXzeDMSGwRJtRVLp7k3ynU7GSLTI
bqamflQ8SUvRkYDbsimUFW1mw2OsTx+MgEJ/Qvb9+ObZWty7AiBki8MpzH8kUDIa
0RIFYIsK9W72i6Xl8oYz5cfxSlCezYqlyLuxDch8WUfI9qKM2BAAlZPoR7BExaF/
ZiiTovt5RL8rL9JM94NWh85RE1u+7SbTdaofNV1GT4jxK5H6IAMGyaOzwSTr/U3l
zloDfihUdoo983hXrO6O9Mi44P/Kz1+JxkPzvi6600v3zx0VHR+avMcr17hvi+e3
pvrMwscTJZCdkiEe58wPkqd2aIfjpy9w0Eyut5DFxNeXJX9AV8ByaGYVCki73SLn
A7VObueJxd7hiy7L2RhDeeDFdt88GDs7+0AlrTtrTsRnxIE07NKxNN9+YtlmK1Ti
J2oOKi8leDfKZK/QSHhkkOMLVL0oxSt1QHG5Cu8U+yxLOiKruxqb+aWekFtNpjx2
aegh7MwhA3Mm9LCpgnr98UbVEyGG1HWXj1cIoEkWgW+KM9BdO3fYlFwqbF185VN+
uzBMFF+Jq/9A/qQCj4ffStEhgy0A/XkdROrw6tsu9KGbE5PN5C8ot2tDp5x7L3Rx
ZRXY2KO37yU6WIO1bGy3mj1lgHdvkCfudN6EQnB1RoJ+Bry9VPP1XYZLwIq+bYaZ
8uRVQU51chF5uMe0cnuAxLLT90MLTTpQMeXPGIPa1UvOnW87p1mt3tfVWgrZZwTT
HVG2y8OUbU0a69DSx3O24uTIWZ3YgTe0lFFRfz+HUNMELRXt4xlAqeHOnYImM2kJ
QVxyZeVRCcaXRinottiAv/6f9eNQlWmEp5qH/RLT8lTlIZlBArK70ASDjNAX1Yv+
8qLdC6+1WBg0VGOF3uNMuPEIr5qLum0FgbaIWAvTMd+1NaSCJcFyCqgYHSES7llN
qgHiPq1jxXR1uqCtwKrsj0f8J0ANl8+GSYmSy5K+xJYJ3/PVd4IJeLguinx/NB0d
FuI1pp3IR+PkcF0NN8M2n8eBiM7VBCxBVgVwYlQrfU7NoIoGoDs+tPUAhR+YCfHj
Bzvzi9ao7+7+v+0FDApFyyq70g1WcDvgFi520qAASS6Yj/oUjZJ2qilkZp0MnTqj
BgSC4SlEKPXkOOCV/CBDlOMeO3OHu2p9Ib/OC62tiia3EBXMDbTaQvE0v/eYh84v
lE5NnPCVAeplok09PHta4nabUDJaUOyGqjz7dGLkLa/dq5qW85vNZZQwUynY3faP
df3MP8id7vS6AK7CzE0tuswuYIpv7p1ExWA6jRS28ZKCv4tFpGq/52Ewtl2Cwo2Z
Zy13VcT8dmJb9P5x6pfogAjO3Lc9EBSYJC4+Vb6FQyvkfp8t1fKWm7+G3BN2C/aN
GeaV5Y0hT7nMQ88e57+sE7fS/3d2gw24PXRoPvupfT4PH4Mz6jsOWp92uDaBPWXW
+vPXqgXFsXIejwSp2Q84rMO8Rf/uYiITiy6qycbWLFr4QxHqxHkxEE9SrD6MJKtg
UfeYzPIZOmEkkDrlusHh2s0d9d/IS0LyWOsl/juewhtoBYMPHu5vG+ifIGhMPfuz
83Do/DsY1qsnd6lRAVyh3M+3pqC4s0OvQX8S0+dP4ksHiazVT9tLYJV98fC0IbGD
lcqXkW9+nIW99poRzo8Urh7xOkMonPv7ytCWmCeKZbVFHCKbUo0KOfw/vsBZQZfl
CTXY4dlra5uynj71U9Nj4T5ZLrTI4tArlfughZCPBjJ/ql/J+Yc9A8G2FUD/A+u2
SVHGMmw/2XCE9DGWCnAJyiBmPDOLH03zyLPkjHeLzJ9XM3EoHay8TqtRBtiHcy0h
+l/eV+H0basZedBxde/qvE6JnLiPYAGcPdpAw0r1pnITDdIu1Sz+4Xzc1HDFz6AD
RhkEmHiH99X8ONHmGTbZqekJedral2mF80A4e0fkZNINKwx/CgGK92UEflntpZAr
XQKuv0UfC/eCuRd/DxZfvjOqQRAbiS8kfpdKKcz/Ucih48QnPnzDMdzaGvQhT4i9
OGMcpG6jlWOKw/5wNvJ8ZBFRCnHiGtoW5iiE8rCdANPzHZAsH31AWzzodkK+y+ML
tSL38B8Xa/51tk/POkYRCpg1wNU9zlUgne/6m+7/Z3pjps04FqMWojTFW82XQNwK
QtH9C0RMJus+KoZYU/1+SAS0BUWalvBYJMsuA4eRPwMIT6s7ZgfG2Fb9FP/UGMnt
KaXhueEXYr1LgwxsdgOMFaPOqdRh3VVV1fZVO2cfXzgxZhhXgAe/3V75Bgt+FAkG
sqh0PZm2yxnJw8AxfP44lCNG8eqNfn4ZqwkZtAlVcIJTsYvJX+CE40cCOR4QeFKU
q+tuwktn4y6H79YRA8wgmYM+Y8vvazelO+TJF2PKOmMpmfl6bGYl8gSzu6cFavs1
fplGmsot8WZ9OfHckokll+rdzMQ5NmX/M46ouBKzrbPBRGBQdWBdeImolnL4y0uk
bMWizpeAKq9jCwsH4YWlATOL42EaTf6nrO42DXerFU+ehO68MiaY5om+gQ3+WGvQ
Xf2WLVt95rW7UcW5f/zYQeLWA11uq/IzHzQfgd9qZImfOa4InVpI9BvuiyXjgEPW
9KhOj2OVrrw96vDZpqPS9gqO+bJrV0YrxFhQsOcxY1zftNxOC0dcDDI1Oqy2szu+
zNG9rVjOPN7P8TKT83Wi5oKaH/aJ0cafh3BL3SNsULqMvwUOltnd8qQymgF89EQU
uwxiYGgynrwdwXyBx5KnYoMttfETT2ZjJ7AN7rBmY+wm47BurVw4p+zaTOPixdZ3
T0lMWcZVTs+RjSmBU8rhk97FcMoXq9rYDP6f/X+cj0YHeRotTz5Gt2chEFt6yJL8
zAdRIm/ww3QRSX5F5+DxQ/VQJbwl8tYUFXcAosl94rbJtj/cCDEzo5gDccBH/+kf
chIwWztAnS1hussgWrstjEDL0v3LMB4TWBHx586lxzso1UEN9Y9BNIXeySHUuGJi
+BM8JC4PQ4RAVHJqBkoG3Z+8Ji0rXuC2BXu+3+PVaeZPUasaiYx8PrBw6UU9No8k
X7kI4Gk3XSWjHWvCNV7MKPJKQ5FnA8isecHE0cVZKC5BAYqyHTTaeKUXPGoK9CFp
0XyUgW9MKCicT7OtKSF/xfMUnq1NQ/aHxz318bNfpcabxpWkZfV+j3kH3IqUK5jc
IJBjBROrZRdbWbgisjF+oH0LBmV5T+kGVXEpvej6c+LdoTVDO5WjlFw43FBCr/2g
PBVg3dgYR8Sfd57AI/sPkeAKof88H4upjgcHWkNW+YV9MH9xHtJE07Tb3kEYgBcl
aCWAge1WDuzUeu87WCo2oxgKDGPO5Ay8Y5jxy2k8IiImPGGmlPSFgJiHYG5alz/o
ie9zPNSKzOJXbOiMTvi3ykTpIDbAtFrg+QBzkIGfImnoE6UctL857bWXsoljV5iN
IKf33idaMikpux3JUhzRqKrtTWS+wvax345qu9s8qTNh8hUi8NcFu5r4FLCKt1Xa
VHk/WW6hpJcHMmPKDaZ+QBzNbKFTHIsa5FJcWnEW2gySE2oJLJQicJgESwLTSmiK
BZfjJz3IJqj4ReYXQe/RMMvsSw4UaDCO1enJtKNJW48VLJRiMX39VcvZSgfs/Llo
GCP3IYnrSswjS3v7slaIYWkHhLZ5LooeXdNA5nex9hQGqLHyw7FCPeCSji8Obd67
phpVH4d3hMjjOM/i4TrbI/h7yZmeTAt6HESYhV3ZCfpHWfpIgMRzgzHIIV0bTnVx
VAoqxLqMEWTTVmKDVpJTfddXCqk6056akZ9KQkUIgLp+X+AbCzQ6/GaP2gxMMc6M
4A3GdXOr+3qURezqkEJ1mFzHnHujES2rqx9wLpCYIv092ut1vGgeO1aU7FI30mF0
FZUEaZdnTkiydV55QPOqpTJfqSrkxzuk/bvllN0u7dRkftX8IKX2fADOLqLUOKr8
bUTRzusQdubFP6z4ziu7/LFEqZM9F92zkTMfISmTdo+XKgTv1TR8rf25w3xWC3yp
gj/L0wV2CAeMhfExSUbWHKCMixiGyopHxLaBK7J2qhhEaIbCbmug5URA4rpBF7VW
YleSLMwZCjw19DG7rXCEuNemfXd4kyLVzcIK/TXZTVKaE7DCVX9qOyOvS4Eb6+bx
YhP8YsQWPZHbPBLCScIdchEiEvM77gxoK+kh/nK69KZoeArlb4GxWKNlwyrKcC2H
4kCmeWo63Na0cMUQBnFbvcMleleZWefz25UaLw74wDepRseHYwUheF7n5tL/J2QG
SZjcrfmFl52MfHRFc+r/4eOEzADagBCu7C2CGA01ddpij3mbly+cJTOjOli41RpA
lrMgHvPXJweG6tMjGFaN9SEPK+UYnlanBXAN/+k3/Y7yGu7pS6SrxwhfZED7va4Q
h08e/M22PfzX4iO8mAWQ1FCMAECphvlQbFkS09Tgq2nU1WcaiMZRbq5aS1jpsusC
cgul0g1H1AVVQCOPyzlKzHV2mQxaY0x/i2UiXOhBtnvDHehXWB1u5Vv4CUhKr9RK
t5j2Axcgn8n2f4MdWBIA61CcK+4oDPoe6/hfHd7uMtyR12vylbMdxmYE5v62H5c8
NCSPxqtI/M+DB/I+SiLhu9ZyX7KrbpueKtq32dPkPVptrX2iKrmGzZb45XhnNnA8
GmFOB02MTs6CGO4ido0p81Fov0hE0KjlvccrXCz/dYlJWjAV9JtGrFiKKV9rSEfM
efv/mbVGNwe4rz/7Yg1lR8kAIJO2QDEXzdqTUnyE3UvucG/kDS1UzC+oeXHvSMVd
8yu+So4vA2hoOrT6nEQESNOrxF+9l1/RPlGuRm+oWzM48T5mrVI6GiPHTqOkz7Au
XW4d2wwO01usN6KW9dIlG5BHDhrkO6Moby6XD5ZzGV8e1sWbv1G8+Ff9lLBOAT0/
3s21WlfKmfs17FEvxsHe2VTNqJ5Kp0dVD1C/Q5E1BRAlMWkM1HzaXHKIo1sebp3N
35pj2fFFk/bo3BQWHLZoWfC1ADCu6MF7D2aFtgoth/H467hsAumssTQnx9kPiiny
/9qSSwPh9SSGzJ1qpItAbhzy0BT6NU2UyiTc4TIiDHpzrpqX/mkgQ3pWIXJm0leu
z+r2cbYmk2fRg5/GvGuJg7Xd7rAI0GoxghC46s+JRsnSrT0YC3jEkSZjzI4Fo1gx
VxC8acZdO0bMk+NLfJck6bOJAESon0FvYxK2e0KnK+LvF5nLpnez85Vc0MuW798Q
+c59ti8YHZpr3wkjii2RUqDIwZ7l+d3Zw6QETqAKCkmPlH1GjlPgeCxDsmmSFNh7
UeRX+40B7iQDiHGPdw8toyK9tIl+m8DmJIhYSWdQ7yZ4M/2YleqhPz+8jYZqNJHY
m5UDoCEqevYgUY07IomjmpcUMRSJP9n+osyOH8yiKKYfE7lhldF56SDyQ2tsz2eI
CdGaPC11InvTiCMi+5XUkKqvGEnPn6F9QX/PVuxLw9dKPXrEx9JkhzcyOAZMYRvB
Ol94HdR9gxvzQyl3/NIx6AORB7CkH3eGbBLbjnWFDRjvqv9aSyEogFzUrbAy2rzr
uOx8N3+F/xa0yPAkT3OBHwx51nv+mpl/Em0ZW6wFEpocpoHemNFnGnZU0klKbuXw
GQ2Sdrk037yKEJzGDhSIDnsJwhgfl9PzkmWqYnLTl52+yJl9Abs9GPBi0mqn1adp
iirKZunXR6BWoYxoXE0PRcpC9tgiDHnBLUiBp/ZP79gNmOif5wS0sNmvV2uN9Ygh
4+jRu9nhA2HtWCVtXnOn1/nxyFRxMhGQkBKUcmSS7PTtLio0+eao14yxwm8V/WJ6
1ZY0qTnobiD1P+vHT+f/E5lU0Nnmdzju+fW4XB39Ybx3nBUxlSLZn4p9sSQ0vExK
LG8Q2AcHJbtYVAoXqUxE1cKRwd8FjfsJF5MU+4eiVb3FsVcZb4S8tC6CPWbuAaKF
PkVGEmNi2hjz/2iTb2vHARDUoxmr8VteQBt8glbAnpAMGYikqzn3BiOrSGkVtKPE
RRaWezdmUCA/ZDLZZaY2d98XMAQ8IKIdTPtQCtRFkXxgsSbiawC++kr9WzyFOH2A
KpoWu68i1lzszrlQM9mkKKSH8EVm+I0xSnAOW7/gmTUk+v5/4uRVqssPMyh/7jad
mrqbSpUe0CQ/l0cviYrNU82+G29J0aID695oKVtRNqb1vaMNjuJCrxjP3Rqb29Z6
lwG+1p2pA2YmwiWLNQlY8D42hysdYThDVfO34EGqzPR6fOmkvoJyW+RwoUvP9mEM
eug1s0cUp2YR48h4LCMdl4rRX/l/asqGeQv04JNEh8itI6k7I37DwhPrkelCVCUi
eZdi9BtRu3zBaLeU0dzaq8HxttjB88YzBzhxjU0a7+I/vFVLMEI0CHgkDTRMHc2O
+bTnXwLLCudEpppN8KBMk/uFjdBQH/t6FtAs8SGVv8Bb73XrClKuc1HMBTYTP04H
hcE7jvrrLiGMFpxNkNAdLulbTH0OfJ9L/HiI5FtCCqaIlSZAzx8c+SStB8l/mXYV
9PgKgfgovo0W7fURAAJ/2h3BS7/sH8AAlz/dUNB0GF1bcdycTrrxwOxSR1wrAzzX
ikucF/VM0yogpDmejLzQYicYYOPiJ0kiN5w3/4n3NTU6LHRUtORva5cjvwvLi3iA
jfKw1qNZKP9IxCXPbEA6FOqyO9tDF7vvbwXoEsrE/c8hHFlsftY7AlbteTV4a1EO
DuWhXSg+FhWQN1cv8rqv30NPwjjYPMI7CzZ4isKiXkFCrBNGzil8ZQ0EH4wQB3Y8
ZLUuPoT7ov6Q4quPXBk3F768bYAhBjWbf0qWboRdao8jpJ9hZE8aEzwWKz2GKe8g
oOG4pQ9sG/GXPl1ICB+6hgAASEBs9Xc1Wt29IfRl71pn19GtPTZLEnXQJbqSZgML
+3Ge+3zJDeWWkJ7OyzB0ywImu3w3bV5RkkzMGAu4t1W8m7h9it/0KU2h/FwM3UJP
yBneh698hbQSEeGUK68JeqyAGQZFEGZP1OrAc96d4aEJRjZeLxjkRKeHZdKM0n0T
IW7OaFwhXEWVmPk0+oX6AwsBkcyvYQ372cKUBmRXo/RIcsqjASnkYrVIqCuafWBO
Omtq3ZdqCdx2w1gyJz5Xb0qdii6gVf2GhLYAeXcz/I1VnSF0NtiWYko5C8KemYPQ
dxmwbmGSaFMslvJn+yScljD5aSrS88VPYuWTS/YTRqBrc62pjCl4bsafoBcr9OY0
xP0AmqJm7yRb0bCxwxyP+B/gfTaWjEuFqsCyi0Fqf6iho5jc5yu/WXoUdOifiEsK
jLmw8XPoHzP+O5FUBN9dq2FPo25mCQvbQZN14zhQ2mlFkhmPsfPxhDBc0BFM+bKw
MxRGlWuSUaFCMAsXBouKB0qxkOWRsfrj3VpS7yYzfkE15TUGD2Fosxec3fZAfW4c
8wNrw4/ZSxKyfB4RPNcmeySJov6DJjK1I3zjG4muze3YnUrt9Sn541nPstrEidBM
NLKFzmzXst1GVYiOQgyuw5DTdS5eSM5Jrq7utz8Qa/fPITrmlCp3DyIzBwKGhhah
YD+8DAxuSApY+/Vna89DM4llwY6eDmStDK1iA/ZTCQ+HnLDgSUtE+zq5aNs6dMdV
azShcgFpVIRxNIXD/cJmzaZLK8K4/H5LcqLTo+muSreff6uBon3Z95/ePQsHWVC7
+cUv9dgGeZrx6HiWnpbJZhgm78AhLpS/4IF9BWrtcRLkcXI3b3yHm0tkHmE3NIJy
u2XYU+nyNxRBEMhlhhvlibOlU5zfXQj51lgc21ltrnV7Uess8tqzAeneWum5dK9v
oT1aT9ihnNV0wC6VsZZdI0Cjmji8McyT5gwZ+C7NWHkWpbOQQ9Cm3Zzld+L08fIU
jZC5osyWgaNnwUNO2VjkzA3om04RyW1IV7Rctwon6TMWlmJx4lpZGknpmRI1q8yL
JqtQVwQ13xrhHo0q43+LIYpgTUP8iLiJESKrCNOWQTTtTT4/9CbFMGNgjGBmxIz5
XM8Tl7UBhbcBdfsHEYoWN/uromCqU/ItGp34XGwj4WduvlSB2L7scqOk+MpZ0Itr
18Gf5Qrn34osdlVFjJOIKnr/y7k2U4TSnUtH9RIrrV7PHc28yyWo07drzY81oyQy
HynVntCdhyr5gA5zvTM5KBXFjNwycCCJZLbSOSSULjZvtzWU0r/BkVOkGQXa3zJN
7TdCGc23kWWH27x+bTPKAVelULQDk9Z5JAv5qyRFYVTZfL7Jwb46lj1iF61TvhWh
/pdtz+r5UfcxKY9cYIA4wqswlwYyKBOAGiTBuKKgmjwXxO/29r67s2V0H3lQVymg
EWbo8CgLjTTm7swMyeAf+5dmcgU0bYoqAO1xmhiVSlZFi9mazjMVut9t5tkaojZO
UKvqvo3uGik1gvMoSYMXdRVjNnxUucnE6uhyAi5toyaSn6UUIzaQgeVcJqNylGOI
KV67NGaUV2Ehx6e4uToAzggFHVtSg7x45t8vew+ILmt/lXMKU8S00Jhwttmj8YQz
MbDjAYd3C0npvwKdleKghmPZLhnHWLO9mtslOVRe3pMQ+pj77HdlqffgmkoCQfdA
K3kZrMqRmnarQeY+9DhuqHx5ayjWU77nZgeAKo6S8FSblhBIGv2oVWLBcaRKrrZA
nfc+rN1WxPBOf4FBGLlKhL4U2Y0oi+tHuCfSHEFLFIhx+S+Jsy113MCyg8S3gnQk
x2k6lGfNmGPLHcrGN1Dv/SeiUMHNI42K4WeY17wjoo3JbzJ839oG8nG+MvyMRWCY
M7tILUEbdjEeUFfF8NirpLczWM/GO6B1U7rmkybhxdq2pATWceH+6JyJemYw6Nlf
bkjatIZaWilP8YZ4wNrQOLIO+z34UWLh03HRNExLWN/NbhR3zXp6RPRQ/XUyG6X+
+IQFh83XM+Hguqvwvb/TTR5HhUpssjE4zuqQcGtpUWjkoMO+OQVbiTIi6y8xe/G2
jKTGrtwE/89RB1k1/3BIBVMr0bNGqpXxfGMc2D4qqj2Ymdbe70yqSvhKL9sbpbCN
U/Dk8opMGNYpKiB76pDfFkR6Mag6kYfloYFAfSSDys0Uf4frf6OswCP4MT+FgATV
FXyKpGP6PfRgeSlk3ooAkfdNgeGmRvNA6vQiP1fv0PMQWwBowO/07b1N0MLMaldH
3u/cgZgf3HWTk6534NdkQa0zhLNXP0fZIaeEvNV3y+Z4E6VGG9A039mIyyD91Rfl
RZkXGiotBF8X/tqLgntALxfg8rg8QzSwTBYWaCOJEs/ryv4aaC3xyKpGQ76YLS7M
9jS7N7DbSvCyzP06EqR28B693ywJF6H7PRLTCy2iCaKnRRIQSkvZTeHJyHqT2371
wLC+OcodOI3KaLqCNS+IOD/EGhC74SFouQficAvv3FQRRYfuDHOgTpNa/n+9eERG
4sdYpmuEJwDjb0AQwbMo9FcacLoOmwJwaJZf4399tdeH5vMlhTYzklchpqk3C+iG
NH7KjK8/jvCwEdcNuEzdg8BbYFCQYAPn5qGqWJFthyvJCo4I5yfZrYD7cAukSB8T
nZ1M8mYhaduHmt3x+5U61lVamdFfxwzbFQgL6SKBm242CBhsM71LvR1wRGeei4u2
UYpEME8jdc4H5R839ZXSIA5oMlZzGvwCG3qBPMBn6jljotmLkMPXT4aOpvWJutNl
wqz70L9YcL7c5IbmjGH8LVz6tRV9IfzouSZZeoAKnhBy8nfBAnnDSej3XZY+29vT
/6pgtzUw7LH2spH8pFScVDJYvCKbUUzUXnKLf8u0HiXtEHITXfYy2hVQFn2HqTXi
kdDByIHmCYST68ocrdnU6m9J8difHsJEl29cnsE1sXZkwtrIAOYgu9EIx3Jyhgmw
ZGOCiGMG2OwdkkneWUCfebfRqNu+MzKdrkLb73vtlUjIVaAL36VwQLjxq10Qt6ws
ejjvxCqG/oWJHzzkXCYCrBhcUFy57dTCcPWu/WLnsuyHuffEVARqFqD30F+YqsAZ
mWpkenlH5p+6mMIkEcVwa0Ut3BL3VZfZH4n8NgNKfo6pDWQiUDBMUBrBTEJI87TT
EP0rlR8Wy3FAdmfYrzg45pZk6jpiZiEPkWiKuuIqf0AxZcDH+OUyipywgx60JuRn
MWnPRO2GekwJNjKBHF+rgkkQnDsvMdeTD34gNjYc09ozJtwqbjpq9aTiKp9kDHQh
RrqWQkUNFqRYeOFWKDgxeC8qTddZTIfAPjltBxqRMTuQ0bt4eeQWyo3X3+Fg9q7z
NBONesgD/XuBqQpGP2HDhc7rOYHRvlD7PXY2fbHOAAHf/wJI0slOCC/mRfEc4Hyf
eIi/Rfsb1eer4x6Rl474AXOJmaw9WkOCPuX45N9nAGFUSQy/9n+GmVS27LkH3fCP
roak6SlXVowu4M2xAOpMcSkKXfwZgVoIado/xiBRpUlbjmOe0+V26zyc74G6BVlx
erFUdxmLTgKOBAOrhFLF36BBL9jTFsDp51gbeOQuCConXqf/FXRCkyg2wy1DDU2q
RZnuiDivfzfaHVJjo18/yVruSw1+i7+yWDTbuPEs9a7KJFsqzIJvGkjfdzm6jIFG
kA4xu/cxn3oWoRCOzAGvBDQH3JhlGAuLjliWrljQ9ZSFDGySD6qIb38HmI1rqoAe
StxRIpRQ4XTM/wBygItNDy5l0Hj1Zv75cQb7+jghoa+n3De68Vgc/ZYzTQFWTbmP
cuf+xrBcXtlKDDKaMektwtrYl/3bQrEWxKj12dtAEmFcDHb9E8B7fPBMKlX/OQIi
9eGIfYGGlcdb05V6G+Y2QcyXhRrZOpF+gIZP893XSC0v14IaCaDFPE17N6ZbYERm
MmSQ4r2OyKTcGTIDlAj4Hk3alaXRQmhzSO3z2VSohxJocduiqlI6kZP9ubWKqF0l
4V2AoEPHl89eMzD7UPKj70Pt1Tsf4f9Bw4e3UNOSuKnPFwNBL+sT5ij697XItigz
SArR9C5Y0yKJ6IZJ62xqfdMu3Gek6hNi5jVUoc08VNRptLEsI40Q7canPB/mk36S
1TM3bwscRKw9jKujx8yNlwyCo6ppolg4jmVpoBdP7V6l5bd/njksKd9t12ds3GHy
NkTlTj1NErgbDvZY89+8V9PnEzaf++356cBtA+9MW5iwQp1gnDztgcE4KiZZ+lLg
pmSKgV4PHVHxEcUqERi7WrVIJ8PIlLgAgbqz0T29pXg73rBJW5M9/NNt2aIqNaVW
E0RtIS83j4d5nWbuspwDWwwgm7AystSvkyC5RFwf4e34vQFw10DlnFoFaYNRuTVY
uKAKSp9ARpxch9LQyAXTDnMhNeFBtkahBhv9LqsaYXUzHBBqO3kMV8LwdQMfYWQU
nM1JTDwyVWIJ8fcMaahvcelYGTPf/lm3k4Nxmv2kx8/127EqZIM3ow5bTEgWLxog
Iyyicr+8K9bj1kFZaT7T2W4X50S1Jw4Hr+R0CHHf6gdYeqjEfAcpRHcUXTZQ8ARF
bDSmFz08FIxeK2DhoUTDqTOo26huOJZ+TDHYXefDlnNw8XvtfEh536kgSzWZs/Kk
TVp0SbT8h9tTTQBhzz57r64Xtno+T3gNla54BhwtekH7yY6GQZniWoNWz7KTuSr1
oEuheddrSx7DBLo9kr4CTGRR2NXFT6Ubhr5+swrMksoKI2QJJu28Syo6H4XWbf3Q
q34kgURbG0zrpIHoiA61h0lzME1qO8SQdS12GGJYExSf3ZNr+47CdfZMUiujfKgY
IyyAx+mH9raT3t3TL9Psb/pTTJPuFhYCZgWuTdyevdaQPoOeRh5QAnyvp2tsN2X0
7Pyhb/zqJopAmqntWdCksFCRbGNi5F1MVRWMul4ZdjtYqJx97FewkhvVjDm6cpBl
BYgY1qNPPfin3V0fxbLqiMNftJyhzqRixETNFcYr+91EIMKCmGA1oXF0xjgyaINm
Tv8UEIZ+CVuQwz/JBX9GUGNQLOztzvpjJBs6UPC7Nt+YIx+l6sF+mLnpY0lMrenU
vvqMORfma4iRqgwSfvzIr7Idl4W38uIiBkoUn5lHEidCMy2yTtbcgfDuRsGA/pMA
OJBOnptVkKlGsFsnegARtVvf4E65ZdUp4wfPpayoxZbKxm3slALE7vIcjBSSNOQl
unbXw0ojleRQaul26hWgybmTGiXDmy0JMPKDjA1kcCaklg5tV4sU2ObUCa+OtTyo
dNEuGkYlqbucPQe6NA0x/FeIKaiy5DM0YZq7LmL/9eo0porANS1Sy18Szl6Buj5Q
wxbr5zrqARUiV1xdxLfDtnnu7TkG72SdBdkjTvmV+q/bwJUVFWI2KxfxXhbEnmbn
TjCcUAijZ8ghuSqrcIUa5I4XzQZUOuv+01R8UQNDex5768/Fly6KqDCYj4dSZuNY
VSOiCmd0nlJDnM/Qn9LcfzBcKAcz0oJFS0Abj5iQHo3ssfdvaYT2uMT225z9ttFq
M8ylFDzGcxy070CltkEazjDf2LgirUw86Fe5UHtJNGFV8GApkHNGlqEYSDuCIwH3
wCx1yaKfmuTJYom9dSUv9HAZZ9MwtqGSX4Oqw7ih76f74uazFE4S2sEmGmBqbO4z
O+xzt82i2FqCeET6RpBCdwQPAff78EJlxjfQYxrlU8WuPr6BKaASGJdjuy46XxIL
F3iX80qPfXI4qrsATiZaGKAL5kKgeHrD4DB8bx7YrpXCKUVey4BgtB51qFvTGgzI
joTVk9Qtqs98VEdg7gVhhEUcWxayuAfCh3Ml28mvrkXK+BA14x6UpzfpMWiwuFyT
QUQ1hVRQq1l7NEAHg2NvJ+M8Fh0Hu53UNo5Qs7ZVifQ45fb8TcWUb0Y6oS7tzRXe
UxrI77g9WzJhoc7W7DahoVWhBAamdG4FRsXoijm6vCZv8uefBjqq0pNsd4PIStlc
WU0tWMMH79zSVuf5YLH9Z1TBmVZBHuEfbhRhDvJTjRdy9Lkl2CB8akGimWPljGo0
B3xEzUVAsVGhPP02K3WOccVry4z7dio6FUjpnO1/0mkyYeD3oPxrCygePBZ1xlKq
3MYTI1MI8n1NOoc7XoHGXxy+MFBGmv2HnMLBtFnCENQny5MqiZOaj4phXgu8YqON
eJ8Gj4DIWbmt0sIVKxNDMRGZo2wDTiu3ZGWih7kGWgqvac3CW6iiXsXp66qch7hI
upNzdoqHWqJF12f2SqEhmRpskIembSFLy2x62mLmW9Lg/vogsMsWdqvTpKhzhQGT
VKDwwwTthRcmy0UgTsCKTuKzGEzJrPhjb+n64i2eghqUI89IQzP7+8+RSwm4YAtI
wd1THYDN/H/KyPLTdEjWYdtxmmWTMgN/ldZRVKgBubR8dPe7Ca8Vl4nxb//NLVyn
kpgx2012dmrIVr7nmKwrP80sfNFo1AVE22FcThAsIiOrlrUTIwcM3U/GosDA4RG9
GGImjNN6aJe5x+hNfxrGGQ9d/Xvbkwinhs3UkfBBnDnBepnbaWQOgjyqvWTv+ct5
AEuX3ATlXyzNaoevZD3rFMU/trJNkA79pliKcE4ooTV82+oPBDPpMpdl2z2QXiWG
IZcW4OVIbZIsuvxdMRJg64ke3vSYFf3tVtwXAbyUPxlpkjP8BrxKRlqxzXiChzcn
QEEijkspG8y+71jcBj4bGN0GbOGakDVsEHeyZ2l9vl7aA953R42ir4/LMqm4FOXg
+h45rb/swhrx45LuxMi5VxAi/9X0kuBwy2IHvWPhbiBc1TlzzCw+DshzqJJH+aGH
wye4i3dab5MiL53YGC5340BNau+2oLC/ieKvEY6M3zJRvFeM1htMuy1SpiP4NLmF
eqm2W8g0+7YB6QZU5uQ2q+DjCBUHa7BN9nkSwOlxNYL3CmPtzS3044OPiDsA7KDs
KtuwOeOg3BncIvfNCVPUddTq2WlaHcwjD7GC1UR3KH55zuu4s+/Tq//dgKCI8aaq
gI5fZFc/LBmcs3nmGFCOm4dgmfUDsTQ6SfcKGIhAUA9CzmkNoF4KiG8hb5f1COxq
MXg3rM8xxawHrwdlrtsEatNltM6HKVD1O/BuG0lcejQRYTGGDuj66KvrGR+aArWw
MbM/g0sosEwJym5tm+waEYVRxAmJEMJaIWauMIUBJCTgCIBk6KhtZiWp+U+ejv7I
pBFPvrcOoRmehxaNmxL/yuFJThkFIZ6Xr+JX6IUmMDw6PBPWOl+foKOAB+oxgc29
GPgESp7dazrlNM4g55QVwHpZ3PODWNONUCYOgM2BzbaVQg1/SBDNUmRfy9naS7gr
0Q4BFqi/mU4t8ZdEKozCGfpEBqAgY73jBbpcfSYP8hqx3LSNfunHxVDloEnavR3b
JDYd0qd/DHXyLlTqHdF6kWnTrW9qk8sEXLYr47g+fld0FHf8XkD5p7+xRggTUAXd
lWPdX43c2OE/CJVk+UUZ8XuWBWxcopBDrTwFB4XGT1gFikm4f+IPQ0YFLHZALh0+
g/SKQZnAwlZKzr3HTcV+BXBp1Tf0CP09ltj3MXgd3bvvQ/oIOouos/DCm1pkhrzS
IJsBAIoXOZwEMjgxh40HA9sDjrkQbNBIwO0rrfTQt4AwfVfrLsaMFpgm0KqySRXi
I+MY3oyU1CVvPU7udP9c2HJu1QJQHph4FtuSJuMW/rOZqUSU4A1ihQnvH26Kch/t
ZVyBV7J2/EI+W68BMK3B43hbVn6WTnI5gRCVLY4aetOsurZKMAGeOkapUklqz2Dc
Yg+1/8N2qnGGLDK6kVmXWxlLBov1jtRNA4Y6wHt7mgMsax8R/QuU6RSoWa1czM1h
KO81CZ4eYX5QwadvqyJF5bLRlAVGm4rH/vcIFXpQSko4Ndjeu7l7SsmKSr0pfYx6
Fw/L9AANQna6NnszuobcBgW9x6BUotoUu0GCkSgje5/nvrjdzPYfaYqqNH8ZAOpM
1umZEVyjjhGk+cDfm5mHdyw8sz3Z6WmYuJXNw3ip/P9mnrOXNpHomsNFZh4b2wIy
weLHuStk6gX+m7y1Jlr2XKo9aCbcJpJUF7iKQ4z79XZGOmuw9Nf+QUgqjEcsezuQ
R9t6Ob/DNGCTZX8j94gfBhDvnrdrmA0dyrvITrzpx3xOKeW3fRUzG5MzRYHh56HN
8+gBoVrnJ3rfQAu+bI5rIPhB8+hnh0PpdixbF/Cvqghs1hnzUPDASMQ4FXQsY5IC
5J3DiITP7B2psf0JSqv3mMGUbasbYVxVKUCQSUOCSq9g2o86aYGsnP92WciqssQj
nB5jl2ir5IjrW6rdTWrGnybC6GhPeRdTNu6x7z3WMY9Hz6NBAZKKWHQYpaJOIw+A
lAk97xqEsijqk1kXTNlP/7pN1PbD/Sj9QMHSnJ7SVY/s46b1EwCPGXy8ixtnf8XA
w06OQ1DEIoTJXawoXL7ddUZvOB7s+xIZt4LgGRpTwNDO1lF3CgdCnrQvSdqwQOqi
oRZqjrL1A/rY+3hR/OnI6CEamLKGd6YlPlN14RjoHwVCRE+NO6FyM9mvgn9hxnOB
/iC3qg/ItsZGM8c3kxlHECI1FjjbOg+uvCxcPp2k8VhmIs29CocC1tgIFClkacXM
rOTchRcUXFbNgLtNT258f30sgrHNIHoNd1FhMbf110CeJaGoYnk9ufZ0L9DuHn5A
9y/bfz2ffyiCDJIn9KJTDzU6/9sA0wP7gE0m0aSphAnDyhgK8UMgfqYcBPoc9pif
ZfBJDuxWtJc8hBEmzenGbs/2tanA1Yn2Q3K1IYyzUY46tzjmeq4sEqax2Ul4lu+k
yLC56zq7mnJmdPggXxOTJMhnfgxifM8Jn2IcDT5l0VUJl9PSN+hObAGg7QcywqRC
t7oCdLAAE6DAWjyXh5UxhyzTbAR6LRf6V55qUeG4HQwaHK0Jgon53Rh9+Fg4wRcp
2FYq0UZ0+HFrDUie4n3QRVzQMx60a35lVB6djjTjcPY4iBYPcSdW2lbh2srIbOO6
1JK3t3biJWgnWgugEbz/LQo51Fv9jVTvw7ysRMQH1fp5fjNpju9lyMvf4Cv5oRxk
/6HHeM9oP2fOYj76tqvOxF/DkOxqPE0pAEjJJqdA3GspaViIGZ34HRoE50+uuI+c
qQZQrDP2QV08xKk6Nd2PuPhEIoqZLS0a2upSFGAsJJE+l6mmAhPB47Oxn4+FpdIT
RGgm8YqDjKdtA87a7wLoan1FPFbGmhCEzK2meDahuGTwV90TdLoxUYLBuQZSsQzJ
6zuAbk6azdWr3MjAB+wDjRxMpFEfmxig26mS16eh8rn+Q7v1iXABJrMNhBJeRAa5
YVIYoepoTbcB7uPPFJ1G/Yzi7uewCFZ+hXLv+u+lXLpGqCz54g0xRF7y27m03D7X
BohhBPVj9TJWjOFD3souKWsb+vZ3FwUERHjRX2Pua0t+AIy2ZX5oZWaaDSbF6zXU
pzfkRxV+rz+wFF66OTVUIBKJ3El1s1uhL2W52djrb86F17o72Ov5fB8u72NRw77R
RLA30Ug+Fi1zIpObeXyQG6k3/M6wKfQAQma103kqc0u0uY3nNvy1aB9QndFZDOIw
CKi1Q8aVSbPGA+HsmNGwgojPlA0ceN6jtJNBcM9B41fN3l4WvSngAb2uME1irqRi
oFI5NC2pcIrtZJ0u021hePZdSSj64z0x2sj1Tc3T8+ht+wDXcqj1aK0opqH+AEY2
s0LF7SnX6JsMUvcC8qhPGKb4C1wH2M5sfVa+EZbET7+33LsRhaxuXZ/abJo3DKI7
4+t/3WLefDFj3Ie83B0UG8SLAFU45RzBkLiLYgZCSft+B7rjkXHT8llhLY63Scqo
qIWgtupK0i6kvcq58Tlg6L5WjHiYXCwogElbaRFR5EM8CRTG+O64NMvPYRGLPlZ/
wy96Nip3FF6MdNIvYr740uz2sQc0Wk5XKTKs7Cqfmmpr0v8BTTXE6J7kAtb36bEY
juBLhdXb0vVDJEQYLQAw+1MWFh4Kaz54BHyDIaHz3/HDe6I1Z73UWctI8AE1w+xR
rGNTWhmGfLIS8Im1XmMtilZXl02PfuA6wNpwIsH3RzhkJ2yMZ3vGyEphCGHb5Fo5
TEl6ujYQ0Bj+EVQqdwt/wdRPC71KVyB2KytqySVhok0uTTnJFpdoLdM5K7FwnT9e
quwgUGXbfIxZDU7DDg1t24WpRaTUPMw85i0zR1193pGqMlYYFi/MA6aDa7PlKNtg
PmXiYREf5SeX5JKjxfyVP9d2kxeaDgFhrl8qXUpu/8SmsIzl0I29bCQjQoelyKJF
9rqcbVwStOOVSDMCwIw8fxz69L1atah3fX5buw3Ci66zaxJyGTbqK73O+cIrNt+L
mB6rSC/UKqovFEZuVic/IRfzPFoxtqJ5wMYM7TkqWnrsHp/5BoxcOUV4r41Lju7T
GfSoQLANclCKbIJJF+0vCpuBsYGA+Xs+WsSyPUQEaBcjkIumquDWm9qABz6xC50u
B9p8Rm3frWHBS+jWK6k9aKQXKqMA5/knGEyKb22i84aLH024x+Ft9Fz7puAWZGnC
98iS52oVm53hCVQG8x1xnhGlerWmPKCPFuuMzsuH4ocEdfkI6g2Yxphq/jZe8tHy
EYavG0CGLrpTBuYQ4NQYq62KGEHy84TwRa7zY3yXOznvNf9HYIAZP+16h+4KkBGz
vd0YWMxySPW6AKiJ5RrNQyLX6KsCH38ITbqSmX1eFgkvgSYQ+3yDLA/ixW4EDmj1
rbz1XjAXQsKTQq+zARJkpQlDXcMiN4vMfCHIZHdTudmM4mVyufvxoKpN+uS9rJ22
6F5BEhXYlNP4Sc1I/gloIjytT07FKrf86cNvn7Wh3k2yZ/drOYkyGajXnOjOa8do
h1YczotRbpXdE4MUSEXnwisW16+qCtIt0Mavxcgzb28POhuRozbETUkkybMHOHxA
63gnm/MDCxv6MNOny5VMFj8DN3rCMf4lqpESXtjOb8gHwk1wgGkZmY6J2mivuJjU
Pzccra3T/z/tf3EAGoXYuZxe+oCo0TTRLgGwU1MFZFsJLcwGyGH7bZEsRXVARZD8
YQPP+/pAjueA5jS6zEV7np6ZgI0mZM12jsXEZTcZcaBvg9zF1G+VAHFouTCwFCW0
7/I9bg1dyvQC4JJmM1tWrlfqlMH73yMcmqKLch8VpSuqFgEO8O4kF5JT4DAS9LWO
IxqFM8zMzvrhz46BZRQD301MAQN8I3sW+SwZwUDwYHH8XXMsbMOt0nUHkg0ZfZ4R
47/oPQWtBQeD1bPn9k7LnhKb9bd6jQ6sdCoopsq8OfnZFI0fbrJCf6K1FYwKCEkm
UJUw1AEQhHNRp9sKgZA6hYGca6Xef3PYZ71UxjXS9htRdjvDpFa9hUSB6j98HArZ
5Oc7VZk9iiVHoE4UwFyAJnHhA/epUyLJoobb2UN89jVy9l5OV0IxPAb0wKUnxa6H
W+nbpXM5dT8QG3jbnnb1j6ZdumlEfvMzhzXKSWGfuaZmjpE9IhH30G7tNDlNtuxP
SLrlvRIoUUa33moTAw8u7CigIkWtnO4dCI+CarMLqBdjev7LfyEsb56LxSmNhynP
MIdo9KFzfpTOywe4ectE2ybd5p9ON3IB3I7bcyKNMuZO6xaJJXErxa/TBdk9/D6d
uJ7a3CqxWbO2ibtxn7OWh3j5osQcwANmCNuQGE/W839hdeDlfNl+4HIl43xGeDsd
L3yoH9k2+UPiTLO8CU6aCMp0bD5ypV148G6XvTPHzVzCx17qx3ZfDV7/rzHUneVf
Pch76lSAfP6C32+LjIZ3olJ0fB0q3ORkNoLqCKM1j79Wr4X5x+TdycaUkQJgSH0N
Rd5EjDwzA3OzrmBSCu2FR3mZPAMx6ZCc867bdfb3hIuS15+u4YUhVaAk4e+xAGFY
RBxfAj4kDBURY7+uVXgxHGCSr/FdWB1bi0kIoXyzgpPbj8spXWSGjSns3QZAQz3Y
67Q6IAqzKmU4++SlrrTLcHTq6ZnXG8CoNXcDdh6M5kmoYZmRJlJCvQleH9C3M5hI
4k2EJjjn9cs/72eHfgZ3wY9A6x4k9AGUSSqPZHguB3lG2lKf3HwLgjsDyRdta0kR
CUQJbhM0sWwDqNpJLgXXjr+xtYCfzJ2MTr0QJXDuL4CfhciLn41E2Gpxud5qHC0N
RTi7HfCZj9VZ/47s6CTStzUYHhwZuc9EgpYLfsmXBKxcNMsdMwi/N48CkhmnkeeX
DGdie8w7RonPIgrmHlHwR0Km6SX+dQldhtNsuWyKJMmG3o+3aw2/o+5eH3uCmoGl
SNrAYwWYOXXTLVRkn3lt22tU2XftKwYyFUMwyYyl+RSUGe247vcE2vuP2/Ti9qXy
pzFg6gpWbAntOuy57DD0UsiBRlrIc1Y37ROxXrgRP30FiEuOtlCId7w6wnB8UbCT
OoABZ/m/GqEOpCWn1XCQj93XlBRof/xTdY2KItfALtyA1L4MUdcwPOCMElJ9AcrU
p8Cx7Dbau5C3+FUKQJhyVZF7UgffKSsxcuT0OSNSC9Ab3xDpN/XqI5MyQl5Yycf1
xW7m9LQbkSPRIT6b3ZAVeZfOkUp+X7wvwbcb3ZkOoL/dV5Ad9AOXnmtc0q1Cd6d3
0APyIC9KCnntU09ued+07rB5NEm7oP1L4+XrwM6uriG3chnL/akRFMB+cO1ByMPw
anRq0oy3M8ZZktw+BgJmBWZqS0B+FWxfe/LgX3Ps8FMPvnQGF/aJK7jy+QZ0bPqy
/KOGDdatrcovHYrDPcfuDWcZ3YUBzOxyR7lZ4ELBZzH+MoXpT5p+mahAjETJ2I00
qzHPjwgARkv91Ofg9FDX6kvr8OWrFbrJ+uoejdDrt4+6Z/B441FYgvnnzgqMQLj/
49TvlVOridV3mzD7Tt4bya6ffWpoK0Q/4W+7oGnKqJVisegnKWUAQWZvLHOFGYj+
aQ4uiNh5cXYXoNNnVPC22PAggsl8ci8+b/pjt25i/syN1dtBQLKk90D0FFIsMV1j
La9XWv9HoNW2S4aTRHyoQVZIowl6OZCq5V3cUxh/gKcKtz6WV14868tpjl+UWaQc
u5cGvEiVOg4ok1cR3V1qXh0n2JCVtuPiE0k8pf/ov4yaTgThRCdpWcLQHZKntYCh
vgQjRnL0DFdIuu0aGbr5aoAkbtZao6lAw8O6OQjlfZDJF/PqYzN7NFidUudoMD1h
a0NG5/GybVMXh81XTi3q5R9Yrk+RlbJlnJHlbvad824MLs3vbafDQiWprkEb1C3X
a+QITTqRQo9HNfWDrVQfeWnYUXwLw7vvu3pxI5Uf3qdAczdkPD0tjK8Fcrufkt0r
6Pv2lqtGfww2Br3yFcynI1U0uruONNkqUpH/8/9U/HLwwsVCuwxPelWQaWBt8X/7
QjZntJlJ0l3x51wkhdXkkl+DWFEYk/i3i39eG9ocEupNr5HRsnNOXT2+jG9yXXe4
7ldqpIw+b2n9s/x2GHBcfzE71vlzsG6GL5evS5sYJM5tE3WIp3aQupZYdSLHa4+Z
R1zqmLBp8JyDYarGME1fGgzofUYUwPLFoMNqu2rZSGAkOP8QfQhwL6hHyE8Q0KjC
Azk0G8KbJIzPr2FMOIgMffck29vaHGp/Zb7Gzpq3H0XwpphbHoVM/OWlRRHjD5MN
Ti+zNmIJEz50qBo3kPLEgAWykT5jRsQ7US+1CFRDD7/hmO5YHwwK6ExXAe9OOU/a
YOAHH0OoC07I9SUBalVFRvrjqi9aCrxPaYrnlH6fZ8W6lawmZhYpry81QD5z81SC
FVGFFbCSVSvNxHJlwpJC8dEm0lrR/MeQPhlJEf+Q6PZyAlzN9ItOlPT/Wf4LU12a
grJH9q9sqQUePYgAtA85HzVxST/d7c+djrDELt05K01sJkqda1cBAg51TeSlyWDa
Yninbit0nRjwdwpScLQnZhx4xriqoaD3nAGHH/mQFNFNGIf+VIZJCEAgOkOYC1TJ
wiBt8A9N4DdRFatvIZdpbPohdEN1IsO9XRv2QFMxgnuqyhg0wkq7S6KkQ4SbjOl1
NO5Gzv9hgt0TROcbW7X0NvAIbHhZPqUT06g/IiOjA50vHcIX7uCAM8ctHEAztFxr
dKBe6HNpcKJorQpSad8GK0k/NM6iT7Rkqb5GQWKv1BTFB0g8aM2MCnV+Jp7HMMbh
IcZI5W8oTJRrdTmzGn+5KxBjoz8CvGsbocEN6JVcXcCQle3WZ0u8SlDZo4gl5iKE
Xp+cl8YiW6GTUtzWNhBW9zdXVuKTF492opNlUSY4V1QCgNM2/k5CjkLHkVz8eSIg
UeRR+mBHczRO84X4P9jeHisk28Wl65JwWNuN3TX4C0/QXU08vH+E9Iuc8wmeOPvh
Nj/Y9QvLhZtjJHZSeDU8LZr8UKegcW5ZI2Wz+Mrcd5IX2T2VhKNUTCC6Ixv6TET/
kJFVFMye0qV6LRSiGvPCzMJsV9YynZwA46CpugRIuqGu3dh1NeNWn7crv1A1FGXJ
Ghcuvr4w3MkxP39KrkglrYHJrUgYrmQBtoyGMHkrUw4J24v5vU8NP46lpCT31wSx
0SAjeJ3DQqwjENUFQYcGtm45+GmLNVQT3diCKjbadGUSH6ajih1sdyZ68Ikqqw61
MaQaz4BXS8Ys4hPu1N+15/T4cDPpSG9kcKQ1Fb35DynPpomF1rVfMmSZ1Y0GEs2w
4mjbHnOnnOjGsPA8HBaX7Z6tbUfFk0eXdfZO7UItm3UiBCgokKBRuUEY1Wj5a+Um
SmBgM9rebfnzlmfFz2r6f/AqJ8JruEFXMfRClnJ45aV+n/17GjUkVwWdwGOZVof3
abw4by3Eg9G5NurBla88epfnL3yRy4UQBGVgIJe7ZgNk0DpPzvXrvAnCB1VJviKB
pflLa+4HvnP5KQGUAmb9ngJMoQ0Om+2yXLmwESCTHVJIz8QufpLn+3awwhdmiN9k
C3r4zRRx/KqnvWdFj/Y3ZWY1o90jEwn524M4yh3raJnKtzEOgkrZ4TrjTF1ht5uR
ipWhXTT/xcGTbiyC2t/s6YVWCWL0oWc+F74VqeKG+udB5dakQBuHYVkTzNO14pfG
/2EnElWScQ4K8hSuRXyhlHkUNaSIS/26ujhQFA836QLzlh30pokvW+kIOPWz1Uor
WWrhcvBPCuurTzmOVRD1H4JXMHcqiLx0gQso9z9qd2Ka/v2CDkiiC0jdsfCtstk8
o4A0utiYCozMSESKwzaIEjQGBCQLgoK2OpvbRuj6nBxgV8han0HoC1iRB+iN2uow
otXrcTFgHvM+xCB5Lln5qevNp4xYor1ddLg1MC0m44BzAXzoWcENHgN2Y4VB/xtz
fae49EkUauR5a1lJY55uAhWrOBRbkMMCKmQFJi3cxvSqn3FRUSdpSmXDAImoBDsP
6kolviOqqvziurrsl8wxq3nhVM94w1xq3JUUYboKbsBZ2AUNk8hGJtgygtfILWBD
FNzQ2gVmY+rm1W5i+gkok5vSO1B9oS1z8rYQOtvXxo8CnqJFC8Fv9oSe3ZfYFpDR
iTvKg3bVHlJVinvjnZTLW3XozvE24uQZaYTv6Qr0FUN1KykpscQCZd7bQDft3M6M
bOmytAUoaQp+9tNOOKrzLBM8sZHkHRy/HG3Cd1vppwUPk1We9vAXOFVmN4wPsyi/
GOfof/egcbAl480zd3TglSDgdT159rl7H1p5YX36Ye5dbciLmZqKkM4c8qGIsM4c
VHDuI7sMxLspsSEq7aX7UWv0hsmzls+7VNrdy1XWWJLZkWg9A3XaEzaNE+A3EvZr
xMqtU4Bucx2+x03yaAY8H36tAO/4ILXWY8wzy51gblEHjBdIaq7dQH0AOlAZ9nXO
VwGmxUBvVRUnRiQYSDUNSEv+Ui4mFUSd8qLtQy7u+Lx9cZntD2b78cOoMAk6zAWn
BVbZmwQqOnU+4kL3mwLFULAyocSrojIZLhzemtwCTkm6X6e4AjctQxK8pla/Sxlf
4rU8RljG+9N6cIQY5mzN1z8gnrY1AV36v55jYvUsC2umVBQY6/DkFQEvWPzA9esD
Kmy4iuWSuLTlljtd3BdyPXLUS+xJWGzi66k96fTO4vxgnDukKEmL3CEMdbH4cyx+
jpZKK8okinMT2cF3i4XQz49lfnmJ8GJPhae2L52i22zH5hgVZsQQLPkI7zqKQAlz
41Y9SLh858IsmqNUiCeaOtRnAYUSawecP7Dl264rjlh3vw1/r7L9GL9HHPIqB0Rz
joHTCzBHleIq5y13MZ10jju7KhQyPMzkrLxc5HRzHT36JpAN1VTYDFKbg8ixhwXd
1I9pPB42YsC/VM8GnStlImQt0HEs/nUbm9V9vj8IlXe9X3+H40A9fJXc9BlLm1Y3
xojLYOOZ1HOZ6U/YJKUMcbhp7P9dKK3AOt3/bYe4Eo8Cpx8r0YUzhRL7WAWd+f4d
9Jcl2BIRhDs5loWt41i8qPcHOTbA+6VbpQ3SFDwApQKLeBPxG26XNwogH4Vimpjs
s9TD/hBnWQCOyIgCTHVLnclqzBxYQSMfxcctm0I9HC4BbaD2ExBhPZB+8Zr0RybJ
extMRLIB2x5HVBNPdsdSd19kqbT7nYXdKkG2HneUrA3TrxIVoc93tZZIDlg0lEG6
6eqksxFj/PvMu9gSPIPPOIm3azHjk09Niu+W4fT20rxdxw/HCZHYrFNk38cqagaW
p0+vks7gv4RNXwcfxa+Mgfz1+YGBPgxseZHOQ7bpM3Z8K43iYchPr5FLdsQCc0dA
zMhFWqxWhdk7edGTtB1NnC/O5ttaaoevRnB8R14PxYZosipVXYQPlmb9ITKgDWFq
6hwoUc3dJR8ybgPF171b4dKkjJNs9zjNUgEtkf0OWafJ50c/S7zn1C/71jJ0NApc
QgLlWzLaefQWDAtzjm7lclKvEfo4LYUxa5lnvcZ7qGYwWkjfM2ct487qmswOKDvW
0O9vm6DuvfVd97xBFyVGBJzcu/tj6GpIngPDeM5bw5m10hwzuBxP3o11fauCq3d/
FRsucV8hX4DjdhYtFMuSerCrd62+FkDS6S2YyKCTsXIm5tllGSIm8v9a7NMWEzHp
eH4Acl6GyFBUEXZuNwxKR5/ThsUlhR1VcoPOqDy0naeK0naOG8t7rYTL1w/+cfFI
Ag7G8LaNodv+6xnznRomBeBbDih+9V2C9xPIOFVtu5Ap3vJOyV1mI7jKRBqkDEot
WkI1sniyqzMFLVlZiAwDORlBno6ZpWwyrMXMS4uu9T7NlLriCsvAHV4bVmFPnkiI
TkxBBjo6vNhlng+gpY4/gvusfx5yMQE74JSoew4sB3OF+WEaH7JbDYEadwIhWqWq
mFrmfIMZrcCB6Z/X1sMlprLXNM+ULRkK1JsLmSmUuVrdMFNXRnYMLmL35bHsXYb9
8YgEUIVc2PXy3vg3YWe4Hb0bED1x4jaM3Q/Hkpxscj69gEfU8kdydGRErvbkpyvw
nKZcc3zxsy8NTPaNZqT0aOa9H6s9iZFxLKDgu5TQ8P6mV2yOJ+QTDwqnVRwoFaGj
SE/SuBIpIKIGHPjuxaxIkvyLBfID5/KOqBKgklrZO7TkEM5FqEoWLHJgrpb/pxEE
UQ9+yHmil5CKmpkDgkTG14mSnYvp7zIWE7HMiS49Rrcvgf5MNTMCMpx3IfX3WBOX
WgITXfDPMLjs9ucIMNdvJ/Qqx1dCxyzg1O7uTYGnsvqaXt07X0fHy4yyi6EQhol6
WfIJCLrfZUaBheL5mpWR3R8O4DL3rekx+fj0+nOILTgFvOOKHfeJ+o1aluTHroSF
FzitoeRtQfyEIZXgfZMAfewpUErzsoGVf0feb9VnVzSxZQ5trEl9MvePJ6kjr94W
AI6p35VPrd/rXSNE2RXp0Oy7lGflmQ4VxfLES3UgrCm8dXprsbGyf8fc4Z4BiE1i
2wr1lBQm6QXcynzmb0pWLFXGm/WHqKalzXVT2LTb51/TAeAVWByvDsbnPn5IIrs1
bvZQiKSBw5LSDSVTelTSkr3J4p7DI3NapDeHeIWDggk/i24Hw3Xe48dYYg3Tzh93
w5jY2ML42FwYJHSkY2uv1EqHOzemLqSugpIDBoYOQZEcnxFBsklO5Aiaklf0hUP/
qtTtA+wS9XsE6PRVlc6UUvTIytfVgLe6PeaU70F8crTqKfriBLxLCqN+ddv3tzkA
ng3qPndR3kWRpHPSk7IL4JBO382Ta1nTc8254CRQs4EIhd71+Ko2GCKcSTAT9i8r
8bApVi6X6s90nBu61a5Usf4BO8EENGr41zQb32ZzcASKO3FFUP39dh7JNvIXa8Eq
sI/ngVbD/MrNVIvG8qXKKTXfR8y6ID5L+w1jKvkwrA8afX0SFBGmbbbyqtNfSbo7
hCH4hetNcVH9oC05KRfFZ814Fsl08sxRoW+2vfoGNwqP8f4BOspEHTnyQL56Tuol
MNOGOdzIOOj7UAkDK7FOfMvHLvDQMTN921oetRkY13SaG0tA2/N5G1uGG50+DhJW
+/yl3WdWIWhZQusJL9BQNiBrzj5W0HwO0oiHE8NFVWrMZpCoZ+GmddbxVRaUfqzl
ywbv850bqW2RnVcwArZjRAF+GaaAVJ7bi7UFkj1tveKCU0nIlwDkgdLRMET94uPb
SfRSKj7nsziZiY5DcITuSmteU5SYFcImvP9dM/Tvc34hMMnC7Z8WojM/bjVp1HC3
VisEvLZlA6m8dirEwYKTBXcp1mGAAG6krrlJXyRqXBq2CnX+44CuP2SmUF4WOEbL
MKhloqluPZL87zXC7bDzp4hLIsjtE/FMhvY/0C2EzBCFGNq7yif0qtXjYcZXEfH+
Xv68ffN5oMafFHwsOrPq6zGDCOaMdP9BVz34KIJHQJ0ewmlRkvPyzjUt6w4V/vW/
BD/LN8b2y6xwMG+/JuzBCphjg73BHYcXxe233jYWqDOOFVMd2W+dIL2fijZbbqaP
E/zwXtWS6frAgClWVP7tOPi6sLl0Va/7GPPygYdLOQ+LaxifahwL8Rcchr3McPOS
fLSXZPTnPN0SYZfAm/OPgCuc2k/Ydf3Ca6MwHx1mxKA8NYeTX3WUJyp9E16QjALA
1cQBC1u3BTv9EukGAR/pnsaOsrhCAZNXJ7hT9xYkD/iQyqENg+KOTyCVhkvqaDck
6E7QPlJfazZ+VKWeKwAbN02A3iKaSQgqSvOpYgcji2fVizz01Jo2igk80xCIXrVR
S4F1ad3oEnNyrj6Mi9CvtdG1Px7rAkMaiI+BpwKwxRxBSr47f9OyE+NZ/s952NU9
XKmB0QUmeKtSfRrSbbUFt9y8zT6K78LroGdf28IoixXy4HotHlTMq0Wb0NxzxLYK
Dw4s0kLE8V5JRF5OEZoRv8QRgekQBIrDxcs5NVYsGYWyXojSoOauBqP48O9hNTnq
R1tvzCO2DDxHcQbANKbBYUEsrV26vNu0avhTIy2Mtp5k9nkCM/rfJnp3SHuRQAIo
hxys7cco2wmorCfxCYeCe51sGRr3agAzGKQmYviaYzPpMhkA2YtPAPjz8Ti7n54P
HXC+wPAJTxOaxdvwR/aYetkCtce8JZjtYkCHSDSZYIKjTm9WoI7LTBCeI6PH5FQl
bKYfIPh2D4iTJcsQN04UOcHfTyTCbK8nFITU5vg0lQzeS0Q6Exo7KHTnkT/OVMp4
6/ayuvvS/7srbeAeQA7gXzGTtAXbZJwuos1FuNwLBO/Y/mmKdXY0HSEceNpqUtfj
a6gqR8jRVKAGSgbOkJA7GLCqTCTa8VsYehEkTn5qPfsZYjOkA1VzeB7hX5itTMYZ
nUPDvvdZiIpV0pL2uYuxUd64KaYxnk/Om8JCAxGrpfpg9/LXVwdAt4OCXO31zCxu
v2hjojujeQkMf00ZIpWcpk7gPy61FbyghbDK1eegBmiNp3w7zy6WJN3dKAT9Koop
3/fifVV5fKq6OmvIJYjYIGYJCb4beLPsEzxSWY/UVPnBdUJesZBI8Acg+soqpCnc
bxR1VdhkxsXbY7M8jniHOA2+ZfREFLFa9FgZOVvOGq8xKvgVGMR/qCX4eGY+XaQr
FTyiPO4gVxeBlCnRflLK/IVHHYWZNo0thZQjUbMMwY2rsnlVh3GKf0YWC2KjDoHn
pXVTVahUNYRRtKGmMZtoBL6pB3V3JmTnswbrgkmTxstgkQMX7xj20MFAlZk7n0Uj
q6QTQyx4I1owcev/v/EMKjgMCt+WPWvCXtTIMs4Ei4swYtODOIpiMVEnCwu2H4Vd
QzkaiWA0ia3SGULxNJs+ZJPA/ah6o+R7M0Ni7qh0pe/kWrEBOb30MsiLb06B3xRd
yGHE76rOODR49qPz4uGDIuVfVFzezR7R7WOyMqQwVr210Qhn5sYWJoGTNfpGlnT6
8WqWGcz8tYo/YkDifVp3mp/Up0iCE4RogCFVrKDqzo3L68K0wJf7yo0QiXl8v+cd
tOJ6cjYAFNWbXgYYIpxjvJ9vs8vsqSulVDfzN+IUbvUXjqZIVsLjx5KzGGXm8yaF
ePcMip5r7Q78MoW+TFh6XzZXRh2Y2Wutxv13ve4pcNR/aMIH893uPBxIpd7YTF1G
zemrXLbOcA1jYdJCZKbLJ4zMIY0OTta3pOGj101Lbhkym4yaLKGvniu+CB+QB0QY
LBHSKT14L2Rq2ibITf6RmncZszQNaKLJudWHuILeUpKip5nrmxIg0WImB5c7Nl/L
F7zBatpHsM6PihM9cRm8EtzsaDg+1oJvOOUPpEcjthckusV37o7WIunCu9zvWd+q
ivGeOmRCfxom0Mb522nR+JjmrLwZot+QVMEFRWEyZrsXkUGlASimUDCMlw4u2z0g
QCJAIbGt/VX6MJBwpKxAPWgRWLE4OWiuXhIXkk9Mk3ZzpN3JhxqrNKhaWFKc9XOz
bISljJBgZz00LgPp3i2qeSha/vS6uW/fPvbn+IM+oONG9rCgKORDXozMu13RvXEH
kEyd6yMv94DCQuL7FFrx/d7k1o0phDWuGEwuXoGVobKSQnKKdEv8h4FXVFSUt4A+
D7QJ0mQaS2aVU3Utm5/+1VGRC8w+GEZKPVZ01Yy6uHDm87GO9tvUKYtY+M3nAl7W
uTcabeb+wqON6TfBX7M/zRw8oucIlMKSnC9shX41SDt+yhOn1Op3fpERIEEfyQ7G
q/k/CVN8TSS0++Vf162bcgERPj4g3fobSrPhHHdyTB7atHO4NEtm5oCqZdd/8lEd
wnliyRTN2QzJWQyZDP6idDtpjlMS5KQa/YrluGunOARrzfsR1VAc72IhWqVKmQlW
4j9/VJ4E0tyzJIN4fHcU6FiLrB7N3CujLbXO49hjhuAPH3ESVTrBm9PRalk1owhX
9dS7ODXetjmmj3MginYnl9Nfb9k/Bh6RBIgAH413fMhwYG1U+3eudFPKzEjUq8YR
7xr3JToBvQAJrjLsAxJcEfKlXFcYbgRlhfioBOTAOUibha5Z4oEbQ+gK87DDN5oT
fCIMztRlvOPo1AoXAkI4iIVuhYamE/nncxLRBxTaIQao/MUyUoB0fhOU+Ow/D3wG
+hYzpYvqYIz7A6eDs5baHwwP0h3ySJE+C5Rgy8/msjkrnFofuXB46SqFuWv3zhDK
xtk0LEy3otmFxvg5iE69cD1WXUEv+nRsi3BH46CTI09mnNIIcObaxvsdyypWUwiQ
5vaIuUJSelLoGQRmfBFnue83oIed6BspEY21wCCyLCsrz+AFQD/Qs4xSVn8FVsP+
fh3JPzbbk5F5LQWikw6jw8DXbNcFA5+UOu0vBgPvVT5Ku6LooKAM33v2LLfyhPXq
PNVlVLVI5P0ZYhVLL+hEADZ26Acby/p9dVK/zoouhsntS8XhvtsdrUIaMwF1oH8F
AQ4B7DymOfHuH1afEC1+a5by5d4c2ReNp6yQkzupiEF70v86BDcCBenEIXZzuaii
LJV7UknfL6bvmo30aD6Kv6ZhaBHvrBDLgULb9lQm+JJIOBjoN2gSGQHOlbzVIk2k
Ezz9gvLD3U8b91q6Te4RaW+k5/qXvz9VWSwSqgBwnkJf8o3QThsUV2H+aS+upI1y
79P4UHVxsV2/khBLqTI6+sC8hkw2ZlPL3gNsgOXcVCsWlIgboLTltIypS6XrYSwD
+Kba8slLsv+CBAMiMuXF3n7inryhi5t3wQ1ptnIaUIv0w79ubLJhty40yHCQK0ad
Ljs8sesIv87H+wkfoa+m1TaKl1S/d1Se1A5/BGHW4CEE7gTzHb3ADXy/NZ7h6bqQ
J886Z9FefajRWyGhazVaLk71Z5TE640FrOO0x3WS9I+aEFU6F9cjBkMdvGhBHX8k
8bFLYT/FhjqWArCt+bxErCxJxMYr8x5WDfgc5F3NDCvZqtmf1Zfb0CI0hEfUP8me
YE1XiW5GL7gai7AqH/xZJUUR61/9tHRvvKkWJJ96mNWjsIwOgbSipCO2m9gVLzrT
tWA3tG9dcdz0dBduLkx/AeZq+eLtee4jAkHPg3nvvYWw23u35IjiIhqvLdyVWfe+
Y6xNmbZPHLMi8GuaTSqWGPWYkIzvthG3bZnkx2Pc2TZcNF1DDyxqAZDUWWzn25Lu
PSGyJNJqQvLPWRxb4/GH5yduJixUZMtFbJPq9K0MsIqNSbdKtl1B+FJVK9+C8w9L
CvPeTULHwKcxXtq/xjTteGZlCIxb8+EMezAH8uJbS+DbStXnN1IZo0taBFrKGtqV
GLUqGUvSHqD3DigmqM+SggfAMbTKkpui1DlKXyGcbfsUWWEFJ1PXmYgHh2VY7z0Q
RiJ5R2ODtTOxjRuAgEO0F0xv4Av1nODr8L4gdphIkcP7Z3uNlahO+Tmpku3URmMQ
X90qXP/+UBy5DhZ76LlvTXdBdO5G92GqFVndAIhHx8e0cpO0kEVUKCBfpm0mgYcK
BBnnmgn/QX0vLjNO1bop5UfGc/Yyn71C/+wbixkSsaltKZqOZJoISPsp9yIe7lqs
dRsGUneBu+PtbNVO/w48GqvnfOxRZh8R2/re1Fxj8LGubqcDdKOBisoBRVIZpzP5
fnKqADPa8jRySeh6tX63HxKH2G1QTseirW6bzd0ORdBCykG312LbmU5KFonIYJJr
OOHnT661eXRmXOJVRYLy58ocOmBEqRqgUwO3BA++z5C9wjyUkXTvmieADPUICrpb
pRrydbO3L1tdOiveJxbqbr8vmnIE0JI+3E6EzP9OK3KUVd8GtIGuC0rV3pkU6jdA
6vP4ulLsinOxovGZYyJWHNRCPIULcjazuRKxEiXXJQT5GOfcIfbit7BgYq3p0w2u
gv8uZJaqHfZ+Mf3qUL5Z0fgNYfn6Yz8Ez8Xl6mDqGa9OY5ARt5mBWK2JHTZC+8wI
/LFOcz9iXg5H3uw9h3FPh0J0vTEd3Kc5D85oowHsVqAK7jpOSegLvmjnSAO1zvJP
uJxJGPYo4k8mSC/Ed5oKMCRBuO98Tm6+kdCNwkLRYYr69XbEq3HcQl495vEpPvdM
fkM9RPSh6rDxThfW0wn0xbrXN4ojeur4scoJAjsvLmJAFg4GnXrE+CJslWSnOdN0
I4GS4MntbRE+mJnyZIUS1eb/ObkfCDVHdPi1NmS0ThzRRdn4wXhvm824la5zyBuA
J7bBQDqSD33bvkLsZw1ZY2WcKwKyCYH4bE9PyD3tEgMWhPd4HpSCY7Rhb4JHJGtQ
Gii6WxOftWVKJNOuRFzSwkb5BxDKsGV7EgN9XO1GDPK/F4v8jmQAkfUVVic75HVs
en+Gk/vaPEcRVjcw2i73lgLnIb0GqZ4/aEmgAHotVLvc+01WXUGfkok9l1xdPCP1
PAe66DKg077ObXqygfEX6EsP8IIt1+oLcz9/aZ1TaWNtHCLSpDZxdyavA+d45ySr
LA7wMIuM0uUzY+BkqfGMisJiNJJkuF0BHhxlR42WXrBEW310P/K1KOBUA7/d2IBe
+UM8MMivIzWr0904dm1zyvl8DwxAEXXHubA5+nbWtDFY0GZM8CO6wH8NoypLDiom
3oHpfgymBBbOkznhdsdl5v/ZwVjaD/DN/u3VFnPgWrQJyEsJ4ByEXXKYBBmx8u/Q
Dg4vdLuSypZ+fRMAmZBc+FA2Ec3kbzBCPmbojkjBBb7nabrqSTu+ppuT6/eJyIlf
lQVyUxK7K6yoHaZuRr/SCOmgGv2R61ckZ2wAj46WPqrYQSLiqvRl8dA8y+Gvp/P2
ULnjrrjDVIk3p6AuTSLFEeL35ehgIEAxgog/LD8sptt2TGCSTvQoZ8rqWW83Vk0G
HhLFvfvKe2W7DfJ1+OXxWTC928Y9l5UboYHS3BOIJ1Nl4IHOOQGIfgutw0RSIdeK
5eBdAQLNL9hNqwhFwuxNLm+jP60j3d8VvP2+6ftgH2J8cshzoWLWy4FQdwaX/PFO
9GN7jvBnWJPYcT5tAu2Z6OrPCP+LgQi99renkVYYhs9f7VM/utX/PnwSP8G7qOho
KILakfn1sqlYaneyC4tLbZ3CXRM09kCqRdvrk0DiSKvBGvOaVK1+Pzh/NUPeP8KK
C0Plf5NYHVjOJGTeGFNyIQP9apbde8v80WuP2LzkbpftpuooRUFbvxCJdtxR3QHV
OM40yop3om48k17wJMms7Y6EoO5dIHORhgSpJjA6HBOC04HL5E5qQdEB1FnSfuP5
Dompn+Z3ym+WaVrBXJhjtGUMOpKNP8255u/8gRNVOW7hxrQAhG8P9gyYunb6+s9j
gW1tqfEChVfc0XYkWOH0Jlza5KHojyv/pp1r0U38Gwco2LGjT8q62CPqpJ7jm/3X
/W72/2cIp0SI05W/D/aabCWDrjbKMjTY3gVJthJ9TVxAZawVTkXV74oXGlvJkvMR
VIeaCQY9fMW05REs/xK+P3TyPWp3gPnfLpI+32UcoykQPJM8nUJu5aDByK4LId84
gOVdeYoGCdnInSmduklROrrME6dxK1w+S4e8WkbxZ+EU3/3Yw5XhqlgDZIY6S58t
hMcduRUap+BxokZQ6glooOMK/CoX32Upttbv7f/UukdW4LMv5LMXLLV2azcNa8zG
cRqVAir66JGr8C2uQkTFFXOVkumYMo4z5st1M+2LSwE/9lkj8DxUx+9fGfJPZbhG
wGTVekrVNebHP1/MbD1ZIwvaDmjE8CiMrAQis4e8leYo/PL8ZgQ5Bn07/AOIo0rl
eS8vrM5ccktGJQN/HW8Ot5vMg9hM+8U71CCoFmEgMlAjqITydhRVeeZeFII8oa2k
SwA5RMoGDwBVfeJSwIAzfg+lWCt7nzihBbojy0LEAHGyhK3fjwfxW4Uavf4POCYG
EjHDtNcybMTs5pmIYn/pdL5V+DtmmwwnUQ+VZxQNsNaWOSYOkkRWv6ksgEjKqVBu
3gb0scraH7WAF1+vhp2cfzdLRG1wlDAmwLuEHQeLGSP2pf1l1ORp9hoT8THOAL84
xKeBhHpNQJwiHh6b2Q/A1aYIIsWjMZL7eJxg/4MwRoWyVmA75fX+BcmzD3rNjeAT
njvAz5/T524Hg6lJLbzx6i8OSu+RU7xOqLCEotEB/NgHNNKhWaaCenjWsRHovDqE
nLxKK1+4flIGX2BFEe2YDTzovHrnyOrd2VXa73PUCUkKSJdp1R2hpx607iLiy67Y
p54I3P8/YXtRhTci80g3oJO0xWMLh6UmAcJaxXW3EN3tvjxUhh5DodmTnBneRjVv
o4nDZTRkaMZsM8V4RpG+Y8OVevSbw6hyRMnEJ5fPLRnyUDEu0gZmkscHWIA0vLzp
YTt9O2cWb1gsK0OyipAvukNCJkXsdLI3cKMcoPfct1JMmSBHnkAZ7cKWJfl//e0m
YQRp7jWo3QBeA3MGafCqczEoQvnApH/WGngUXv5Ttcb24m6+Eb7MNAWyyYskspbx
igi46m+lqDqVVAs5vFWIYYp1h4ApV80olNzXe48HXzDfIoG/yn3k/TLNIYZkCmUU
Qv9maMqb3S82++JcHEVNiVOrMsPklv+ide+6WwThdTvulPpHWUY6Y9cOnRwnIhwh
fn8bxqLsqI8Qp1Xrs3Fdgm02Eqs7QgulyBbkYQbfqqWNYnRixAfPeEMh2B9JwnPL
A1R0XZA0QcXW9I70NH6zVuli6x3GhBMehww+wOFtuaosqUHRAvjTFqzRY3ZfxyX6
Yh/obk+oiFnx+54dvcO6qWpk8pjYNE3HGCW4qaPoOTL5zm3CMrylcvArbyZMkUBY
NGAttLFhmmHIF6w6O9IINTECbDPUAwnXPzDVW9SbegJjVI/rqDbt/wxnEecJCuHJ
CImaTQtM0EGBbRQ7d6InZLbqSEcycsClTOUr4Zl+7Ed+cTb/uvWKkiRodOdNonku
H10zIcpeOV07W6naURJCXJlEpHQTmI4jDDL3zfavsCqIhHkMK+5xDHa6HoVW8gDP
3bfUzA7i1S9Q1HspGe7V+AzMZCklB5JBWCSn0+NTBd6o9KwJun9I9ABtH817BagB
ydDC9/r30obcmYYlbf1FeMYqy7hoDiuNRgl4m25zIEyb2kpDax5ZvWCuQDXjqsgW
VjgGwNBk60aWRa2sPuDCXOM2ftioIo+hFQut5GxUE28LFWfDtip1zhn3v6umSj9I
WJdijHfBeQQL1OrfDbyKUFnJ7b5gD57tvu3h/ghRGXfHXQB85E2PoPK18z/JwAiK
Ht1DgdlD3C9NxQND5o0KONYVX2xjhxxkq+aWgl/ACns1UEz0d7mZd+ACfrp3vvLO
NAx6/tdSbM+6rebRleBkkirqFPi1r2m+cHducA590guY4E415RbCf6zEjCEuKhoT
kr5vXvUwAg6sNYlN+WT+faZvLyo2v7GE7YlKKYqz0z3b/aTV4cMqtEHTPXH3ylXd
cOtDvEOkr9/iZzc5laojNP+yR4+dOfYhnwGL2JRbuRvHwCB7cSzty851FmH+kOA2
6p4pNt7DhvsL8nN9w/JRM/fAz8hj4qAFfwGS10fLe3ALF10PO8XT+PK5/wrKwj+l
144Ybhjj9/lkdcz4A7uYt6MHanFU6bbqyJ23zwSOLe88GtXg4iT/oK7EsQbZKFJ0
UiJJDaiwfLjd9AhyTA4vBLAsdjB4qzoX71SMRX5lSpH9Inrz5yJ2D2yB8iyKOT/d
UexXQGBpT8dUHv56jJeGHG7gDmPDasH45D8Wx6XXT7tQBL5uQhrIhdxArzy14+Dz
b/Z6xz4fanVJObX1BZ0ot3FRFcEztt6lwBxYA9PNkbLZ6CV10ekf/OO++Nkd8PtY
JIZsC6teeZx9/lSxHm//m1A+8gkxceZgUr5M8itsEorppRCsNT4bbTwFyGGNVsTn
EOkx8AlRABSm8PR1XrkRaKOEd5ShDWwuZ4br3qC5sfiks6ARqmj9FzhJ9SBY/d2Y
5P9bQ1DSbVCkTbYmrKanShrdLum3xoDh8p63kcetuTJL+0XJHzXAgD7q4WaVbAMf
aWzB3MTIkaWhNRTCICy/3/NHwDbEoZO+ZJqaszLuwcc4kuXf9KLPaEnC2S1IbiNa
bGznrDSwfgfE9/pTK0obB4nFkqU26E7YiXg4M+WadLf96lp3W8D7Q6VhswEDfWtg
iep8675evYf167WodgNGVoJkp90zozsuIyvwceLM1kGPGnfgR4tSr6AViekvEhcZ
CIhkE8gfAKvio3T2jpMpFNdlQsfxrTCsBTc1zRKy9mLpNH8R3B9fND4SYMFEC+6A
eaq4JsSRNIwcVVWmga0fIXfYZZXJ1frjYLT+clM1Pg7jQ9xWMbCCPiMVpzxhhiTe
uzMLjeDPq5sqQGmggUI9xwlyraka/S5p4CKiI8Z6uVVGmfCOmU5Xi4J3icbpjTmc
k3Fayl1G1Tphv64lglo0nhdAw3tzdT1j24GWauNSkR9UIuao6CLLpouYizMn7rAL
aKODGOyaN98UrvMX4AzwFmr4IzcoWj8YdGvOtu/H0Rx2bPD4VUAd/61PIiyFHwcz
0anv2LqMBhCgPAczzICrh2HXIOUq7BhHofXN/+ZwEqURlQjUb8aoucvcVaujyvBm
oMs1uWr3jG/tFbdhTJ2lMD3rz5o8gG6VLCze+dhbBexyZPC6aw5mqFFHxiegU8Um
8AKa0pckWOEbnRugHUydPw2IN1f+Rwa4Od2z41izmuNDpxjp8gc5DR+Cxf8tr2wD
AHVo7EPJ24xy4zgw3UG5bRRMFkdRjomy+G3EH7CEWNDcQ53xVIkOmFEKKbJB7u42
Xe3ip2Xa1pcgFaMs8banvt96+CCgvwa3pMJscdQ9pgLBocVfDOJEM+hZ9+Lg6Ugr
sX6BBSS1GYyWcaJ6AMC5l5N2DDkRU/HVlfOq/3n/KNJrzZamcR2U2UnFdOhGZyP5
yCxfjkAQQdqdx/S7HMHPDyvaM1C/5j3cKP9j6U6i9nTQjKkDXotjQo3YOAbEFqCy
xhgMNH4or1NrBMv1at4oUiCQ8Yj6P6nGTWl+CAP2dfHctIxqEaAk2llP5ZUvdRvD
RFYlSbpNfOU/6KxDm+lhwNfY/QByUTmapiE8gqYszYDerDaUDcq5msRfGxxpee6a
A4zaaldZd+PdG4gVy6yWljsCK92PBsWlsVa3W5n8TjBvMoIwd23zY3dN2eFPQBHZ
9KnHO6miFDSNrOGTgzm5GvwLwcNhqfRo95yYgpTDO1lAY6WKzJbCLZCFUdEaDYRW
ClLjYjQxpgqlkQROAEXFjYOkrxPoxjVqOwiadZaiNpd38VwPHKdFxEohuMwJvqsU
4ObIYrszsR5Mdz3VkZHKdutK11v/oQpRX4szRLWhCmfASvqGVzCNrYLrJUh50Z8E
jrhec1qVhqFFlbUJbE8/C5JWFTiwvpB7BFUqmlRgTBIQdi0IFQr0BwZjyDvlsI2e
smG4YEuoC4Q9wzbY7iPdNThKp0Uwz/WPN8ooJz5liOWO4LrYUEvtKtFwpVpbi/FR
XEyFWeljo2z9fTL2N/tUTY/CMedshFt1lfcw6Y7u+TL8zUAjFEa6Enna28w40Wl6
N16otXGzkpgIPgJCxwiNKhsGNpCIudHeQYcKnPqAafgFfheJWLpgOd+noDpVVpsh
GQ0ggTvEFPZOp1tVKCahFs06Z3KVkXltpv3ryMfboqGYn8R3YRpVyjmRgdl9VEQk
kCx75umjVltc43ca7x6dCTryhW7EnOmc3JBLMCrHGMJjaiJXZfIlEwyxgCy741/z
5NkZM/QnKZjRfxN1OsMmEDZ7RAIS3nSTcvpuNbEcFIVDym5ZUoaki5JWJgyZPv4F
sMZUrmuv8KQvkoTuBNu+ulwPyr4HiU8S8yDm84lTDiIJsy5+id6yBiLOHdIBrPHc
MiG2RgwEa0mP3DJR4EvSqN31hAY+2WmOJv6ovRCYM1qZz1UrxHTQSi3IChzdlqsY
rCqLfvkTisxuqhW9Jh7dyBov7lp0OGvNsZM2PEywZgulHb0jVlmkXA7kinYdxQLX
aZFEIxy6NKMO3vZRxFEma+8ioR+pnEKYGrAhIetYvTrbCGD3dKeJKj3DKc41gbEN
YXXCjyaFvPnJhq/1JJLLIbdPHpdvAfPuaq1ulDeeuBfnDS7xqejRLjy0MBB7+IZz
M+LryCS/hFsQIJZw22p+t70yuEsZBnPpxH1jmhJbo2WEqojS4c8EGutqiamzsuDF
CyuJ9OG0zgpyPHuntkSfE/I1hk4N8KSdou+tduAz+jewpYDhz/whoc0pl3LlwY1M
ZwlMoHBdPbVxxfdV6PmFv1Lei9TB/yODR2TbgAqfMBthfY0o3gN3JyjVqo55BnEJ
L9rNHcreSgrJZ8HSy2frWWj4s3S3QpaR3iappMKc7z1v3l3itqEzd0QUvS333zqB
yilnV5K8SU741fVeeEcIdYjU+TSfmHlDXzInV73e27QJoT1br/hK+8aWE0/2qPsN
2qXmG7JS4vmW0hIewppgRb0WdDwU8acZnEEGujGa2wkEII95RZTrO8ED1Gxuksh1
kFRaa+WSDXEhMcTbv1TBl9k/enptPrnikmEumyKLHlQUkxhfDlNxQajylXDE22/6
udhzlMt5bJAzNiC/Fcbz+XnIg+pNgMJvUDF6UX2B37k8vkQYpEwEGSuChhKtRYPQ
Rrxi6u6k9fout/xxIU/foii+L3Jm48KbBPurToS7584iyp9q02ZCZ7tGqzffQmGe
5c5uR/YVi0P/8BAUDBXBCyGguwwYCxqIsucGALzhAeiXhtTknibuR7Koj7FXBhk9
KSssCeUBXJYNp1oyC05fXSMG1tCK/5cAV9qTNTjdvAOufWZoWIPdZv4FymjR15Bo
xc9lCg66/Aal1O2O8tq8UG2aHqTQ04bp4epmuIWBJOkn0rCHRimvEBIfFoZRKqtZ
GeZ7Q9lv6fRQO9ufHcTEcWnLGfzlc4WfUzdDc8/fi8l2N4BOKZua1bHI2F8bUMel
wDdgePPGMG8KaRagtO2308QdY4PGz408xMHCDwV+gRR0dvgvY1f7ZbvcuS8Fm8rr
Io11qJuuoqoqVz3NWWA4S/7XCG9BnnqLV/m1HLSfxshAf89gHNY+LKLW9MHdGaZo
2uzuBhEUp8xetblsBxrEqC3EKgKehxL/NTP4dZlmjAK8YXXthn2Iushdc28YsxDj
+cVxXqphNLhqCsdT8/tmOr+CNsLEoHn8VTvRBC24ffxwdH2V3OMhdoJRmAGUJieK
ByXRMA14ZMAclZnyMgf8Y6ljBUofDZG5yD/lMasa5U9OJa3vUKXYZRPVQ+5cV5zF
azYu17U/ZRmMAtu4OVNq3RguRL+Yfg/woyVemufAL0Tmca5W26ifjtORz6qJd0+h
WdpKFVDclcrUk0ht1l9CV98qosXBGtJV3cB27uRDIlc41I9g53VeF/ka3VsDwk3G
SX2usivmN54NXwTJzQAOsEcNjdCgr7PIXdjzmVdj6H/MY0BH2Gjk6AhoEESmy4uS
Jy9kw35Oxj8ztLO5b3enc0ESGiU88oiOnA5ch1oM3beNvD4VNX5WVqqssVopZ6m5
h2r5SR8WUY6LFThzXHhZRngvXcLoROupXsAMBK14itbrQUYqYTEiA2lrdMmLnDJx
j5DzIfNRh4c+pulTZhQS0NQud/ZCu9MMKXDGA5e02jsNWK6MmaahjugDgwmb7mGY
YJwDqLG/DNl/wmhh0lZiEddWu9Yo3Hudh8ppnM2u1u5/7vz8zIFVWCCzgZcauFmj
AJXAtAYgBAy0IhZQt7vNC98c2tEOfpvkbMVmPViesQvGofK5jD/91g7vzFVtHvvR
MeRf/XIXInsCuIiiOBWTN6Z2r7zoKrEI4gwKkQP31gl2TebnqJPcV4/IG8IjlyaS
62I4ct3HMJ9Z6ILcIVQlUt1tocCU1Es/G5o1Xvyb6MKqZ0Picsovvilg2KxPAJbL
1sJRZ1ZMn1UTdtvIAOgDo19P0BVC4tqLeWZUuI33xO6v3e0c+Ymfi3CL9jTfgmev
olmj38iA31YIWZAp8e2b1V1YeeaEMQwayGJEHpbyvgdLO7taWAItroPinRV9SSkN
SeJZYH2+StT4yTY0hYv5Jk4g1XkD7FLn65wIXf5syp1QMLTWET4CdK4XVr/Xc1El
I0JFLGG1O0meNG8Fot9KMTBDk3UB57LRQKgL63sblxtNCOu5kHS6w0JlVYyn0a0j
tkzN3XW6HDNv1C2HTNDkZA1nlUECRgAck5xJpcKLsZ+oV4bnz0pPAucRMFtsDcCJ
MAWsQaBuIXuwgUxkaY2XsLmspQkrkmhkSW2jluFYtDHPDbIf43nsWN/+vcc0WZJe
LdrvLuu8q8JmnbWqyOxjbZh0XaGli1lvSnIxxYQdwniOZccQQnAtU/A2cgmsQZpZ
LEY7f43IhkrMAsd7JL8qEBJmpNytBIy9skzwZ86uOuzvFiOgtAobDPkTfYHEwOJw
pkERtBWdUX8M/mzpaHnzuZaDqpKN5wW3q+Kylhhigbhfk/nut+VDZP+GXNDx+/4P
Q/PgHUjki9w8ZPkE3JZYecwDx2V7R7knEFi6pcVuTOwpB6CSjW3AUZf4zj1I3rMb
qp6oTznhRG0pOZ/q1RZ1J6hHlSfHM9hqgXuKdYrS56HMntG0e0DSyqs6L6gkC7SF
IClSt7nRLgrJHyuF3zjh04p85hg5q4ZBcG0tG2B6djIJbXfWT761n+tgbvUwVsBe
XsUnmCfuR+bXweaTd/9xoDKc81lzUbyzVHj00JJEtglb/zEyt8O6LMN+DO20V286
TjO9UCzrJTf4L4fZImyuXlQQSfuys4fVINdSAxE93c5Yrli9aA7d+nVfDAhD3mxW
IGIB+2WFiDq/c8AMlao5chTdvoGhApmJeU3/H27zTtyq0IPoUSwvJPoaFNI37Ebp
t3gtBmhnejOF4fMBxXWHjYFjaNvGC7SSbmp89VyZNMt80DjrX3zCPcVav89Z+UwB
46sXeXrN9tUSFKsZ+kZ21ChE6hn+1EVwQBIFve4icE1M3JbIfZyRmIvLK6t7ItOb
pYGJux4p7eYSykgczqgVVmO4yErQiaCRtHOYi52zE2otIFhG4xjMzyJxZMn+9aaw
N+uCwrwDFL5bQI7OViFvC4jsa63zvAaAy1xuJ8+i5cbV4klqo74JBcKrL2AXsAYE
MBX9tbBOC+AMggsOXYE+utJV+qiBw2hPHSEkywY8rNAMQjKowSLK3hFvXGzKgTAi
bAUJNGhIc5Ybp341HZ0z6bFxoUFM1KczMe4Prckwg3QUwJJsULCzDpMSdOha2pXU
6kiYCAKEIeyC03UqOoc2sAc7huXtu8waS6CTuhLCb5SN/7+R+avaRWT5XAcBZW1+
v/xoqzizUyNwPXXbob5EGVqQx3tb7XD5eMsl5XnSWMIZIOjuPGEg0nXIfS7cYCy/
ZzzC7rjfyraaJbD/VzAHfN+xkkUCHoadEA7Ze2oqPhUvOK9MZW4CVj0mleEWRx4l
mAIYJ/+ty6uAPXl87aWlcIlJVh9LFs/5qtXQs2Nxoz2mVLVnpBa8whejhy1L4iTC
a7Sxr2ZXiBjOjXWdsBR4z9pDt7JjY9byOPMH0fs0Z52q+4W+u306r1gEvx3AyNVp
Jlvz9ncW/zltc9mwKc6VHcwKjkJWPAd93NzF0g9g58//CJhYEpuZJGlc6TXwYoY0
3MZwcP5+1tb5L3vUq+jeMdWc3yuEUOdbcdnkH2WMdXbELb55UZPtDBQz0Zr03u8t
m+iNt75nL8Gx9r80dyKcOe8tdLQWxVjX0uzCSe/7UziINq9PpnEZuLSZNxoDW4p0
/O22qw2eLflAtc8MbV9J7/vzpJyZ4c8Z+7GfJAeemyplUqRPOd7B9z6gdzqieNLF
fjNQhd+LrFvGy0KAAkMsCDwUXMMco+a3NCl5EOzNb57WyvJcd0RxRWcOi1Zlu+Fu
b9KS6J0ty4Ni3ikV0keF4x3KmQmRWQlWzgQP+0i3V31wITnx2NfvwOXsp+YY26pE
WK8HfszuyUm56ouiDH3nSoRHplJNf3jti4grJ5u8Smmb3EZ7ktgOQ5eIzXo7S/0/
N4ALcxWn760jDaMHfniDe64MF6eXORq34KhmHXglZf+vq3xEiFjahmhOb+ss5hiZ
s9FMqSxulhaGEW2meDqniMPsDvptEQc05a/cNlG+MHGZyBzTvgfrzp6hgPEgqY0H
5uBPjPGsdk+O4U2RcsRqSqpMJ76OxSJfWx/x5Rj+a3YHbykwb2ygfwRiNsBuMFs9
P013kPIxh/c353IO9yKOMLiRYgFJIS7XuyXgJk0GrnLZ/Jf3XVv21lODIEYBxkZh
2IpTJSAbYsSsoG12Hc5omtTWP7kvx/Z+/NsFRLxO7LrmKHUswro68mQapDIkRuUA
aQc8vrppb1z96c9Ts26jOq/wKcfrjU6c51a0/TENgoUzJzpi5prhZavcBtkbNbm6
yYY9Rwj9oQ63cxq7GXlo6w+hf8Q+KkTMPgNeZ9Q5AmGx6IY68Zgzx0AzjrF7psGY
v//1tC4+X9uCjDW3JeIhTYs9HVd+hz/DN6fo6OYWP8hZinbCigD+LPlF+OhTWLIU
985ldWY3iSU5pSNOU5s0JAZIaAriK6Y9X1LJqWadcGJdNEOJdpR10w7KTiwbw4qi
zvRd7mEdYG39kOeX/PfOpC8CZL6Yfc3jI0zOxiTH2qVdLQa/G+oyd1U9MtzVwjFP
tDCIyr6+BNtdVYNTG2D1UV3ghMDAg4mx+9KQpYq6mjSaay3q6vqMTRbLR8eL0NGl
LrptxGD2IHWRqcw/29lL6qyJCUzDhu3ZaLbyS76m3B8OcXRdVNQwtEiNqlSsFPRG
XXWUUxdS17+DNbLXgJ1DHBSKKnkOofcJUqXcIU2Hqkmpqyp87T1EAKffaDKyTgsB
LlBaRiG2QABGFZa1z9ER0hIfJ5e3s8/Yv9YgNZkHihZSgWnjlO5B7z39xKDwizEO
br1UaG8XqH417sL/h0GqmHuSWPl1UqTLKA81AdqCgyUeu3cb2XMcb2ibG+B2K5+F
5xv3iDvwSh/CS6Fyh6nLMaoCG/MYqDY4RJn9Q1VAezTXfaVaxrWslpbBCQ1Li19j
OtrCXNEzePTFPc9/nzCUbNbq2fHaoWpBk9Gaw0tBdKz6Lf84voL7Z7isGL/YoI2F
W+IXovT3ZkE47mFE7xsf2pmk5nO4wl6CFHurTZMj+1ZUmGKxy0GjHL9yZu6qNbBR
f3VK22WmPP8Ez0J88Du+hL3NInhwEVmFlEdK9Evc0M5EIQWtJLJsW5vOUDFXkmY8
bjTG+WotjYyPr3NTZG0VennzYVUBqi+AUYfiO4fqb0xwUS7K8Cf1uxNNtfzj311+
k84vI9j9ZlA7eTkOOYCOxJ1M4yTnAoD0ViU0309R+/ZvVya4slTlsHY2pGfYLYlf
ab3rvrI8AN5b9jR9cdLJ0v1n1H/38yJTb0KvUEb4KlLOsDP1sx7iyUkUztsaFCjU
rklsJN9jpJQEzvVQTFPO+g1rDKM/QzuVzHOMwXT5KDDbNMyTh2WJqci/u3ueLHO2
NLIUSaOYnoqAI2gV69PFxm4QyWYyYajQyNkjx3V6Y2qKob+B0PWMxJ1ME0RBusCC
F9qx4y2zmeGSTVGHuMX7OAbVBim+mZo5RoHDYBr//3rbd3bS/re7vkpdnO/hosIw
lJ1kSPf1CC4lNIAlFCa+10vApIxsuAsjoVHlboTufv60YqVlz1sf6OJRzk9f+d8B
FIqHc4y5jocEVqEwiZbEZPByVe8P8Ic0erRwZcUN+oPPw9wp3iy1aQHlF+1HCUPW
RoxpO9IQ9DDK3QmektK+VV+ADHA/7bbcQL3epGQe1XEACnXmmlKKPcf6HvajoQmi
dX0Qn8OBG4+2zORFfbNQ/v8/CfahH7dm/oWk3kfH/n+RYeW67HQDmfGG5uDl51CX
A/VRnI/VvV9nlRr3+T7pCkxZZNUEoXizpx4R7TZYByzfGA7c+wZexY1OfpwgHciP
ca3JmUz/XBvMUVTj16H1MUo5iyGAx45mt8Ybahprj5CEU9pmOcqdRBYZZ8nI/i/d
eYGRRaojfExnkfgjstAHnduVm9FgMwIOddZDjHDnC2QzbNox9Uu0Xtuay+zbHgXR
elgjJXYuXJ7THDsYDKvGpsWIGdNJ511k0ue785Mu4nVrp2gKihWye770hpNXJr5u
45lHX9nhGaa2pFAUYpwh6m4cVDoMbVtzQ15XfKEJ5YPQku/w9gqbCpipddiJmAuU
GjuWAJBhhqgCDE5k1eedPmIMlCmnmlaSS6NtprO5Jn5P/OSdWU7QxnvzwnfLwcE/
kbBawgKd3jaizGvJ3znobDqlhnMx0ui3mIyeYsVaaYmRVUItXtmb25ZNP2TOIWIR
IUYmLZ1+YB+SwKtKnQbsmEVTn/SSvp31rib3XPXLCvsOKLcnA7T5TEmuIiCH68u0
XY/gdYhxchgtls3bMugBDsy5biOTo1O1jFLk2a83JyfRdXiRbYrljvc8t03yJ8Zc
9CsITVDXHH8hO/1rlwHwYe1/FhZTI2/ix51unGeiw5bCpqFT0OC8OQskG54+KZs4
oa7gnpHndq4UXRlRdAs+b9cy+ofkYGwOduZEGzoFj5XPCkIO+5tjc8I0rGb9Zksb
IPTgPMcvmDmSvKmWnCPyJmhHjQTVIgAuqM5Pgzt6SUFldPn3JVPdlX153IN4Btk7
4AlGaJ4tV8jGb3fDNjGx3tHC7DKKYgafiOGNcILjfKyXI1c7gHo81syvhQM8wah5
Mx5+L6XcncOYtACl5gKXXlsD/JC12QEDBC6mNePv8g8NYhjp7JfvOzfaBx6LxlJ8
t864wW9IX4Y9kRoz9KbzQSTZ+aH5rSwAhtltyVQZ1b8SwxxS8Ck8bwp1M8KXJ8Hy
0je6YCDVxmiUDlCTAPugHrfTDywzidZGwkYdiKa6gBLbJWAvSjGsIrvTqVBHnT/P
nwKaa+tQxBpF9iJFEZg7HOidPMwTrk0ffJNvh6wAcwr5qbuY0178QFo4zQMEaxZU
s9SFVDRF8pZd9KMdrl0P8/GwZf7KCk8d48r+EDfqf1AedCvHATLoeg2L1xIYyI4d
OxufI2FlREbo4qeHktFm+xMWg2d+NWfpttSK/bI7toZ3/e3XSysjGjyhjuJ0IklT
OR1PdZ/Mv4wjEAI3Pai5CvIZDUzQJOibOAyxVjw5mFF6oAN34hVjFCCbWlKr3qpH
uDtYRelROKMFEXONMyhs0QyCpbNFrPO8IDxEtCMBsXQAvIuvuClqMJb6MLUQ9NjG
RJeJbw8Ys7OjSJzcZ7X2KexhNBFqye5FffD3X4qIK6XygDVisFCRDx/XLSx/8opY
b2751sI5YDvYWrv0/CY5CXYjb0T7LW3oQifUvvy4PbAjRIqnfSxKMW1XN2qiO7To
eKBFohT3dRTi9UQw24aDoqTV1iupD44hVCI1jDlX/XDjnRAhxrChQitG764DWbrw
fxOTw4+6aimmrlMMIAg56bvtUc24QOU0neteA7KOlFal/c6XDyicoOQEYQaOHmN6
PYY6qwVZzqz6A75xKVLEaCPxn8tXGssZBwPnLvqIO0M6xkj0XH7olhKsH9AaOxBy
tVGPJ8srSzGSN4k5jxdQNNJUbTxnR8nr7kMNRajt/gb8SVJpWVdT5E0M8CJRWJUQ
QhVsUXxgs2jGD2V6nvfu1QWDfBozQB2m1Ybk+styGReZCx8iVSNzShNG1iQIGxrT
n77PVp6g6LAZO0bKyxp9Z5ya3/yNLxrLj2arzVfKhcJyF186hISOPr62CsuPZBv3
rqZFlAEgbvLUGV/6Wyrhif/BWM+PW5vv4P+ot7K8HKCh3UPfI8b7AfbLwCw1KafT
RnPj8OPKWTnuVeo8FAOYPse5B8dPq+Uk7jVgfwC2ua3TDBg5CiR3n40lSlE+Z8wa
Ob98DFsGiEwqadmapF1jtzrHg5v5Gb6qsOrcx9p/mlx0UebQl373RYDF1qvSbHQ7
ZbE3BXL4NKzQRDMtd45s8yw+UDDI8LDqWylLrTYV41g1nUvdTcpjtZyAQt6wYM6p
vUktv2N/P4yyURGrEYTUQ5HpQBdkmgZo1NU7RYg3BLmqlB+PfFpT/Pt0HA++ErXh
Y6nhiQ58xw7eEJgwirHfPzl7jCb54IEK5CLK6KR6DsKZozwV3H5UoXAWVDr7qRqe
VeNSbzkG0546H2j1qkzuiOyxCtoQ7oAUxkWEBaVfZGWlXcJvzS6jdYHOb4mqL65E
Lejfpo3XZoMaGagg4K/TJm0Co6IZ6t+TanYqDBotyg0z3uFQH2WZp5TDke+iRPvR
dCeGCZfc3ZixvNGJtAq6jDLNoDzXpE/N7Ppbh+iBgOjXet7bW1aubpLMU7sgWqS3
icWPWid3vz+bfOGQdad7Svz2Zb8OKV6IUpiROOrphGGo2y7NqFVKvKLPP9Tnpdd7
zjuRkpf8jDDk8WXgiX2ZX4cJ5fdNMyuOXArZ1MSPgQi8Ld2v5hfSUvdIYA36AewZ
uqVs5jIDV+Ogv3q2p9loGRECZkK4tPE1ivhBIUdjSqTIIzBJFBiVkhTCDfu8+4iY
h/2e4a7z6H5R9fGqSePgtyeHsPeS2EQKsHBqv62Ble7+seJPdu31nUlAyTO6nT/L
f3v7i7haeAovVgdmJtbTbASWuFMRlfrhWJmGZCdPfvSnYFcv30Yowrj3sg0lTw34
gPPYzAaq1z0FArINeHSBmItNukS5JhQ4Z5os9Yz2ke56ia6E3uCbUVjtTu/5VRBg
ph85zjQrPoIDWv++RYWNM47yneoEvux400xsjmxsD39qEw+JFV6c2dGVdcfP2jLB
bBd/f9yF91vJ1uaDIqB/9RtlRz2q3FL1obYWVaNuuCCeJ3xFPjTKD6VYQ2EGHc+9
GITCDIFEF2Ew48g6mpyNA43uV5PMbwcZ6emCzFyRpZs796/EQxDc6w4mzzTdT7lA
plRkxjhHWY/zg/8FfpjOMTPlxm+3ejUMJtBKpceZrWzBkhwRANdrrEcp+qkOwmVR
2QwEKo/g4FMue2b/BpSg/wcTCzY7jFc7YdS6YKOPj0GxtcAx8Lry+/LWejFFP6Eq
YOh86nVfhBXyxXC6M/1Yx43G7oJADtWnwu7SnQrz8y9gAlO8vsADyxeU3W/qq7QL
44tG2o4iLfCfgrVnQ00bG7uLYHVnyOknld+oA3HwAABF/GYzZEtq0k8STil4aPES
wCGvkAEXOKDyBl/phmi4FXg6QwioiTpHTHPqZdx1m/Y6vo/gqnXLbGpxysWDElTF
dEjtwF8W1os1vpbvFraR8URU7u7vS8T4iKheqKqBxH8skHvfPnX145rGbHSJhpot
Ya7k6+g2DfkQNldiP1UxY2nR3LjCB9PRWGKulHQxol0x1TD7lKQMP78kyUfGFR+N
Dj82Asg0nJsbe8l78vZc+7FupB63FzYx+4V5ZQWilxi+nuPeY8wgZY5ms86ZWi56
xn3M8isyQugaQGzkGH+33+QkHYCVw6ANBRLyz9IGr2elv4Qpa+NznTAiZ580Q4mk
Y9QgzWxb+vNg+eH1wt+u1PQcYAKYSEQEcmPRo1EHXk2Vam8US1d4n9aTFp+OxXU9
hURCxELhbRa4hyhobTGnetxrdQg5KDnPcHl06cG9IJXe8fJjbjTd+SrH2kLQLnOK
p0jhMO9BG0SgGFMAJH/eOQJn4d41H3TSnYyEcQtmQV5jNQqrUKHCyFWMLG853wZw
S20ByI5V6ic/YPbr1MPTl+Y2PZBjSHZT1/y3BB5+ZjWW5ZhChyrFhA74GB0p84iY
jsUJA+KMV2w6+qW/INu4KtIfQ68nIz55p2+15OyxXSXM43VN4qz9buXeI5xUWEjf
jmcU9JwGWPAL+1ospl7qAGIV101/H/80EMAVQ9vPv0Cha4XU70CKRprPFgcSI1xw
yXUDU2OlvI20n2GBurgJYzNrV3VlMgEQAPlUXL1ppAv5KV9JAZ4IHgCeulnX9jKB
uf0LeccaetOSGorrY76CgEQe11DJcmHsSwKUitOCQXfo0eVHbejWfqVzRXROQp60
wlwChQU+CeqAwTKoGcp1RQ57/Vrrj2QshS6XV2JFKWZ9N5uGVmmG+0FAfWDH+0jR
XpTCH1p2CBIwrdMQ6dIrzNO3tfgg2i3Mxwvq4MyU24KWMJb33TVocvwglIqXDySZ
E8Yh1zVkC8KqL5N097LQdZ5Ah5Swbaop9t3FDSl/jI1qAIj2I/90/ALk0In5dFmB
MpzraowhwHT/t/Jn4iwuF4NHZkE0kFOLdQAF1MQjIyMtU50nw2ruNw3THfsbqEqg
8TNJKi5bgSQKSBAUpA1evmEDeoq3kA1JYENLLRtdOpq5bs8Hg6hETT7NjeW7GsSF
/cEJ+Bz28SZeFmThRe19DzA9tbsxASTTToAtOcYXoxiaz/Dk2lljG/3wUeFepoFv
4Oh8q4aE6Wxn08wYE3T7wv6C6qLwLY/8SDASwtml2khGZ2ez7yCw8UA2xKin+7nG
TTHBBhfmryieOU8U9gmNoFw4cwapozFJTY/6PEWM3FkSIwBx2jFB+DAukna4pHtd
i0mQdLGU6QTEuxfPMwXrfkiId7ZOHLDL9G+9L5B1POntym6SUjYLk4vGj2Q5FZup
r3tY7B9M5dnOJtAvwNW96nzFSIcHpYPPmwHCG75c90hAao6dvPkMl2VgSMDPjUxP
Rdmabaz5Dwccm7ddO4c0c9ELU9TQNgDmUyUxtY17u7zTkfL7q+WXduai5RYL/6fs
X4n2d/Bgseq0OU7BWTFSCnbOGvavG5C3n7iHCDsshMZuG+6Kxv6+yd1Fmgg1dBvD
eTyA5DYgt3QDIFvpEJosMAQPyoBDeVrxMGhxltEBaBDx3yhDZcGZM51WIK8dYObQ
Dy0LnGlAKUvtspBygs8jXRHdliqXBX5Fc+Cxekfr+6KPyn9cFoEPdlcnLhNV6Ws8
KPBXjbFDnSRlzRjH81l+1coPPla0WDi+WXGjZm3Con7y+1QrLAX9F44/TwTNOS93
VjOMMCTaTvcUUtzfzqaPusEnbWBJNnXlanU3M/aNU5wjB/y4kLj4ndz0+2lE1Wjo
PzoYqCGNuKcjpH2yh3UXWbPIuhoLBuI0A+PMaJ7gP+tAb3oofNXzHeoKqIZai84i
a6Vh4UA5VcwZU2JZiQaPZJgH4ymLkkGBggDDSeO8ytB+6DoEjefvTY7Pl7osf2Fo
4HNRMQf17BrqvqhLAlu4LseJVz4KaHTKUJf/L/RRnaxD3MVJM6oaGB8tdGeaGvrT
gb2vswNRxc80j/6F/JWYlv3YyQIOz2lqPB7lvv6l2xBeGbfk6vWYnEbnJ94n+b6I
67o2UFjV8AjKiWEcoJ/abtWOHoQpkyS/y2KiVe3/QEM5BwzChx0lQBn82Vou0YTt
8BpSB5yd5Hjejp1srrcKeFs0f4HQ1etxyeUJWUqcfn5jG/ujSa85rneKJJgjWxa5
2G2+llBKHoUReOpcjKtbGLK1grCLmiNKmmguO1ozVoMfnpDsf1LYKDCchxVlIuKi
j9YqlL6FpMNm9Iiw2JKSXGLxJEkSUZiI6CkxOXKN+2EuIZB8hr6DzOTNYZ9tJLca
xhy/cgdYpGU17xgzNmqGlzaPv7bwwNBHsPrKFcrRwAP4Ax8V9gDOMhouXEuLfYaT
9cf2vMnd43VbU3J8mHe5L14swjVK1IyGQIWqAb9EmZkI5isNwhQxG/ueMg7Ih/4z
aI+67r73apu0RWygXWSLwFfLEERacsjCg8stF95akb7k7usEgTRaP6IPVmMxOzG3
8bARG7Uj3buoAqNv36apj3iiHqt9qnwiqpVMplMg3axFmaKvHNJetQC28M13vLGu
E5AfwpFNARsGwZu/pB0bSJSQ8+IDt+RY9ezK4FtC/5y51h365riCWGfXC47TWKvm
Vo8ee6pon4414DsPfles9dA24c/HOsya5HFoWYZqVc8rD0HvdAdw4a0UEprnwu8Y
I0U6WCKN3QmOK05EkHmIcbe2ffTWl9e3K6/mKN4Hid0uPAVQKthX/F/KDx2x6s8N
6Z98dF6b3rFwS7jb/aBUXwtt1RIiZ6ZUBJg4+DTROUnDpwnN6nXkKqq7RvC0t8bX
RieDzlVar3bwmzuNelJhicWghZRhL68Jac47ukDbHD691L1qBUIU5JpKkBdg+2lx
R15cXrA6gtjWTxTdtd/N5reWhgT8IKEEzTWj1vwaq0Zv+BuKChXmsNVW2yqsrcvl
2klznz0bKJyBHSsHXTxqnoI7BH1CRt/nLdHIndy0cqG0U5fmQqVw74uU4hWxcGvv
9R1BosrPebnO/cYgDwomkOKSYKNsJjiPrKKn7WogU/E1WllJ6vRJrE2oKOT98Ycm
kSORov5WHfCAScQ7iRacwpNrXh6zvWCeZSRJ3wVuvlNM1FsZE0lO2O47HO3efLIF
RLKvDNPg3yRm16j48q2wpx1QC7BsC/uC8Nka0BWv45+3RFNF/aFbeVeYna9V2a2x
6RCqTjdGKkJcrlZ2XCF3+DBPZEnMUQWt3lrixvouIWenGbhZoD9MzF3duMuFFG96
bV0FmexOxC90NcPCRWL4q7bXYWY2FCcsU7UltPg0KuBoWhN/SY8ldxJK2RMly7PG
vdzZwgn3+CVghi2xUHpF3vpSEBExK9tFQoU/VFOiUm1JEgmwP1aLAkWisInDchzr
n1YPcKPyk0Ny4MpvvZhTwKXS8eb+yGkjKARiItkhqkaerwsMPpJs2RNMTjDGl4CT
Q/qiJ4abfMUYZhgmTotKInTVn9L13X44olEFCCulMAOvGj98+q4flE9UsyhMShGo
33feH3RkuGrYM1ttyrsHyGZlQGJ0dxpdAA82VwedURRDSNfJhNpV+J8nM7d86XV1
P+MJgHFq1Pnh/2z29xC6fFBQe9vfWYyw943oI0aTGPYy24cJMcA+jOO/3TXDrmEV
Bb3gEZsJ5Xc3ZWCzTswBkAYFo6ylbKSjj1FFOShWV0nJ/y4kMJTqGo3hjlZUveM4
M7WItl2XNBEhUq+ojKVy/BiEIICqDpsZadZlMENkfHN65/ERul8I+9inCi/p4vpD
GWFqXXaliak5eoblSGXM8SpA8SOT3+omfbJ58Sqc9wfgyIpBhXGjK2IRmUWBos0V
NRu8r9aDF7gCRDVRzhRbqBHiLCvUtdGspelbxT+ZPoY2huU4MmkiVrEiI/kdYoa/
UkGLMLNli8coA9CMcISW+m2vulDC36gyCa3YkMj6RlT7AQFhE4Pzg59h+Jhcoqmb
ChA2XD/OC1niMOv6I7CuQY8clCjZK/I+qox751JsY3gszRmbKsCjdhb/vFeZqjA1
WY/cdDGMJM6x8St4vVpeKAG09z1uF4CICVtIh7cc27ASO9wJuBenjSs3gxL5KbeS
EZN9LkZtyiz8qhyy75tobjrXO2G3gRuLVtjZRg0T7tcJZRM3iLONNOeJwRWGcrbI
WmiCosayOzn22RJGP89ot7tWi3nS2Y89IERO9Li2zICruz6x58SQWvY54Pj3xXzb
2LwV98fohn9sJ270bXTGD6JjpMkKpuNEkcAV3cPWNYNuWm1awq3TXMLlLcaMg7/O
phWCz/oUrdweyCpuHO8jQLp4a75cCakiYKFM9rzxxAgNivLUxl/fEO/9AhP4BsUX
kMWH622lY12T3ci2GCqQu4j2zj0mHD5pi6XP1Mz99Tp1CQMbzefZKYvmHXx87CLM
sEUV3W3wHLbbR7D1cnSGhUtul9ZonaDRCXmg609ufddWXKxI93l6VrfUy0QknWzA
di/0C8YLVqMJHk1yLKnJsBJi2Yv1W1BeCKyJllRzFcnOD7evREdxSen8s0qOYx/z
Wl1ombsgBPxHfI4ufZO4t16mNGkUM5c0irWJH6su9LWry4D4q+EBLQqlJ9qtQzLc
wVpqK9hXRghMuxbZfFbFVxnvxg5xdNUlGmJ67NH8yjzc2XT7y+let3H5hMMZvuEK
BB0PQHQmYzsUY/0/yn5NuxOQB5MkEdBH+6Q3zC9FYpD7/X5mM67Pxp2ZQnm9Dibs
djecc3q7qLG/QIlO9z+XquPsFnOtqZ7ypLWAm6jyLgOSizy+wRzBjErEFKL+jnJv
rlvkK0U0sB+Qrv8LDuf34G03Gh9KCk10UO4dzlpbEWQxKAyMTn+OpCTp/fBuoVRa
UDdXce2M2CVrSwr/2W+0wuN1tI7YT4P/EWFEbD+Lr9mSHYYJeBWnoxn35vAaolRp
XpqlqkZ6zAT4fmDwZuPPdGts5ZUSzMmPYEAuA5J6JRwryqm4Md+z7ha9U+VQyu8j
ya+3ZoT77EHib/rlzUpYc/rTzXhEzx5l4X1ps5gtCDM4hOj95+rT6gPBl7xmzIXc
ex8OcuUuUodZ6vg7ezBKlip5/uysmCwAwmZojtPgBMHvj7GL2Au5fEL6er3yNN+d
wMuWFy11PsKYzrVoKcHT2hu3oNsXkgHGM/SzrIZONL3JvP6ziZgU5CR1eTCBcDjW
w7tBvUuXP4iAh8kMbPBb6vxNwyag6OLZ5F7Wq24dTSidGRf3KRBunyewiEEV2H89
XJy/6MpxdRbYwUo7jHUuF7d//jRSYpPCeDL81h3ItUl9PJzBs0yMxfAB5AeOljUO
q9GO41YXcu7Q4GBjXwFXFsbRd3AeKzFs4NJPIwks47BIUlgRoqiYfWKc4kRXUVER
6csXC6u5JPVeJkyJkH7uVN6GMy48T+QV86E88LgVip2TyXiK+/+HLVIFBdkw+7Ri
5P9VeQooyBcmw0/RjQHUGkjJINtfsZG4NCn4LOMfn7akqLSogTC9mM5eNpee84xl
2Ogx6gEH7xoqJBMp9ECoz16KLlmu81PQLFsD0b1iWlGXgqSinTJELDZFE+EncB0x
kZv5arYNsyGmcmt50GSBlugzA5EcXw33bDCHEwHMZG02wzC8QsvpPV3EK0aJgsdG
SksCGVaDakSwzIoaeL3hAit4NRaCrj7lp7JBhrd8ZaDuIbEkMzpp+KF1dkObFxOW
VgEVbX3Mz3IXwWZKcw/zlc14hv+ByUZlOBZI8LI7+qU1Rb93w1hZSI5qgzStsEvp
B+89+d5o9VxnN6tZ4xYeXNZkiN+6VsUf+T0hFP3JdsYfqfM+SrMoOiPff5vXqvAO
GzqpbOC37vYXm0imAjcsQiqLIItZ7e1Oobxl6Rn/2zE8x5P02wv4j/hyedBlM5Lq
TTuU8JAHnjerTTpKNP//ak6UM7IWOKyaumH8olkEzaCYl2IhiegVyaj3dBfcreob
hZzEiC5bGz41Njv0QvWfkafuUBFvT0cr9QsqmX3UU0oqnG87BZ3KBLH0xRayGnXY
CQsWb8OrZedghMYGUApAJcyPeh+0Fa7BKfwGSYrWS+V5AQRvY5zWrauca2RCX4FT
p7VMMhCU6VOUaP+po36+cmOS7xOuTcr2Hw3goi4WbR/Rkdfq3cYj8xwpHJi+mj1G
GKWChdvoS9xq8HZEFhaSJc2k7Oo7cBBLPHUHwjCJdzEQnVO/y/5LjrSVTeIjuLZ6
uhB2qcC+l3wQA/gRdORuOtPpe8aY+BWfQksb2tm4kdHWrg0dRmeCLiO/s72fs1/F
4QyHgTVmmL4UPxO2ys29iJD+e85TZEpJ0pvHBawkQo0GLGQy7x0XtRuKFoBP5C9w
HTs2J34k1AtjtUmUwiUxYyOBGFSJj45E0oRtf9PoCx3SGdM4xxJa6FBfMeAYP8Ci
YzcNOgJdic8L/l9Xl/OmH2cbzdKsOLs5isg/KWrjeFp/vLod8ysirh9yASV0yeHw
2AlGF8zOFNewSGakpqes2Jr/2X/tSEJxeyrc2MUIOEhVpgZrQg2jhLkOwJAYaas9
dALHHn8SCMsRfwpkX2NPSZOuNsajL8oVrqC10QtySrEIf638UQTyF74tSp6Z2EDc
HhxY3CpfYmiH8DSiut8rN0LR8y2btFb+MOoPHFFjw560P3xsZ/sbdkaQqjr2BzTu
vrrfoF95gbNDSfR2EPGn/eI8kzbifrxhn3n68egrxwLtXohR1zoHew7MpKIJDYAS
dSDzXk91SR5SoyS+NwfSWTi0uZa+ED0TWaqSQnrf1WCEszN9hxRPZogBwQjgWcJY
kTGtM5LMhvIXDivdNZcAnLGYC+KOHFq3WOlmdBhc/LFnRgINqCQuvkF+SoMI1vUR
eMuWHGCS42FpKnoULmAywPAeY0r9AqrfDrA76QL0dzuM8L9YsX9ESrsTeNUlF2iz
BNQy8ExZul2bUPs3KSX0DePA4hpB6LBcf98XTjtGUvKljGHHJnc8O9pKp6sRiUu/
d2wXkCXhGtj+cUUhAoqAKbtrQMf2y0jnYQDuB8qnzKxaKryEZ2McJAieG4IwasiL
PXj78SDDaLRBPhmM0HHMpYcRf6PYH+k6thCJFwCD0qJcwgGepH5tVtwm39F8kfEE
Oh4LyEFEUwUnc78/pDUFk+XyrI4bra5IekC5ggzm56n4xWL345jkxwMpNrv/R9wT
u5VKVK1S47aT+vLf+ZMYijsScoHEoB08bYCrp52/YSQ+iVqCofgujBKODCKDbxMu
SJKEzQd63iO+tPH8y9viv/i34lN+XazySPpej5FFRpr84XkyZaxrcDzhTK/W9+UY
MI9jWrDuL9S/CQG54Pt1J6Fw2YLF9GaPUUcqb4UzIGKeVdIqEfMRilDIeYwOzOwi
vAqWl+NPEZEe0ZfPhjkaSWMnfuMfYXRPOWTI22M+gX/kk/PKVymuKkSoQKJ0mHJe
f+zYQNk7QODBuBUrxIq6UzrjgcVT6K1/od9OPx7lLDtfm6gc11RjC9HTYjhqh6Om
XK9OAKRlJoChqRvAMhsZYXkmms4lhKMAnMt12eQLgvbTwyFILi5UUJCuowZeOzUD
Qrh5eNSaVyDl9wvtM5FP0I6gw0BcPD7G5CaiZWQKDpUbtO9raKb9yrvVf449KC7G
unnA3YbXeD1bJ905gThsUG6PXWN8JS5lvGk9UOEox1Qf3GdPpF12y6M1cDt4bPhn
LbCuxPfUQwhHh6AZapLR5TASxR2VYpKJ1hYUNwYTQEHg9s9sxGjVC2IjTZooxoxR
rf7pge3zdc+/t1MDLM7mYq7sCNOMjy26IfRg+MdLTJEsdSreaxaEyL/KN5OkP36J
HOFw8WYsOPu8MVd4gJG0ItBdsuVqhKCFXCGk4joj5mdW9z/nKaNKciMePqhEocd/
0h++4j0YNDpb4TVWJWWgn+LvmHweUIxDqiB4wJNGq6WeERiHtzFcCHyRcwVMi6ji
fmZIH/XZ6veJU+136BxF/VmFayDKo9bHPGKFP4h03gXYPC3A3pYkPx+fBBXw5qF9
mIfA8JcbQputCxYUagCsaALjZE2Ckkn5AXcPl5jtcFTqP/Ru3O/QnqEojpfv9vXi
xJtcxZZq7MbVEZ7YlSYsc5zmtfQBOjY1BCeSn6Zby3h9/4Hvc6NOBixQpiXtdlb6
CIML7JqLWnVA1tUEWKlddgBDWd81OGIFC7cYEdxWTP9jFvpvInpSKwC5lpjzIfh6
0Hkdc4TkrX7ftRIZy6N3HTPwxpDHVZbqRDZEihETFSlHuILqFl+R6Eo7++BycPDc
cb2ViXVpuZZ5evraeoRuii2vT2U+hovWNsXMhksSUTUX6OPqMfAOh/EE6G7jDRXX
CTMfWd/3BmD0YR4BrglXMmTVnyh5lNbUYJ6cHPYafcmElenG2Wval+zLWdpu/sok
WgIlKY9iBW/oz2EwnEQ+APJ6U21LlK64cqJ87xOJr7bPOMSOTT7u2iiVx+I9Q1YZ
ba8fSulhDLh8nYFgo94IYJOuQhaeW8a2pacZl1wssrGwn6GFnk0k9DVXVzDkmJhb
eKiEDgWTl2hW1rR1YT8eva/LKPNCxJPDYvcH1sAV2owObflCJ9/dvxSoHCxjmmeL
yNbEzhNZHUGc987WA5KQpsgLL15Uf1tG2Vnt8zVxuVozYyJ7l62i1lJ33kWsGo7C
ROkUt/ZMG4MRhKFWq8A2+PpUK2+JBpux64YPbBCBxob8gJgcIe4HQ1zIfCD7YVH0
byRdhHRbaZdYhU0eO5Cfk02Bzwf6Fr6yh2PPQgsnvGnbbfX3h3wCZsJJvpJzEzaV
4d9llX32rffQomQhdYmrvmESSzb1yBPDOwBK6Mo/oPzLa1Rg6t0CFaQgTrt6xFNV
Hh106vNRMJlWoFlA1gcx9RCKpvhWNo18XndvyWhvb7INzaft8wCER+Q4IgzK9ocb
LFTIlHHFo5PLxzGapqXFgAq4vIseKruDn/O9/3/Oj5njNubJoXXb3MSrH0sA/l06
54yl8keBHHawOvMMr6KzkjvKsysFa/2b1e2lpL/dZTZ/RtvAWtrmq4ZlNq2eLhGp
mZdpsH8qvrrK1bYB5fxTzHE8viSlvwc0iUAzyZ55btsbNqOedNFS4PFPlkUk8uGA
M6cHXi7c59kGTuS9V9qotcjriQdSS/lGZB1DFQQ+FHr2YMY44UY6NHhE31CzX5cK
JxwGsL2fM616a9jO01Ui+QFi/iPLym0J3wJRGQexDBWXQ/1aqKL+oPwH3r58RJT4
v64WKLlzmOqNwitELfC8kzyR2uPzk2Pk0hHOLB8oxNJtSR96iPwBFAJCKzLQH+71
WElr20I0xN50zq+mGNYxO9XxiCq1iy6ftMe7EvPZTU9LPx/bSVOMXeRZ7cQfiWPQ
bdqTFPDvvm4uhaZQYtwS2Lg+YeJ7ZOgM6jx6wWELRLGoXzuouimBbI8PJiq11/ZV
al1XT/xFhTN7KPok2VAwJgcuhMVZfnmRV89J2bXt51Aum8EmOaf9uj/VOnHeM8zp
1ERPBf9QKn6wHMV5HPfKjp4v4TqJdN/M5GkYPKrbX8q2ELBXFiLP5FnoxhDJjZyF
y7mbe6gmfuadt+y4clchJNCKsXr8xkhlPoYx6xfgUEcMehajCQOJVvZexEQN8n8h
qwJ0MQN9TNRHroQAzxM5ezqa1dY09XHZzKS4vWttRSL+5FrNQNP6QejvgLBHNHt6
gANzx1fi3y84zSa9W8trCBr6oLmc/PFHp2Mnvuu+Gbm/kJv0AXKpse7Zr8wMkKgs
/fGpMsksV5y1QWH39as8YA8sa0Ql8d+k6EoJ4azuGZu/ja49lADtRs8YRkvSFdCE
c3nBZXXeEMSOcHPHKjT/sm4C1PhqT3M+jl2Y1JQ3HtZxG649q0/4c2Vx+yGQjkMF
p9EOvNvnfmqJF2rJB8eHyzbYsLobJtZ/6Aue3AYcxmRIxJliLPWBEtPF21tCcXVc
wh63S+TnRoaSwEkFFKejgs2lwg+Yet2Kz3k/eQQYDcOoQfuVRawsqoVQzKAHzaLF
E7HajFDAT1IcdCsfKhp8Dmah3rIpfe0BrRIwWSOrh2F+FUWtxjYZRJlr/Ybgtmfv
sGaxPR3Yf7JbEO+uL8HwvH0c/4mchcACnYX0KtxVNqk4EeuPN9EFjzwGxijkNupO
EwYOv/ZPrbi+A0+zwzuRSbkGQVmSMzUXhYKdPLhgVQR9rXDe347FsZNuoFwzqqOG
q0wtu2b1q9sRznNE2y3O+XZW2XbxR/zjw15vO2YepY2gjr0w4HsX2yNFxaowKR/g
E6rrVJGn4lEYI5Gh18tr6Q8yWmfDltMQCKbzdt6f5/SjQjR41lLHBTFQtUMz22fh
OurIlaL1/DZK6F1ZAzwj15s9XuFWFD26+RVFm52oOyp5bl2ntDEDiwUNDNcARtnt
oYNm0RwmFjfMLITSFPOznNB1iJqPssEckQK4yNazGXAh/8sDV9gUGCA7Rt7pfuIB
uBaggSCivgiZpNcqiW1ogy5nTKCjC6awQQMkHzjci0uaa1rg/ltklgdB4KSi6Guh
8dhgoazV4rMjPHI2lLtowIT15GpYQYmEBULEeLplaw8+Wq3n48emDCTPhejavkk6
TnQD3rIs8vtO5wNU0TfEYDuV3Qe56J9Hy7MI80Kq2hLo7ALZBxyAZ6tyA7glJ/PO
3GxdGvihZrhl3eVvU+8XDP+pFc/pvF1UqIB3tLZs0Vn0xmLT+Cm/Z9NfKhKay9Fg
ZjKYDkekX58G38dnJ6jGveBItSqRtoqhtiDpKx2Rhpt7uLCotL1HkrGzVGrojPZJ
3fHcLMzoK5vFZB8TildhFXEyEL2F8fjgQsHGhaiJo69Wyy7XgG9XnZIim5Zdwr/+
jm9B79cNtJE1V2Uln5m/I2F79onfQaNr1GCmWRufBDxqy24rBaNBGO+dYgwnzYbs
TvYGDWeI8T+3I331H4Mbx9g0KG+bvKcirYw7uWpf+OvlgPHCyyv/IWEdZ/7Jj+YH
DlNlDEWNGb6tRTm0Yllr2BNDfMx2Ax1RRqemEF0wrh2uvck5rDLOx41G+U8DffND
xqnXJEOR7Zj6uTsp825iED5fedydTYhRjXHbtOXTofJ6ru99FKmTF798i39K+kHt
4yf7LYoF+fLQ6Jp/GxdEhgUp3s/UmXVfkKGbVHGG5aJm7Gzx2MQI7qRCH5SKcfeP
IZSwNJWC6DgDFlIqWsdo3HT68LFrX8Qx0gv4mSfs1XEOszh145JD38CRFi3G11jZ
klfFx0S8cWOvnPcRJ2h689pGBmXtZd6KfpPVET3IHiDpF+9cYHljEwjwcV/oWTw2
77R6/CUXyNCrxm6Cf5IkBdcsD1/lPj2/6TN3dN60vA3WhLHPawwUuC8Psf++yBO8
LGHKqi2+aU7YhMvIjpp7uyfqmuOA14Z4WMCUHXtqclDTPUy/nAGvu2uJSkRT9f/r
rz1zg+WNK0hzy/tZAqL0sEoOZ1tck2hTNbll60fnDlvTciDS6htSfcK8oUNx3Hep
5hUM+c+IRQtIjwKY/l5s8JGvLuUh/Y+1HYOTebUpSrI4qbUhhXEuhoKlh0Osdnep
G0kMt6Sr7WLvTguT/AvqZMqmJIKaU34/X8cPyNQuoNlSHWxZhn3DNWD3qjxfvqhR
F9UT4Ix+w3r6rfxmxTGVkQlShiztaj88FPPgmZLGMa3Ph+YKD14sVCwoha/y93eo
inZthlLsLi7Cr0fGIjj02Q4qMjhszgPBReJiHppXw6vg9YzZrti1/O/LmL0FgSZb
77MdTU0LHBaBkoTsdsbt/VxXhfeu6kdajOIeECMuvbeqNagx1cZOlfXLg1jsiOGB
ujMZY/ZCdmksdA6IRMOfUSAnkKjS7u+gddMj1UGMQrrSdvuCSFiYj+79eAd7yBbT
OFaUSNi81uD6TXChUHlZf6sXjvQiuSyPuwi5qFDKH6S0xJYhs7gmPBgwRrxgTdNe
VGu1qQpzLPBEupMtvcgvcKkYgjTCidWOqxJT3zMvbzekI+I4S6OPfDoQqaq5IFrr
5/N8ggsSV1CyuZ2/m06gMNgQtuQvgqOd1Sx5Z+UXVJImtz5nv261zrl6f9auGLtd
H4/IrgOnU7Ow3iXtoHWOf95fAM/Gd4s7jEopYiZiSUVf0HLvoaFK4NeO11LYISSb
XrlJZFk+4aG7GxZYBFAQULjK4a5eohfDVhhE0NNSP53km4dVFiuMjLVpg3mAZtc+
Sf4lrPMrnxtg8msmXZ6BJRyxMmxIYRNP86wR3oMMLjSM3l+9aot6/uGHhiCuzZ9F
I/rHUxVcxJuGd3ne5UHcqQ==
`protect END_PROTECTED
