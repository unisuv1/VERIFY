`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vro/QvqMAkFIzpdsfPGMCSF48UK5RIv69JVeaPJWGIZ1TfpdZqvJDY35FsixgFQV
4Z1jsODkGOeSjboO4YLF6CvZcwHL7dA1/wngtkLZ/js0D4NaWOgJfrq+lzk/J0i/
yXPwPo5ThZfAseo2V/Y425xz7j+PtK6eSYo7kqPP3l7CSKy7ZbogbqIdCShD4Z7E
0+SrABHBl0dFeZ6LbiBfaQJJbsucTxiBkQjJ2E0PaDRhmatcEOKTiAVOE/oMQjE0
Uhi8j7NVNaSsn7IVD9hU5U3WyKtQxKMbMXTJqpykZHD1OxEM9PuPmLxUVfS1Au4I
glcBcNH0+FvdRLKwS/zTk6vfJEsVYYhgY3lrqAmkkZRw8h1+cR8ixy/Looc1mqKV
mU1u1SOA1/zkV2gIX48Q4Vi93rPcGpnIADimmND0U7b7xaAaKsgJG/amRpYxDTTg
gyUFj+8AxpvVSDs2787YG/3m2pZnXzLDAaOZUngujXIxcFYSxfjpMShlsJHJnb/h
GXtd4HKxdcmaxH/tOgCClZR+RpxlQXdII0NDzQ9PEIBJXS7ZjCox2wpHkZ3GBCSP
cNYI47wj7I3xQZBDkxE90bPJXG9i00iKra0jmkZMB/7DGCsXT0wxWj435hxZ5zuz
e6sTFJTyjRs4tgL+uh98jNa1E51KRk6zmkwS/ZMNwzc3jj6/6z0TrovK6WPiIdIS
gjfp4oCbamTJlDdF6hNW+pdOQ9SJugoH4e6FdOy0+wiIT7hMPA9v67+/RyHpZDPj
DIgr+kTpDHbvWbsE3B03Bp/vZ37JxIs5lZw+iGG0kdEcAIZihNgJEy2IcnN5exRo
dTZ76NyXBcOXEYI3tDvtBm1tyBMubVZcbZQRoFz9GAv6rzTyR3DhPaBnei1JW94A
SZ+Cv321EapanQjFPQZx+2rCKKU+xLwpONvg7/zCXFV8FWqXT/eHZjv7I7b3JJmc
GOIVrDWOskOqeBcYmgHNfD+FUhyTDdRFeHE5khA8/OiReEkE8wv6bWSKkax6RzfX
BOPP1OdcT1ZYylaM5g7Dyvdln0deIj+mlAXTF8819ckoaHbOG5dJju7w+nxzoHyl
ELZf7J+5yv+v7sE3qMGiUmkIxRDrovz7nCrSxCPAddXHq1OGFVzRm4v6crfKEIC0
0W7I/B/0qZ9wM3q4j13zW11Web3yAYBJRfkKrSHj+88lmotobLAag+rjwKpmfWgV
Jq3G75FWt3K6MK2ps5cVPEZign+LDQBd+Qr3Inc727Unz7M8qj9KiH3q7ujvLQ2j
GvlimpnlSjOeGjFgU/pzXqnYMeWtP7v2r0oZUAF6SrWhDAohrRcOJZ6Vfan2/a9X
xs4iAn88TD1g/vSPFbJPIyJ+s/f2ZFu2E2ycFiKp3Atj6s7Xpb75C6ai/Kt1mUQh
q9qoua/WUtfxogr1gi9XGXh1vJ/PglsNe1GL4UezcY8n+gyRjlIainSQhYt+T8SC
GVkz6+9uPAenQKUlPB5IRLAeCce+tMC2xBZSfCErcVEd/3L1FQ4664aAjQGKgUGY
t3YfBjDmqHd8gCpbvAbUZzXW0YDr9Ng+8l65Q6t3QiEAoCDgg9sBlGODTbZw2otm
LxhBjoi01XMzDMKQwyWiNcZJlSdYuKgA2FOqmYxoJESzVtsR7vRiYPpKlF2nZ/yw
16ciIhI/Bon7zI4KLVty/yDFO11m2mAnDQQYfirfkq8=
`protect END_PROTECTED
