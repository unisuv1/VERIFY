`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
W2Zw3RNiZgMb/ZusnMMPyFz9zK4z9afmZ1qFaQ3v0AVekGO2kyVdPfEdHVkoEB8K
CRFk0MzrAkoTzUitOeIQ+z+7K68F3zaUJYtI+ItM0A9YK8NBmktKoVVeAKfT2Air
uxM52Jzjs9OBkj9b3teYev/v71NJIvTdcvlSLexHFAidoPj7oPLMYcs5QS7BH9u3
tAMFnJblhZCZYUZcb6OiK/mBE+n436FRmnuYaZnesHOvEfRVQSjJ36QVyv+bCHe8
Qr7RQoB0vL3NQwIahKoJ4XLbiWXTOGJeXE6W7L4ckrEBWXR17AuFznx6LT5A8J7B
YARxL9Y47k/nAEs68GP2jPFxZv42NSY+WiSlCrObTH6cOTbxwJuArJ5Rt23GHxxG
D5Wc1Gfv7B8MO4BLj3ew0WNmQIB1EuPYFoufvENoO6c920r5LBa4+1CxEDAyA6N0
84O7qY763hA11NUYgaZsdB+Wm1CCo5W2r7Iew118EDxjE2PhFqJxMVFLMQQrgb3q
eShGtX77FqkQ8quZaCLLHZfFdwU2bbUBgW2rfzX9GxQ846Vr5S5vbJ2Z0dxOMdvb
PW/bIAxQor5gZ9FNQIhZ7l7nEkOXdpsEGqaVK8pbFdaiN4RZv4keUG2j85LCHya9
WXZyynftKb18WrVMsg4ajvFoPEmCWoTN8Jq6D1nYAE9Yo5oYKYPlHWA0sHMeJ8Nr
EmDFWfnqlEPNhfZqafb/Vr774FQoRW2fYDFtv2EIwMkLNedwe6oZrZusxfVeX3JW
pVMMyYm0hGFCTjiZK++8EIFWF8X5GbvsosOjfPXvIbfW8CLRoAgdhTY0VSTCDU55
/+UcRosqT2VqcU0YTQrH5ZpP06hx1dyjnf2vNA6kFpdn65EFQ593LTwwseRl+C3s
3YHnwXUTwIqpWaXj01qi//rGWaofdvXdztFtqnGIEpvwOYlm1T0C9Y/Fh/H2sU6k
/Sv3LpiKCkoswRT0MNtP5d/PbXgOkKWXVOIh6tiJZM4NZQhoIuiJys4Fixq7AGPB
6X5Dp5rpzKQfl3E6FlR6BN8t0fWpUB2D+Bt/bzEdMpX9irurLKag1k/DZ1edi18H
E9XN5xppN3iSF1X69PK/BGLXMf9x9JEkGS5fspNL9jfXBpOMvfvJZV1rnC+AP7m7
kgWpIAyuIF/noPI0HfnQ7ffqg17x7Vg6XQVZPbvRLEOxtL007l7dGH9JY4r3acE9
SH5oGUsu6yu+hhxTHUhc2wU0UnIZA9gdWCdMxLPhjofhCgZvWdMxCKIvQUnbwe8G
iW0avVNBWmE4rZTgQReMxZQNSIMDuNts0lAHE5Zvwl7JwtI/O0M5/UVORgRFmYV1
Pf3c0l1VLvIyynVZ36O5A3c5i0b7U2/PGJRS8Dne7L58Ll7Hr2VcWvCP1xVpfy1J
NBlvwbW7SJ8TwSK6AA23EdjmckaSGv4U2j4R+PEydWlApayuYvyhS9dNOv+KP1h9
Mwz6bV8+Bxr/jmqsLJXv05t+HkMQPzzM6gnaXn/KocnKKpGeS1Z9SpkBP4cgJxv5
hmD9/nlxvFKp4fieWjEke8TdbOGDyFTgh9fYBVziDbxD8ngzu6FOG66Z7BSZUsSC
pcKWEStPltQIG5jFzkJ6X+RoPlcg/hQxdX+8XFTko/dMf2YUB5eOnGVswNm8FFws
JsrbBW01dQTrKLLz3t+CjLSd/pCCOxnLH7c0s8S0pPHBqJ8nMdbZRGrKa3Zs2DZs
8ML6UMmKiBwd7zawETkDdhbcnjuGYUWZpLPMVY0EJQK2qhE8EVck2LokEAJA9oi1
6xEAM2OqTQ3tOEAsCq6LL9eofyNnSWjywn5A1MaPrA1P53gComGVTVNYA+MrxabQ
ljQtpjetcIpARVLnh/3BOJsdWlNDnQFmpfbl/AcnbsY6td1xUArc4KdB/t63AdWk
hJVCYCHpiuodBFc9ITdLqS8jcBaPcnMywhJuI1oAVzwUtKwre85L2CLkuQrbmzPM
TGcS9o+pcptnkh/DFCO/uR3NVGeepPDtOgxbMNTqXi8v5joL54CB58rVz28JioVm
/nFInwm2shnTN9paVgfKLTtuD3VlA46T3whESRmS7uk8pURAZvA2PaT5jA6NR6hO
v5qnPIBE/cSNOCYIxV19AvFoeGt54OKmGQl7iICQb5rNdZuVSlYjufy1B2moNXSe
UR5f1aUG+LV5Z8lPftC3LQZmELpahckhIIq8EDCzwtJbmG46APVvU0srvpMZ6wPq
SSQFP9XXIy8NsDdez2ntpvMZXjqdkdOo3tXCjoacD9LKMP+Fy4o7bOYmOVaR13Z3
s1cnjMIJjKoCrwFhxa28LT2QzHyGrG1E+AZ04G/coeG7SUudjL/SovMYX0+xxnyR
2GZYCqF5JJuFpkmm1INx+SRWnFs/U+sTQ7glPgbRHCvHK24v3fV5gpMNE4p+8te6
mcNG5CtSgXPd4K2/1pCPrRpv2dovpzSkNkwUsPJ+/Mu5eyw7WQQp534A4kXbo1Sy
2qieBhfbRLpjYG8u0dDaY5YymQxkRAbsHEaHbuOrAu/qS6uUOc+R3qXefYvOk/13
2RfWluGFK/mR43blAEJ6bCTHVJ45IHoxhEx40ExRJ17aQlh5mJvrnoBTAuoAU1Wc
cHHHmBiLyUSNA7BOIP/ZZabaoacPw4Va6OOohzLCLYN2TeGfLxTsP3ajPlfOKQzd
OlqppPY1/K9xtgqDxQbFbbEf3+UfB0h7eLZzjvl+wR7zgfEveWUqs0XLcfO8WW4C
NWzFd/G5ZgfPCWcW8l2f/ojW4MN+iq4f3GzPhkdAa6gLocawdcPqZCaMeAcFo9f1
YAnpNP7QZWpt4UsyvuIuKbmp9W0Trwc1SMN3cKiLyJk+TADKYiIhzY5QmdESo6O3
2Vkr8hTw79uhy4CGV0DbhfPermQR215v5TpYYcYBk4PDdAWt2FeblUUAPOfARjQY
mm5KZzXoXVfKo4aO7IJdVzEmSszfd9ld36Iq/wDHIfyMlHvkHCjCnJuAZqyj5nA9
XXNSkeVb9sF54y8Frn2YgbkjrxUVD7lNMZwx3PUPBvEOGiDa3ap9PW+8cqv5KN7R
yXgqPDaAR5DHt7lIuCkwqGJl4yRIDGIqccDBRMOnNt3cmC+75hWH8d44/uAXajbP
9qLGddowovL3SpxPXTFLq3BMVp0Tcp8PVbr0yihRbbGWonfNRH47ocbqNa8IDUls
FlW+qSQZVroufjrYfRrp01XVw/+D70TMuvd086Vs4EGNnZUQQ2NnP1SzFKIbv4jr
W78tDDxw/WBMJ/xDUN/43C0NuyT2AfhkozPiat5UMA6KvbGI5kjhYA1sEL6QnvHi
+sz9gsm/7iTbstOc+PJvM2pYP9M72F67rpZXjczUokAQMNnbN3+zjQKytNKBBsA0
NJNKFhC7Fett5Ee+wIGTJ1+5B61mbb/1NapWeK15ivKwID/Ortigso2ovI+VtECM
54K03Sjhk1PCpps462SvcZ9WWRMzZ3JtHoigHWQW+5sdZd0fwHmJTTyejyqAY5Ic
tKfe8tBgByff9ddSbaKGQMQ2JITcgd7jk7+bfnYBwd0DgD+1ekia299Zn8KwYt3D
HxLK1sdTxQN3E1lLmtoumq40zh9ZKT9aP3GxW3Jd9lY8P3kJU2tIQkfHTzHkMJ7A
SGi2aPZGxynCGJ1vHhmja92b+UO51M2kt97V8QAfyCXqDa/MpPpA/HlLq3piHZda
qfAv3dCQmMJqfkG3/3OWrdir4eXvdItlL/zFEZuMoZEicTLsLulLH01b7tJvrZau
qt/SccK9I+THsJQiRlUVO5ZxphKroTielaGAnRn9o2ckFzW53UcdrgTa+NvUpMZb
qXbL2eYKTqsM7/cL79yyWLZWMWUyBaOGxg6UkTIdJMuk4CPB8DAzEH8uTm9XYHAm
f/G88fPVpsyrXCzycZKjCcD9HgNz25Rggxw3h24LmOAvWF83e9tNDfqvUNaA4kdW
Y4TF94AaNB3lESc5ep7hlNVmWFn65bY5C8feGuHqVyM55ETeXGSdCX4kEZvN7+zF
6f+lPIx9WxR/rCmESkKi9lQYh/TLeCvgtRngHh36I3p1udjfJC8rjlDc23dkYK+d
cIg7Gh9g0oPaXbu4FIe3pgtktLQ1jdlJEvs2Z8v4iV5gbhegsZEn8+JyOSFNvfbp
RifJ85pftJJIdjJ4cZX5UKTVpWpfwXoTaTFpOx/pSzmZT03rGen4n83djKDeBAUl
1Tppdh3j0e6JEVnMDYAuY4Z2PROviwm66My5zysYerwZBqyZxyjq80F0WlCkaQcN
zeb+P3EyZk1DqfCGX/1n5Zc8fWg9Nl1SXFgtuUkk/cIdewdmCfY9vfuKBPbXbug3
3Uls3HLU0kE5X9UfUV4o1hlr4EVLU59bXIXGrCutNrOAXjLmFEUDHyzqR8JFdXT5
1tGx3aG+ChDtTzjwGdgiECgypAgTqy4EzkWLSwJgZl7VQa7W/NV5a7t1JTAz5g2K
WCVEEF1zBaac5AOnGUqqtr7ki7i5jS22i+bHayV1L3cjSIOdkVHAiU67EzNfQmwf
mcoGAg7nlZbtgJ9TOMsGLR9oyfqLrC8rckzJW6pCGa6Y4SEKnEOPWhl2UDeCUK0o
G4awR4R/fI3SqvAok8LPeyk52yqdhubbsS/h5aU7fFkWVbJI/ZP+W+HwUO1QbKOw
5JfQoUcWqf8jXeRjSeUSUIHXXYVNtifbQv/rG/zirJf4UDw1AssrgQxIZsip2680
ggjqjj7dTUhlnmWNPFuogKA6SsyOVA7sAaEMSufTpsYuXW1wRLGBeUcQp+AHq4LR
SEFNToIDzh9Pvi5pIheJZlLD+eCqGJJ0oLoioCFqE0yNTwD/c06EC5Q33BD9BFxW
bg0j/iv0aX2MwFYJ5RADSmAzuQTHQBt9ks7xnGx5qu0ck6wJ7RvC3QwbZpNHTtYl
t5ToyPuOXSxgPyMxeBqEAGMl1p04TTF/MKX8HGD5xL4RGrhNlOHP5ZpjzM+RF5Pu
TCoMeOPy1qA2LaXA838NwfqHDy+tZlE2+rv+GqFLuk5/WFeNH+XtZbEZlZs9ppeS
ls6kkUZjZSQ8AsHhnvIIAHfkvquhMs3i2+pGLbjm+ubfKB2UomCj7ew9Cgphi8xb
QG2k3GOD5M6A3oOTSap1DY+PuLbbEl3UpyoeN28h2U98bF53BLYEFceTHQ4ggMO3
rdz94+JqitnG2o9ftGuQHjQNEkDDLvSeLYzxowr5HEK5okZaeCByd94QxtDiM4vs
hWHJTUvh7loXPz0O7b9nR4u1o8tKFzs7zU+mhYYh9j6ZA4UnhyEXIwlQHuZPnv9+
OiFxT77w472oj9eEmh+bSOtiNZ3SIRYT6oE9suXLw6JDQ2bMv/quCySzFMfdK5or
Y8rkS6HcXEjQ6RPuq6WRCLjo3PAK67x+lm83Ks9/GzXwDGa7jTezV7nbW7MzT53R
dNLH9GTINb4AHK48L1IpD6+qRF6U+p3ugvWEfsRaBP1Jj1I9XG6vA4NjcqtVFQWv
ZMW6sXEk4HArA0me4AX16hBFJKASRJZkILxyke8VlTaze+XGTQTsVmDAH9MwDWid
1Jnfo7Jqh3irMXmYFMXuCY1PRbv9Pl+msbSQiNpgdO2OGwOYBl16g8oMxBBiygWn
Sahd79rmsHs0nytuVs27PP+nqypcKjgyl1cXw4RKpXqcGi61jMJ4gwC2ApSi+VaF
YZXEpI1rCLsSEAdvt5ZEXZ4valUW5EwpcmY6oggm6CnzJuEK0xPilGpvG62aMFfM
PqIQETYykbb14I33OguWQkteJBA0/A7aNSY/gTiSendWkKNH3iYLIrz2V0lGxEiJ
IZHlXwPBOF6JvBIFuG08FFdotYfnVWTNwgDncEqYGAZQt8KZru1zQjTtjhp5ZSCl
nI7nEHMQapIbmQv54S8D9QSEqkWOr0GBojxqZnNlCQIwLahm9ZhlMf3QWcacpXKN
cwVTS4/lb1edr6v/eifEi5RMky9tmQ+Y5lAT9/yc3xnT77Ro19ebrFB445pURrSK
niMwuLxDapqknIWdf5Weo8oCfiBW3POp/fy4zfbTFyiovHdXJT/H2c5/89NZ/sPM
oGHqgfcrf5NMhe2hrCj4SH7LxLAV2pIJB+vpyxqP8DQ5ylPc3qRiVKIBei776u6z
Rk6uBdEWIOAKZ5gBkZbjw+DZA1pbIPLvuVNlZyhlFU1y1cRpZjIQhSjdMrzHHv4W
BvJHfFkFZnUmruM/F1iiw4++ivkmKFiNnGimFf908/hvCufSvc+KQmqi6ER0BkO+
qI1CRuKU94gszSb6oAcJz1zliR4fAISpdzH9jZ3MgnxhOfMiQE2s1Fvb4P1KFesx
BMjbpMWJoyLBR3AA1cUiGuWlgdMes/MbQ0HpRJIYNsybtziO3s7+T/kWX3y9c/T0
6Qy2/XE5EuA284FM4YG7FE0mk1wGt+WZmQsZj1aGLV48LMVRc9vuSC+bJQE59iiG
zyNeTxr6TrdWB09IeVSBxjUF/V9+msKZvlSMe0zN3jdxnDv+A0Hnr76ax6svcSA3
2KHnF8iZCSJFPvuCV/8oxRT62OhkFP/+ZsMeVHYe7Zu1CtGtDHQr7zZLz2Ln93EI
XjzT8QdsjAnBpdUwc0NlodNYrCOV01atL7IYMOiiAUfhCJhphTIXtWSvF2Sc90lo
KTsL15x7Q6/aJU5B5vOXZnnhmDM8sEofg0V7jq/6ITOojXethqFhZsfatVriy8Fd
hb+wzRBxCaLlOujYYKMX4UvExlxo2u8NwbGKO0HoKFtKIWoGcdbhOKapW+PLX81e
s4lcgrkuZfGuU7y9EqjFfVsE2KduK69FS/Npj2N55A0bhhVBPWvUgyqUJNZ3IaWG
IJsi+H9KjJlEe7yF7Ud6JnVb+UefdGiC+4axKRCWZR8Z8D0eF4JTgD6QA4wAC9S8
E8+WAaIlxQsHfndiNeVDXO1DSHFCtz3/j9C9+1MMPU+q3h3GNp398A1KQmlQseMA
zGnq7Xjy0dV85b9MJsi/tAzN9afOzMy20N+SOBoL6xl0L8YFGODebj2LhOA9R6kn
LxYIuMkVHvQPGsItgIR3Tp1hjoe5vCnnOkidUxRdlompLD4YtL0OYSqHDAhrP7sa
WeUFQtIEJ59mDyzfqKgCWZNLZNibZLlOY2Z7g4eQ3IIQAfFZZjlpX8umyJ+UD1yi
6hRBqJMXXSyE9wQwvxx9zlpWa8PITYafnpkrVV/r9pEJMke25WpTWO2ChjAaNgfl
0lfabXFl1jzsi4cwu9/L8utPfYVfm8bT8keWjkn5iSMzVAvF/230tTI9kfj5IRlX
SDVGnftknflRGUwMpKwfMJN40bLEq8tW1N8/KaphlNZPCRfc/5RDPb3usy5E3VvJ
GsJOap4hfqXRPIERvUldBMP/eZynMCpSB3Djj1nvBjsHx3N57cpRCD/LaxY3ryDn
H3k9vVXE48dlFoJhFH/W/QC8HxH5rFRl2gBOYSEBpQQy+Bruj5l7I1WwnZ+oaA40
ptGoedRZ4ZvVPs7JZismOutmTgg87GwqTAM2ozN5IwLnnWaKZp3CP0hmOvZX421x
lSVzXZrXZP8GdXqgN52u4YMBV0YHX2t8uid33TICx3RlE+gP0wjDe8e9PKqKVVu/
PX+8g9M99/xh6gmbeicFCICZEbJe/qPH8mqk4Luxe4z4Rv+Fcd2bt/jJo/LUx1Cy
w5i4wDi3P/AzRACV/K2PzUybaLsV8S+Xc9RW9l2bmHNJnHuUAuLuJSOvtCPlAy4Z
vCC1zMIys0W0erGtOGIj8t0N9leyMK8YR64vAIq+1z/JC3zEYRDCNeqJyRRjq0YP
gmpfwjezktJnVvuzzpS83fhYE68H2z56xTSpuRNHY6u0oUua6JUrMPW/2MMqIXNt
j9098JwKpJbkeOem0Waix4qftssB05SVw4gq3SchNAgyFF1NzkvPJRHDyObd+Ng+
2usiuutr4O+i61P3YUz59/ghjx8O0QAQSiZSn3lcKjABC24k8x4BC6i0Y4su376p
iUEuZ65K5h9iXXxuOSTKT3cWv7rQQX3a23U9NqxQ1FmMS/F7FDmxnuQH6xZzb0Uy
xeXnllG/DOloDyN4spzrm31UbQMOjsKSqadr8+j23kaGDfGj7fpHazDy5bt9Lz1C
dCJ1ztB550opTlq6NWHUynN2kqciPkuvAzZDIjBsE8HbeYH0a0ZKUcPLY0gJd07z
oCpmMJZE7+6prkPOoYCG1z05qUxMVNX38kttzbrZv8OJLkSewDw/lYuk7nSFCnMt
OiAmrcxNUbnmbwmxR2H/ZRBlaplUdBQc+0sSeGQ2GOzDtAHaz2LEppXPDMU76myu
dLe6ZCv7bZSdHEkm99zeoUdyya1nOcf++9QtC+lMpzvgOHTZXEJFyD9qHQHIlSBl
czQpxl6mSssoJprxmhXMoLWPNrhH9rt2XZo38xwq7z6QPlPSOmCggOh5JEPawKI7
c3Z4CYnExCRAyq++/anYwTS+way0i8x2X8EXnATXh/Bly1A6tncEmll6jG5rxTjS
8st3150YiC/jSERSuW1LAWG8YaHCEuUx4uBQj9/VCtpYlFDciQ6MkuJhLCHMSPwx
wE1winPx8wffUEQBhtMmTVWwTE0dQwKCJ2ltZQVgTr1LS66xGJ9kxqhloFrHz86b
Sz9fv+REKqmmYJCuUuZk+dGcaYHkIWv6GXtIykrqfTWrkl6pvT8Mkr7OEDa3icbQ
XbaboXcU/Il6ymldIMiQJkYa0n6n+nfuXe2r5pek6Jo4QkkzFsdq/LnliKIEiX5q
y4h3x/LgDxUu7hTI8joizuZN3QI6r4/0l5kAoDHKlL60FXQlbEoAcq+fs4zIWkix
ouv+1qnYmvOU4XgYdJKGfET+GJK8vCdi//4G1anx8CvAiOF2H4HJQMeWCDLRUThg
PbonpuP09EGgITowBAoanMXxbyzOvVw/c3JYPxWRRqGp6HhK/Q0LIrsoWWPEFnF2
1Vw8gJJKppaFMeP58j1VDFMsfiSDi89kq7zV3JcvVMnbHqbzMWjWGaX9gw6I0+D1
jDvmXaSThO3F0LCXOPnDe0AXKm/9i2rpzr9pdO+8h7gHRPDes5n4wv3xmS+8JCvI
+2tmzhamAouzrHfRpieF6JwAp28RNYg7HiSzQsq/JZ+C6qUpmW5OTeLiKNcwg+Rt
ulIemZn2onyl0BnbWdV6rkZF1qNkOUQ3ajFWRCDU1bqagi60SRoBeviErpWX7YPA
L9OZuudCUxW32BzUVlV+cIETz0uYWmYEh2XgJYjRhrJaQ+9wbmX0NQh9kZIn4tIE
rrm374UqEAYgiMQsPOFaOBB6U7XGC+F8wJ4jNQG7m34ooiBAPgCNi8ufKVTzEt6i
1tU7injB5LIpUn/n1kszWHaljKHRLVmPvb2rHliiK3Q9j8YKgHfQhglLQxhLTJOH
rtV7Pas/owS/sU4UcoJcA6HS0GurAXoQizSFpdYuSx1PO8M0mF7tzFiP7dznUPBc
x5CJEPPuvmgZTUkhOF7vRpjzjHH2spMGTv2rJjzPZ7DpyUiUo8U9D7Zx2K6hgHFT
Y7mnq88BX2mbHZN7pSQgio1FmZ86jgY0olXlqKpifBP1Q80Yib+r96IlTbuHztei
YA5u1oPBIS7Msju7TsNHOjwKoRO9lOXHUaTuAMoW22cJm7W7dYbXWjheRAERhK0p
8ndMul7emlptS/OZtqHWqA9pup6D3HRCPrNOT5U0BuinQ9x9uoP5E7LHlB9BESxJ
nIs8eI1yIYw4G9maG/lU7zYiOosWXEMgl2lsPKOqGwLJ7USEuS2EFKadX6paCi94
ROVjryxbRqdZLcP+tLWcRrBPG9Kih0VsNi5pZGRgdVaOLFHs47SjnCgFn8bZWT8X
b3JqvN+R+hIGuuPOOcLGEiHbhsHBobE81koc+qoZ0jkAgoujaK60DSOewKnTae+E
Sm5vOWYGdRsps0Iq16UQypHLGhDmc2HLlTyGB0qoHmg+WFua6T0vtU+HLWEk7DeE
vvGS51PABo2bOVAQ2QPBPrMBqKhEMACX59pjG/+OAFvMhbD6cWL4cmYj+5of+zSe
vK7Lpilx1k55VqIhEiQy6oefUopwRUwJvaJVO5pkNh+7P6ucI2B4Ou48buGxtNTX
7grrvXlO7ueb/lU6Jhl3HYd7f9CRcISufz0VXUGtVc6X5SD+EDDSYTRJcOo0iX9d
WAqYzGKujMyXx0q/Tn9Y3k+WANMFNRcv72qugRVrpfbTesGte1GCMsV8uCfur73C
Kywy5rJfjBdNirt6oEZgJgMC8i92MjL9Sd8OA++S7JapyRq6IEZZEPnoKzKinrHa
1JSZj8CMe59xwqlIqVX7fnio8ryNR10VTJWKmiDDH+YdOUhO0CT/RdGTiLJ7GnfL
eaTvaCIQdHrgDMPqLUmdD5ichDX7xMFaVtZfc6KCcbFFNBLf0djDZ1gFzOIdnlX3
IvRAHa9+KPer206YPE+Kw5ssoK0sdNM7s4k3wcsq26swEuwbxDmCIBjriqvOE24i
Rqv5WYb0U6rGEjODyafzInYchOXX2WYt0osiOnYcg2xPGH8UQHE4AXx8hq75JvJc
tg+BM3Mam4r+MUw6ypv1kqfnjSZO+LJQLpWuRLEpM8L+HTeuJA/9IGrwfP7QkZUv
dqU4m/9Jf14Rh0X+25f5WiqvwOT4UaF3uoKAqR610KqxzoJIE+lgjYeP1BURsbPA
qUtFfkvwNiFQiIM1satvFZqxeKu3yziTFgt0puXk2q0k5GVhZtrWMKPX5MOQGMKx
hXrBgHfZmf2Mmp6Ej//tKo9DFhXc21gY/UKSBQ+eH/F8pzhx7fMzeJPGNkTjziUz
2DKt1MrhAMwmcBO89SqmgbNtECukEjIG7jRYbZqQc8HidRH0ZRlK91ofsV5Was6t
bjJvlA9/i8nGKXCYrL0SWrq3qoaA+JWxuhMqOENS7IMGpr33d8Q8L26kZbodYzm8
F0Pjo2ZiUnMx2YmqEWHYaHC5ohc9t50+xDGzGsyc0y3IOZDoo5DidW0SBZZQFDy6
JWnNQLNrvkP6/XujoK0r1gluAZVHuZ0enHk1yDgQZ5Jqh4aIpDV+84u87Ia+tRpc
+L6Fc/bXVrS5nrNlZrVZjXKia6/j5cR713KPRcr1d9Z6skK7t1YwMsdcggE5fmgP
z0nJNd13UaC4h/QAo0nwcZqiJzwQS2Qef/HY7k8tnb22GrJTDMb+aCGgkaGeKcwL
SOfdSGVYUzETNk9vmZko3FRmvtgD4XqPYtFSDaurpGqgBxoa2Xaq8TFnlqFQOsCK
Ywe7H9D/auTKO8RVvRHwL4/xGUKm8TugYKDtlqBV7svmNgaVCKWS85rcpBgm9TpA
adU4IFaRsACf9Bg8CfsmSWCjvoxZmQn5MMg0MoUbMO+CrMoZ874+1FBvdsc0C8JA
DvO+iZwMu/zKOu6IG+ZdzhLOhj96/DjDOyMMQn+/omh4X9aAdVCz46qB2hdXbgSp
I0b+lSlipioUhqi29FV+mulnKid6L1x0rEp6VIZCDvaRe9sXFte3HDrnJi119WR0
1/uOunDeToAh3DHlrVwuM1VMfnozGqtkcwoJkRXgWm5leBuj5Q0L1oIn6RJF+wWE
dTWgeze/dswi2OoES7Qiedxw783o2XAx5OREIgW9exMZ+kottwD9Pcz06PwUUU+Z
HOaJpLg5YUv+36zGIjuAsMakJwe5YLjenb3VtVwOTHjbH1IbnzBzgO8+DtjlOy5e
hjmfqVo1dASg4rQm0F3cxZDYD7NoKlGLjMmkuMlO9/W4yhmiOrVih5B/nmcLA2hz
bUQZauu+sQBmfHY0hlx+MNK8+q9YQNN8j/uwWEYmul0fPp2KEOsvfRJR4LOlqL8i
/syF9TbiDqmpoo9Q/GC66agMqXb7WrRUjkeS5LiuI3vp+fRXeyfpyFaS+NTpuLTh
CVHu7EUDi2x0g74h8ClEs5KiOBhnaIkseZdPKp7LIx5B8YbF7YPOP6ytJ/4qOGzU
83PusW99W8wYMfJ4kKucgiL9jmRrBLbHj51/E8rzBzrzQTmgdKZBzULpYo0fCd8Q
YyUv9B1KL3EF5RfYdKx3dXGf+qfgbo6T0K/lRpcwUUsZY0764AbqwXGdVngnz3KN
mAX59FSs9xNoD8n2AuEZkDemS881ya5oDViM5dK43w0eLUcQlkjV070v4h8YZhKz
xO6mVu7kJW7tPeQogiji7NuENlM4NhScxcPDXhgvtT0szMTeTvD1WL+YyBUtX2eG
MuNeztcHKwWQZcWWICY/s4JFe4/aTHeWv2wLAvJzFVrZZTCJ5qFJHEXaUXM+Azj5
KDKLZRGW2Ngm0O7Ern3iXiox4P6/nhFfqXVWVzLSlRgIprnTABWpa4eQoE1ya6k2
6Iij/bGRxDyaZaDsS/yEvk084Cm64H+s/cQ2qy9Z7WnJkt4cXiKwzwOU3tNSxqzs
nioAztcdPbS8k+v2SuaruluYK2yYpze2W3RifZrOOr+/L+b7hJc9njq1r4WBt85f
eFFMMhVgfWTSkvxXiQqWZby6uEkOcrWlpk5i2ZOI+cYCjpyALSorWNrOuidyXc/2
hEmW3Y0l+kObsSjm1CdfSYwgyDOtWgT8l7n9iKRL43qyxaKVU8b1Zx35883/jUGt
Azo2IRFuh7LnrywWwis4VbMYVIY+rmFlJyTc0/IBMynokht+9fvV+EXrsjtFGQfg
nria1YWdzLhltKv9ppE++4JYSOkJVw1KcLabOxy80ba6/dNkmgc5wgcbC/n2ERcJ
5vcZoGy1b4/w6ENTUY+JDZjRIZZWe7X3Rx3EYQAlX5ibAyViXYhYXwfTzWByMrAk
5h3F0637/k7TLNG8R0YWjVl0tPR6U725IniUqjRE77Ckuj3QlhCfmmW3uNDBnsFk
0hJ2MPkQBDRlZBx7cHdD/G0YPlgZ+dtmCndwarsfj8hi3tSv8UsRsVAs5NDwssDZ
yKZim1UnR0de9Y9LMFrL1qSMP7xe6EtPJa6uO2XbdzvpDLN6pl3ns6QUlUH+f+4o
CnT8//LT4rrPZN7mIV0yvx9zZOx5FYJU6u6VAtw+hWQCPQJAA/yw1Dp/tuioywfs
+7J3I2VDlIX5PXT88BaP7zMYISehhihfDiXP/u7E33gnV1ic0TiWBivHEoQe6isE
NO3+iZRf/CKyAONH07YzGjvx5ejEOAXppqsxsdINlBiOGgonvwVDpjWD7d6taCq9
1kPQ3F/jfV/uDKbDu/Tdn/0B1q3eccEK0CzQPnd3o7y29S/RGk74ajfczGQlUsCI
1AbYQty7PpevsCb3CFb+f68U0IDmxKZY+zB/RUiPXRLOlAUDNaLfE3Ccyz1KiXcD
8eAId4Ra0wbndTNQ0XUBeA==
`protect END_PROTECTED
