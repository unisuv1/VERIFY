`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
QiAnCw66vb4rrWMsvVytnJ+P3NL3Cn2zIbftQyzUgb0a6GFfBjJlLGkVq0+5A6lW
MjOLKqdwAbUwFVCb4H0JlyaWAtijQ+WDUh3N0tDojzHFO4BeaL7XuSMjqX7W6rOD
E0GYGeQDtXlTCmMRQaB3qedo4PZzAsQl1AAIN8c5iMH05AEjsOXQQjAqNRuVCSyM
1NXttbT1gBNb+dLmuP3rwAuQ1N6A5oFG7oV3rHAzru3xGp17ya96t9II7ILf3NIF
W8nLMh+aGksfgJt+Oznd/xx8a2SYttmuqTMdpFFTaNNzF1ryu1KH66qGoOEgBcgi
HlnKsovJiiGLyaLAZzShQ1YS7tuDTFAu8LU0Ok4ac13sC2od1VoVDHnfbxD0veG/
FRKql6g6x8qob7FBsK0W//b4q4aMjMq2llQ6nx+gXWuirscZiBE/+tpLk/AMHdZv
fPcvMdzbN20OvQ27czGBRR/hhzHTKj46/+5nbKYt16Tm3dfACjz+0L9p0X5NKJrB
2WJ54KpzLxCiKIdVuZByTt1A3ZKo7XpsTPRxC0XtdmB7zH+Gf/+l2YhCjQlzayD0
QkiTu1B2nVCWcGFXRmGelxYnbnJ2UD5FD+0MNRYKzwPr/fgd3mnU5sZ+LpQhqoK1
tj+Muq+C+6re2CuDDK7q1GB6axFyiBfpXAw7iyry9QBw0+JsZ+857RCbVzYHHwgv
V5HgsqQWeYxvV00kgIBM89N/zQD/z46r1FW/lMMybnm2jcRoMhMWCgqq6OmHUd1U
GsFVX3tPdgfoVgCcpEqf2NXU5UZ68t9ViUYnNVm3wgNfvizeh5la+6iiHHDDyWe9
ZidCqfw3zmwPykXmNEydKg+TWll7d/ekk5FpTLnXjKRbWdZszyrHqTQ9jivjM37J
JDtzCwrvg35Lh/nxiDqIPCXzg7VtWOpR2P2jks8kB9cQ3mVIJa1rE6HlKahlKi4s
KCkteMJNGE3ogqH8oI/8BLCkdh65K2E8IrBN9s1HJnkUrMlRuly9oy8Y4I40Bg2j
3hy2nmXp4JFA6aPsxIa9IewTkUiXRvZK72DXNnr4dc+wT48oGQIEMxEKOXC8HKOE
6SLL59HXfi+NTyT8Lr4hAnrGlqletd0o19bJDMWHn/EjprakrBYY7IZa+lc9Faz6
SZC9uopgGJpOahHfleKdd3g3A1fkhRaf+Aa2Ax3EihJqgCBwtp0dxFL10OzC+/jN
xuzGq9k+dPlW1Mbff+cZ4g8TL6BsQxLjDm6cR6PGjo1G2kPJYxDha9CHRDxX6lNr
AmiRRDgQv6E2DBFH7QZGre9vO6v1SFrQ8hhleJ2ZQjT/Ur2aDjA0/n0K1XHYrKFK
yd6Bk9vnb8p/nL5kb+CUxyqZXz5a563rKfWd1X5JxOBstlRTMkWEHJUqRPvCIw+/
IoHNY1ECgQIRrCVA0+wBS69F6fV84Z3TtEZ1GfjJ79/M72HvfzH+7UicbZcm1iYR
GNF4sMtv9/GFjprMyt1M4zFJEaYWIdWHvowN0jGH+txCgHIv8SOyrYKVAsB+UP5Q
+s2DrRcWGHJLz1gL3Kz4Prir/jNDkYFTgJS6jGgNeBZFjg4m7HO1cOfHFJuH/jhd
3o1mtQ7LSJkrbULTNDYLsEycl4zfZeMNhhgdRW4p5XKg5Lo2hT67LKEGR9R0POTd
nc6rOVMikiQSrbPEpp8VYGGjoaUj25GgBAPlZAjDjgE9u69eHDsN1Gswn5woJMYu
hx0hvVWFkCA9pSOsqS7x7DoatEcEi4gxjQ21cNvdMsJsOyhKgoeUmrmGpuxriw86
NeRh+nCcSBAAWvEv4zozIc4nv+R0bMca/EJcrdkMtJjxwlEyzk7QuLGu8v6xD3gX
ltsypS5ETeAQPu5yIfb2FlahMsHEJ7bxux7cLpj2xOAnwtk7NxXAvPY8Pw4DOQYM
v6CXPFceZdaFHLG0fVrw/pmtZ7zUh17Fi32mjNzf7Bog0xF4wY2mPWGwXNLzH6uH
dkzLl3OlcWKbwHQCkw1HHiBsoMZg7bcopdBwrdAClh5T6lGmmnjVKilcdF9KTj/C
QmMHmR9qDpkw28v4Kkiqxpjz3v/X94MjqdqUW2UztPYD4W5SMp9gt+Gd2d2Z3uiq
SnVmnfJwnLV5mRVbxlvUps6C8/K048DPKb0U3OYODpDuT/P+mogF8SX/alggsRFo
hiRnfi8YmZ7df6a3rfU/9kfz2ERdyaVgKwiP+Z+y0n07w5h4HpAViF79KC/ngR65
93b0Ii7WVaV1fj1FdPqyL1J+x3lIPPXV04OePGVwLypjPJbY0zlrMsuFbYznXkOo
GFhQP4tJNHsJ31gF7TQ0N7wgaPzMfhNRpKH4Hrfgs7swS/cN2QyjcoIWX+pxQASY
0CG8y8ljC3S9AQpd7SxGwjhT/qdmiv9kOQixv6cyoYeVWcjP94vYzRhEx6z4M0Rh
8bq2VtWuLxxoNWfRIAntFehk1/OJDcntMWAr0TDfRBUVmB0Xy0NCU9qQ0LenS4iK
V1qq3U5Wetfwv7ev1OTU5Ct9Vrm+cNi1SzSdUDaH9uVM5kie4H+BuMCPihAc52wR
bHIqJtBp1VTk+38q43MIm11sETopMNlVix3ndpGFqxRyfJr2q2PmIYEW0V93EjPo
QqFLBj6vxENFSg6QiwevRUQYFxhFDbrgH+3AyY+onYWm2b2NXERINWMdFJpXleL9
+TQPjo8Hi6QbOEZ8282OvYcw36VdZWL/KyEkLm3TiNBC86VKwx4KL91e8rtTgmRk
AQMXTPaZ9VqlCf+MoVbD3pmD717Zw4QFR/TepbhxkSCZnYGm9mWsvWqbR8uSFD+H
71tJb5vARlGujDZt1DqDTmMXNoI81XYh3nNnvN4wHGowaxW+oy9dc/vCPwC8lE7q
8EreWjUT7GaofpNO6VM/1W8COwhiO0CSyHHY+d9Vqjd5PHIzWNRFRDA/GXNVa0Ak
nQ1yEZOCrJRccLMhZpYTaYStu2FrFHy39aVQUjNykmLsLkP0tJgys4dlHA4OslC6
sAtEYps62XBLt7zt/BajkCyhE4a40X0GKgT24sVWV4avNaX0AsQVyixc4AgfQgN1
OYqFtjYXJpolzl6reMxZ07dRtEUHbT/vZjFENA2eu38gq9i1CW03trLJaqLGs1A6
csTQNW1OnhA4jsgN/0prawdJHxEKsukkKZ3veaPgj9mWe2L0JX4lmJKaSrMTIelq
NDSt2eccE1ynD3eGMUbNfrq9mGgHL8n0n3w/M8ihdnwpdmkdVgb9TBythgyv8oyi
xpDTPhLTVkDCfYraRDQkCKPiRYoH8KR74RrLqOC5lZ5Frb0hT1SnM2i/mq9eRlh4
HgYUL8ltd/hyRKj9/JTSi75tD0ri17mPtemrGMWGLMy5AVOa7icTr5/YX7vQs7Ts
2DWu7w29Bjj+otJZXnlsg0PbMSvO5XND5+/j19T+mv8OoxYEOCeBsWolXspUmCNh
h58uL0CwtyrQ6F9eydlKql6P7SendBmtYReW1NX3dNE+S2kXgFZ36WavzwPibCPU
G5jauy/aNcF5WfYU+HaIJ4o5ywQ/v1z27MjxCqlM63WxCG3Ou4Ok9LisAgl9vC44
H9awaIxdU3ZcX4Zto3oaqnZlCtuvfAy6WRHPdvByyBYY/dEwVsdkyl0V2Fy0pM62
e52vtpwN+p4afISEeXDHgUjHd+MRUdH8cS/Pw73CNHz+JomXxXP5dHkREEkwgllc
V+q2X4WmcegvoIJT2Dkox6zVSowjejTJFPOSCWlo4v1ix7PdTrcxwTpvqFTXz3aU
IcIbu9OVxv7Vy4+gqJT+NYdpzK/+EyxJNYMqC+/xGVZRUo0qgyq51QsUOIlnoLRh
xlHBLg/qNxc6R6Y9pylpTol7PXOzESpmrrqb0tkioplv5naxHpohphzoWLE9+FGa
iZqGbtflIQzreB4FCmAUobtAMMsN/OD9ueseagL8AYdmUFQtHGZjNp6d40twVoY/
D3siqjH69m7eH2SGS8ARmQHfnrYoUFfIJ+56pNLMQxerjKgbaMtjaHSN4IW0M4Vt
hTQQmokfFBTZb6Qiw13MZhsgrLD5zaTG4X6ouPA2O4lvfSsEjAEWFMMI4fqAVlG5
mwWUzhRSJ9408s8BIU/iorYF1hF0WGiNOSYxx2ilAMcE+rwGspMtlwbAwgHsdxQU
Ugt7+EXnz3HVSyfK16/kt/rLIHEPwbhTAQ3SzMljRE+JwPT8h+os2QNRVw0lgT8l
3Ghf9dA/D7O5iIog+ZVz6dAnZIJFgJTO434fra7yIQ4BEoixvKr6Bg0xzBToFRzr
wbM2AetPrP8UP1d9UEwxMBXGBbxVvyK7/PvtMb5/wZWkiZ2jnOHUbO6uONsfR8+/
aECHMz9t7Bh/72v9IFGxFpGf3DRmeTsolCVBaUsk7VWqI+1zK3db8B/1fTjuOabp
/gEPCZkhutvdD3P/n24427obyD/neTVlEE3kTc0OE1tiKn/CpZRald4gO9h42TYT
MX9CCdQ7IDqYjlFS1EVpQX6U6lAfBhs/XHMt3GCHSKOHGp40/5IviK3WTclLIvKY
aUbzEsVa+DkQ6l3dpxw8E5cGaYMTo6pdCzJ68nyBxlk5wainAAKwh7apy5o+nPi9
zV74PdYAVidCVcaTIJ1hFF3XSOu/1kUzBhP8rLuebj2JUkbe11pi6v/AtT4LTswo
c2M6c18wzw6sMA3+eijiZUoewQJrvHIovBJ+bnyyA1LMWK87n62pOIserbrDGYVM
nOsKoehVGtRtGtU+SNsJn0kEBeEy1xkncA6fQVv4KIYpfmEHsBAOcZeMPBmlOutE
Woo3tQ5RNKQ8b+/LYbzIgtz7h9dyx7wfvvJQdQgqjQ4Rr7hjDIbMb64OACEBresP
9drvaQxyOm1TUf26kiUUSv0FQQu4/EMg/ByRVponJw1BxaJF0CsNWvxY5yIznzT2
zCJsupL7y6vU5qshs7zXsxPGwWClddxPrp6/aimI84DANTc100aU7UAjRAdrxLaU
eYj3pbYHUc5bFpcS2wNehaYqTNTAkhDTWzFOKQimf/Y1roDo8XgB5YNiR00QtEG1
ZsdpG6V6eM5BIafkrDWx8r9dgnq/B5lVgYJ5ELq4UAr7Ab+oycIxQSc82L39khIg
rMa7FB79GBTcpZcGG8ckzR0hZ45eE9UuiRSCPh4RRAcGRy96p9KBC9hQRwP2Y0hh
HlCsIiS/MTDR6iVWBEZNwUXRBJGkbs4CWVYRaYMI9ZJ47emfnmZuJRUtfa+8uP9G
5ZJq+UaJHJnbIgta5RslSv2ZELki0RRnigISR4O3eGPbI4vPtClYWdfj7q7eKQlU
fhOkHmufR3Tv6iJkHpU/uHzYEWvWYxAnpBv384Q1rT21ERaq24f1AUMHCN8843Rc
4UgaDheROfiwn1n7MFhSu278Iu/YTNhck1f+9lM0Cr+98xgHbclaBRTxubB5s3x7
wCL+ihPrPsAWL+khgPh76n3qFuNFF2OxBaF0dnf+ZGhiH3e3FVxs2umxASBtCY0W
hf2+Ml8IVZSf3m5CXrhFcQ98zqOcS3flSR9PG72oEK9mxsXYDk6/cfj6bxcZH5BO
idHHZcls4SnWz2XhGJxNpaI4XW9LGrrbqGbALAh82H3/ujwO/rWraZgMSENHlgKc
wg/wdXA6d5YB/9Jv8xDTzFTKWraH+YJvguXC/BT+xL+MY6XXVEV7w7hQQnQl6SqC
kpt+45cssNnfipfngEFT1ugZWRCc33zOdl7CGyNm4sXlPq5zg3ziVGw/Oq+yynO4
PEMij2Cch7atm2qHHC+b0oguPFUjxwi7cTTveaOrL+uQ0K/Ccr4P2Jlptj4RVZbk
vX1u3wnirB9ANUYbXjrf8TBPrlfiYIvTDmM+D7V1so2xiChb9oGDT086BzoK2JN7
4nZVi/wlqOjFAwo1D/Gf65+EjwnWkUcg98J6vyhvxkB/CnA8Eluly6iOD9I9uys7
aghQmlzA3LpLmguqEsg1cn5uFEDfZ+srwxu8pSVXLY/dkG0nEMpfmcw9qmk4IeHq
NWGC8HpfT2x8u1MOnhQv55CN81N56Ues7FNNRnJBn4y0kEgadctQGcS4+EgS2Gvr
53fewFzVnrZpbv+R0h5MpjjcenImzzbrEVpgvyKzY7VWwQAAGJGb0ZgNybHrNT3a
WoPTPclrNXuAPD25p+Sd5lZvL4Cp+e7jemU/DIcruD0wXEWGtXNTfuajQkjSe7bs
dTE0Zdj0Rki9QyAUaFDSllKc0LHIFDpD+HeHnQ3HUHrn0qkBpy3uzf1m6GhHwBJC
STKrX236UH/gDu8AIKi6Te3quhX/ZcxKdlOzG/xQFkPK4gYjeUrplbdnLXmk3N2x
CvWnhDGyS8aJb4qe6Vw6t2a3xuixzXOfdSUFtTIhBWAKXbDH7SMct4y9n9PonLpa
S63dzAS+3U5rO/kM5vJd9K7AmEowLTSmD2bz5lY0KXqIKK6F4+2RJ9kwA4lgAzq9
4E2/ERTuXIjXUkkDSy5eqTUoq81y+BQY4s8JjPLysvS8Wdu6iGxshmevEihUaACN
PpD9aehBgKxHAtdxiaF7nhsBWkAk9NFZZwlfUDT4PAE0G479cvF8eKDD3whjxAJR
k75AvqCn/Jkbb199zriMWzr+9lbZCPpEZXIAwd4+NTxWAcYCrUidKbwUoLgB6Aug
b7adeFgTdjiHglP09Fm1lyJ9UtjWeBJ4VQMAn33IkVc2AePvSUOE7uTNaXRr11a8
47CU0J9Ih+SXsakZAW7daJsPILGC7objOZMKn0gDuTaRBGbmJjcWOB7lj29EfKNG
Gm7DizhDI2katuVMeAAschvZ/XaAfocUIrcod6ewmN0xX+s0jX9Bj+4Msu1s3uRv
D/jEjyGM48urWVILgHHqrL61gK5mfp8ZB6T4+Pv44L97D9KhHNSgJpCF81fviDON
lyUX2P3P6PswrqPBnRMaFrPK6T+WgPRPHzdnlqnSTkohLvrazpzj/knP7+arB2JE
YG+/wyFrgnegnfEDFpDT3yXfXeeXUlEsXjtwDPIvUKYBmK5ju9tg9qbKj34O+dBB
VZm6zwb9gAAU1AA7V6ML95ZMP6frVWqeKk127J2adN8Bqbcd2qOu/iBMXiLqhygy
Iq7Z+b5sqcYuy07td4nwRs+hUvTn3tjyhkRADVt9G9fVWmDXygGaM5EBDXPmu3X+
fr8odbU32kREQU2/M6h/oBuHgW9BbwfpLyWtvPUuK2SRMFvPRenl4yp/459mubFq
fE8Wdu0UtjjDOh7twsjI9pkrab65lJpzxtS9pOGywDV/MPvs30sP5wwvGg1N42Fq
ekRIaXxtQVVlQK9wHGM8wQ==
`protect END_PROTECTED
