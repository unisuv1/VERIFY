`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mifuenn3fvz8zroQlVzTPJkGvsvLQctA1nEA0Bo8Ubd9VQcsSx+L0ZGweB5icm0u
FAMLtU3WiBIB9lLSP8RMQlTzVoZy6f7MGxevUCug3OtXEo9J/4aaYJvSHHuP71nA
lOWW5+9WiJK9z2MkShKvaC2nBbVZaJE86qvHjb/W7swPTZsI/ST08HFKJHO5iV6M
uzBTBJwwmIx7SGUSrMWBDjLQA1ORGA+N+m0voE3+EuCJT8ju31IlQ05R4jN3+1fG
Lr5oYdNj+9HAukpt7+BTK7FZdQ3X4nPc7yxiBZanp4FdlPF1X8SKU5ljTkL7rfM3
WRzMoStWj2CTzLNyoVkngm3XAZqEnAOI0kljhnZoGiS7Dl5D2bPSX5bmHIyRmIou
ugrfhcG8XnZ7Gymg91lXV1rY0JQ8It2d7Dg5thaw7QT+ohTXQRub3/csVAfZ18zQ
oTN1F/eXj7nidavlTRBs3xm4rVnUz7S2B3dCFDsW6HKsC+FAU3g+AWcdFgGJ6Nnn
kKtpz1mCsMLdWZ60EomUlhRyZdAECfRfECvm/bvCZKrbh7HQbaGfO05ybYfI0qGr
3XyeL8FjpARUxtV9e1UmCIi6eDtfrFNegVjGzEnG3T9IplI82M1Z/lCWhvakTNTZ
LL3eZKuIXeiV787SQxYRWZhDOe/EI1KJy+k4uTFdnhwliR5+n4gLUyA8fWBgL7DC
14y7g6mNtbJMUdOKV9bxriaPBbZbpjbYxelb3u7NkhhzZHt0UXayPQwI6YYmZLn7
ebhRfzUKKNr1UGlth54DNc17IbiBqqir1vZVwswmhius0kJ43LlNzP6d3qxcubJ2
nqmb8f1msyNd+TYemCylhZxwiAQuiT3LpUBZNiTKoAQXuIxXeS45ALzrwqU7wfwu
wg0v6Z7hFtyANARW4XlqSWtPXotlFfIcyzGGhDrVXGS3XZpnfmZ4Uun9R3zHFz2b
WnadLWh9zaAfUEQQf2rZ9hD1UhdkQllBHbgUgu3MTn0Gl3CVGTmMbKG+cr38c1Kt
RATBxWf3jSOhuzVN5zz1aY/OJvSagX3FxxOlrH4UT8CxFufFYdPoZtePGOoPSC53
w8CT7XidGAlCW+ioLXDk+R4nUS42IduohrCRyF9YZiWm2Dr5p3lHMkhpN6RyOe6Y
NF941x4d+UD+UGCg/b5IvSCPYloYe9xkYCL2n/weO5OdrSCrKIIf81sWYG+Cs2+7
vxnVLSAjnvMhg0ySbVSdWNro1uBlKiKLZeb21XrVDyUF49ymKYrFYOiQN4687UmL
8YZ2Wp4ht/KKhaYWW0UtA2lTEnRogeNKufA1j57zyC6W+FQzixA+1Ypz/EkuKm/z
tw0OBxHB2nix1PMaTRPk2YreJWwRC/mD7Bd5nrh7UgtUrBl0y659Mem4udivR+HU
iih7+oZIa2l3PJ51QaKMOiuunX6mOQXC5b5k5rT7uP19up4cRYVWW+21jUhk4J5J
d533dvFofbLdPxo8ERjCTylJ7OSDSzXI5aEgH9n59ro=
`protect END_PROTECTED
