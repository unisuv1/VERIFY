`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
o141+vqeJEKbrXV5QsFSjBgQQqtYBMqIabTYp0Mg6Llemui0eh5OlVXXjgPXPcuH
tqed8/Yx+41GBSvuxQWRcrlHdRy0Zx/ZkEzYFhCs0qUAB571NtiwE2Us6/s33Fe/
ch4HFf8zSAxOJgU4230ogXNWrbYao+aSkCU6evh/DeHco7LzxucdJESHesBUkBfG
yTJ/GRSX+lNnWf4uCKvTjbmrG24lkxxs3RWdytmYT5KOiX/PgrgeqJLfpE2W3Jvg
/M6xk2JvORogMOnZSNUYngCCbfieowdeAab83NJdBMZKObYkrPHrfBH9Pj6EVfND
c9PUF6tVi0UAIzdQI/N1y97NujamjR34UQqDO8QsfUFayLL47JSRdDeVjnU35+oV
rAMF0pFi5wIIbABxPE5u8NW45COgycrxYWNY40HxkoO13tIokM6PwiFShO9x7LiO
WGmo4zPH0LHLxvJxng1ymUNdhOT9L1gZ1f8t7DRdjCtEmLfBGZc2g96BaR8gk4Mi
r48R+vR/frwjT3/qgbkCbE+IqhHTyZiEuoWJz9qwaSBJYuHetQf/ulHmGrsITyfb
ZoqVx6Q3rEKAucRf2+Z14aNZKtGmv43muszdhTcAiqU90FiDI4DoICjhEiFXj+aF
jw/T2LkigBFC5rdiyFbu5RKc9w8XC5/oZzX/6vlVwUawDpmC01LUOZqWqrkdiefj
fptHBAdI3KrhvV6ayXLNRJb+xiPdtdmvrznqi+qBUVyeD03+dvQ6X21emKRHAFQB
IpJgk/rR9M3wd12Q3lJHFAbjaSnfEVbB46DkqRxTn1fUglFopQfvHoYwuzaPe+Ru
x9w+4p9zPPN5+l6rFfdj+nql0JQB2dKnDiUBMZUAL7Y+k5NrsetlLmVOOf4S7JZX
TIq11tlx48OtAzT3ST/AAj/KBM2Dh5/TgfzqQF51jm5+BsWMIynVUt5VICbDtFf0
pKOUrV1jKxZKPow2eElDyKtt1G/QnegBaA2Kf6lINuLhn7INJI3bwcK+mc8eSzVA
fibASXSIc/D48NPdOxlPkYLjnxuuBw/7GvwLbWCr3zijv0G1dtTzERy0dagF6yMN
gvD0lYCRnODGHbTQn90D7tbUeq9IZmx260+nLcbYQdwxvZ3740Tdhjp52BTE+xPU
QFLZ8ItzXE8Ro2qCtqg23X9CLkBoCn9NMTzxjdczg/evpFFXdr6LzID7dAFRawDP
yXEN4pd1HE17IeAoaSllNzh0kg7zxluB2bnVKdop5xaKmxh1Jq7i8qisE9EqEaPZ
IDN3F9uDCxc9X7NmaGgCyLqpVkd/ereo49xQZpA+KxlN0JX4+r47JOt1S/mLp+Rf
TMnlrQjlMM+umInkSbZVveqvA0nUfYRNbS35J9OHnmr19BM+9A/9S8t9Ct5XCCXd
8Z2YFKR6krQ9AKW9QTn+a6bx4gzqFnbnLMM7oNdu8EbyFp0x+d4Dce7DxiBwFN9r
9XLr9mcABGjwBPDqk3gvj5RAoQbZTflJJoHMTEGXAucPP6C+lcohFHphLyWYPQtE
nKIa0XTPCOOjf7NTwsjYig==
`protect END_PROTECTED
