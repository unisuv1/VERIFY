`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+/xxeaPw6pfQOPVSFW26pFKFaVZxjtIa6cxtNJXiMQOsw31noxO7kyuzsHM9qWPZ
y2cMvuKA96mb5xYlvxk5yxGMBKD+fJo09sRFK8uQo70URh3MzozNjVkJ44ZDjfty
J9WYm6WVVxpTEFHyWcJZKEshZk6RTJM1BdMa4yt5qvy05IRuEr9SZiDHhR3X4Lbw
dV9xjKbpTkg320pSOOhJRN8nyxCmoEI4Gp8ijUstlUZ5CbLRi+tWYwrCDCTOySrT
lkK8PxC3tIv4NisJRgb6pEdTEXsySHzK255ZSrB4ZNbFmpCmOxfotT0CjWluVopX
va5xC07F71e8aCm9xiS2ALeQ2q4cxiNzSRBuAMC9F4a8g4N4Ff5ajJQNXxqpiVs2
Kbx+BCQstskTFegjZD5LJVI6VQifSbpQsaQgIJ03+5MxBmAvuZKh+IXZpz1DIm9L
7SAIu9XHLdAFyi2L9vZv/aPQQ8XvYVcmuVaqwcM9+nbHdc5n80S+qdZupGoCitUU
E2n9AFXELde7hLSw7GGte5Fu8tLdytP6BSUn9rdI8pC51yhqfcztnKDVnQ9scEPj
DowKPtiTvww5NB4sybf6ljoLkEXluX5Nw6qHzK63LWkFTJ1DZAztcQ72zOIjYJlh
i5X7Ka1Y7+2ibhqF1r+vlWnc859LRiRhpEKU0QE2jhPRvjE8vmI3dmNHfppr2xE5
/tqD4JRvrN3zhT9CPiQDtpnKocbg3WlYS7JlUAJwkuhtjybeCKqFe9qyiNF9VL8M
rPIJKPGeWk0guWaVX1AIxVmRW/zZMefB+J3UbIvORsF7qkgd1xFlKGWkDYib2Mku
LI+2kYEDEu9owATSvK27xLSLIiXTqL4WPs19sE+UkElGrQ/0WkWmZsGzCLgt/6Jw
32lmgWfg/M0Vnv53vyitFqwDvJAN5h6jeEptfMQ3fux+4xlW+BA9YlV42bpnveTo
W1f7OBqH6FaDV7f/bAePsJ2POIX4qFox63Ni8OvVekw+n3Cskjx3deEv8U2loIN0
BvFB0fY/jUTyvJDU7ejV4ZFieSlFYCK3j6It4L8x/Te4kuZ46dLNlxxMemFN7M/l
vaTNfpin4OpvByZ6u3YxPaVX9w+HhP3Pt3U+ajZRkM6I8kF8GOzLy2+kGFN2GG1Z
F8DGlFtnPn5FVDeSSjydR84zkfQdIovKRWGNXwkQGQxgWmDIzn6/3yUMZn360OOK
gUNrW7imTApQmCPthPXPGGenFwHNR9if8ltHOc0gAYdwnGjoy6XDUoHHV8MQ4BX1
KbbZpDH7ZJsT7+2BxifKD2ptKgJbA//ujjH7Q9LbZIqfD9jj/nDw8I5hjgIc4B89
vkM4dhMOqGQ7ia52EKjNP5KXQOX7mwztiADtV/m71WQ0Lax//DVtzDaVj2mNGJcX
/nu1Zjpq2IoEzSaewJlJAJGiiS+3FCOQj3nsFfXEB0h/Oi992bUH4R8k9ApNHTiN
+AVsyQ3hhBrIVAi8KP0h4hbLynMAY4TkfjxaKh55Dl3N30QeYTJCNKL5gML1bFhx
a2VGZIUaP3yqofsDJfnJjiLi2yOW3wim/NKubCNBcZsj7fur5FT8Tw/kVDi1YVhJ
fqprUceAE3jfPPWnQnMlErYKetku6Wj/cWe14uV1nWC56A2nLxAR4nTPzoPV7Nnm
Pm9ZS5GLrfPW+ql31ao7GkpdY6wyKjsr+cqho/xhIWfMP0Ioa0ir7uT6CyWDkXn9
xKrGQm+Uoe1+WhvcXXyvidsSAW7VDw0NWUePaQLByTsBcAaMY4fl6BWHxIkbqiR7
POlRrYrJNHDSRixtlKRDUpb9GgHCHk+SfLYHeccpfkeS7Oia5inJ/yTTKpmU+cTj
7fhSnhN/FLBWBJZt1eaL4v+6B2DclWQKPiK/QPQBLJd7YytNQsUZ29TAIgUEeXXC
SU1TxscwcUXXd9VLITBh9h5NfSRWBniibaASh+J+7djVd7lJ4ecxuBQKOAuRYb29
aOUjumesx70MTNmIjt4OOpGnj1shzb0NkmpSFZhShSLnsC4Hah19KKaWDCO3+WRA
YIGjpR0wrME778lfUMN+ndjQ4EGgEQ1Nw5RP5ldwNCAmQkQ3rLmJymXkuaQmDOVz
c89HrSCYIs2zYbVHEnWTL/MW/o9waXhwNsUjCEwdjjLzFTm8GTXW3DXcvc0sgob4
KQJ9bd9gT7RAmCqyZB1FRRndg1k8KbF6Tt12E5H9Rjv/p97YUvBIWHFRBZqeqH60
LKBlzAuZJfNcKFKORXuuw1817m5jP+MTzHV9oHJz/0gs3TqqcjdxqnR9kCfZerhH
0CUQZju5HKPhkSowd9ZwngEnHja8JtUccW/cAWj/v6C4SGWvJn4azAyB5xqCkGba
2fXD5y4pF/VwYvZpEK80kMmeEXpqrNEj5UsvHROQCtNDBQUb/ZHHA7iNXHNe6YN/
tQquBbXboR8k0p26V0IwPvqx+RCgNLh6LmHnymNakf+R0yNygVIr5OCyutT5ROWr
bVvhwxNnQ+aEWqxD+6FC2KFMRXjOmvUEZAGupQUyZOoYD8aJNAjvqNkYHQVzBj3y
ESFTAwO7Fz+tvr+39hx8UF60ZoeTL9DBdgqSaEi+8pd8M0q7FiaVYpCAEWPdSS7L
YUgwMffO8WeNIZWeDixz08S6kN0fli82YFjl43tZPLs8e09GdVeSMtm3x8T7S60i
sSwdSLGfgXQDTYwbkv5vJs6rt8xLUAzfi6l0X3HetF85bh1ib5tXBX60aEQjAssF
dnOLvAOjWGiVjzuNvUVl6+OxNVif70iyvvW+lBLMU5vqyRMpNDwIcDIQvrNcdS0W
RV08NvxAk4tjpNEYh1jkv0Tv4IriXHD+IIZ0FaI5sUwSBciH2Qkf9CUTiX/gTUU6
jxQtXhHswKaLwJfsSztKNg2Rfi5fAOb2bofAX0vFaUyluJNu/+uMa+9rcPtbot25
uFAZCkQu2zr5sieA5sj+C3M7CB0YYBSnFLshlYi5OkWCijw3raQO0HSFWGvMydOE
89yR/atL53YUzRwXj+ckQkCPYtvQrO5VZy7aAjgO/V8XJiodk2WQ+B7MCqmRdtGM
ENsvD/WqFBtSUkOOUN0UEMh+wjjZKTxQZ07oBtuPvjI3uwfirtE0TDNg8SM19J5a
E6XfZlJZ7yCZS0litzZso2//9bLzJwV/ult37XKcla3ew41JOrhhwCUs8AMBKvua
ajEAtQpL7u+qCd4mLwfV4+Bf4zQmo8+8bsQwUQ+ofjkurnhr6AXGOP9zHE68ZobS
zn3XvEZMDrBNz1+k7vvXRW6jZBV8rvG5VU2+hHi2l2Z6+mzXJUhiZA5izITKi2iC
eDzS5qKZ0+07xlMQ1neL964Y4TtHSXYrJRkl4jjXqrTSnW2zvYP/X4Tuizym+K5l
+IyPAil4K0y4LhUFH3et1eXtpAiJ94nY2i1qZAh5C8egiYxZ437bbOBF3H93ZuNZ
O0ZIEbgHp4+wowgKx2vvm8Pn0yBX4Xf6Ux5Q3P6Hmedkxut55LU4KSVqCoZd7Y0D
Xzill6QZ65t3No5Wz6Tw/muuaqurDnqUpsRmRAy/OoRgnA5iqApcSHxkDEaS2djL
7OYIBvH4HQOqx39I8xF0t/u4UAdjv81kIVAOs+dVFtN5WKE4vzK9YE9xZTy6utuF
4OCkTmCJ7MYqw5I6y1CtuuCsUECHA8BDoiEZacpB9joKNSTc7rJek/ZjRfIIVrZ7
pAhZatbO4vDO+KRPG8cdnW79DV4yEmwgk5kCgz+uUuV1lcufgrU4shpw/WPCHrIB
SQ7LVmy4ZugnFs55pbbZ7C1hundUfuo/9NqvI4qwrtfpl5BrRbnFKl7YvfLfdywg
SQwNqeGMsVBqE6M89L3CSsP++SFpKHJ7zPCua7FDvDrUJcBVUx3k4hVXqrCBRaW1
z+42A3NxmS6e1oF6pSom/PvPo7Nuj+HGDSvkKbqT1Nbquc/+hD1dSHlNi7ZNwg8p
wdopevQ6ew5WKSmQ3uAhcOVKx5vr9vQi/ZlHtvcjkzwnrc0PxZU9udGDjwdd8Msj
/nHpIfyOSnUkm1qmBUUUWyhzcYKIHf3JtAlK2Wp3rG2Bs4ap8eZ4CgdZpPN0S9VF
9gK02bV8rYw+ALWf432eqa/qOCE/RdocnxLOpgdr1/fsdZnrIbB9dv4m+AMgpYZM
CKS7di3g/MkZ8Ov+sCxgIPQylgBoMqX1T1hNkHVdWd3KRvtHABbl9VcXEvATKa9M
M6GS56Mtanraaq7tqiC1tfdWDltuVZucolmnHf3j9L6IuoKM4Q36oYhk1Np2Gfdt
CP1zJ72L0KunC+IySdw0SYjr1/b3XmXmiiP5Ngj/EwKTIkjazz1WLf0y5p0nojoO
TQKYjtSxkHIIo7fk6JGipQ==
`protect END_PROTECTED
