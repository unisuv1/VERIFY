`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eVgWPhj2dSbpPzdiRFITfzl+W3rf2qYMMmNie5gn4arqmAx3OAY3BaGav4phAnlg
UooPhI77uLaACP/gx9OYEJDq3n+X4c0X/hDiyDrhPrHY7L9AWHX/meU8Hr9sQ6XA
QzLhsWKN4ITXZa8Ml8xxqnmTQaaEXdfBuHcB0cJAbniAqg6jV0X/8F5q5dcGaT0y
gOup1V1NnINukf3hocPXfiK8rQnWL1nqqS/++XmJdz5qTsvOPIHOu0a3NNJb8i1G
DB00ByHTYzLxVYBfeRh/bqcw/qagUjzDFWlqQ+ihumxU3Gjg8COrcCo3pu4dCniZ
4iDUUBWEqLAsW/mASEU1c1UsG2iBWvX4gtdsU8FlsersmsLP4pcHfM/ivGyKwbFj
w6Ih8Hw9e/vIQs2GMjP7aee/7JR2IekXTaOz7nKXooEBIk1fA7G1qkB+Gzi1cGwu
qQB26B5ouhTCxfeetkhXytnlX7TT6t0WppM3MGggPklot31walnC5WFZDCCbVOhV
ohLRjyjHSWkMTQZqWEWA1VWvSb4r+Rj1re5Sp6kKbhUCs/GP8wWOy4oB+Y99PgA+
7+8MqIDXApV4eqTigk1IAe84pXZiqkO0BzIKmMSV7+Zs9K63vhtlcIN2Nt7ivCL7
5AaAOoKwg6rN1zw9i1qAn6mTaiBYzAAFx6UozOhrC5/MFQrHBjUXMCpmJm4G23tl
zBtuyIIuIqkCceBzlM80nIRSNgs7LPVYCXbmhbr0eCL45+nu+c2+7VebxNxomf76
S+5R7lVrjGIu2UayHATupSyE5t5Xpsr8j1eRzm4u9vSxXD7aUzy2x7Klj3mWNTjL
omO1oNIFh+LIswdpB4PSaQRf5D/sBm0ubGjzQkSlpHVSRXp0BPTiglkeybxMCM/Q
+mRfQsH9P4lb+e4WvXbp111Aa4Lpyl/T5xqOagPPBroPrPp4jDmEuw6bkxRj0o+8
jeml77xv3/Ph7jvz9VGyCNklKQnL03efDqQybAKDOkjv8gfyiFjTHHcpNGNCkhOf
SBA43oVedNoVH3RNZL3Zvmy4qsW8ohfRqIzyj5Fx/MQzFoGTmLySC2ubP/1S3CHA
rdIw4MEHZy6NGEKEhSpxXZsl6zMgFJ3t67ToQJWKf19Xpbx+nYNkcZ84NS+ceeTH
yaE8QMsP2qqQka6coL1PDvxv3l85YJM/YKO76HhN9kJc4awINvyhPao7GgboObRQ
O7O+U9gEwOitPuhhr6cfc6WvVWrZnMbSK950DwfMu/u5Exb/S6kF3XuH+rzwAIIH
fTAsXODOwe1tAAoU0da832T7OLnbzEmTwVl2lxaLnLcBHT/Id26hUbSX6aUosTJt
yf3ozuFdy0FUQqkq+ZItMWjZWH4rCGPG7QWfZZVIqcZR6xTDFQ3Ez825ltxggCwY
2cDeksjDx0JbYrGohrkjbCprYQs2bQTXTZWuY3R8ByHIUM2yBIIzVjzqnUN9pkIf
`protect END_PROTECTED
