`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
y4gU25iTeQlAfRy1okisOhLV4UrUzxxOTDHK67UPqotyiZDErUhxs+Tn26eqitwc
zu02pybwblpom38vL9Y6t4bNSqzaFYqrnX30Vqq6ncIC4letbXw/uAIuGkd2dfdx
AnxkXznjTyw/K1NT+7e0ZmLPZYSxJG1GLnwxTRwvzwx8XEqpkB8pXBWmy0qniw35
tKo2m4QaxlflKqepGihK9zrk/2pYhsoSH2dk23/W2kx+WJ232QqoAY2Xxpda/NrO
0+fwD9OR0FdoipvIqRDYCMO0dfAnNRpBq0WbvgYwg9SHyJ1wXEPxwiPHq3nQzRSs
207EWPun4ialAfobvi+0kZeurVbAKd1UxqWMLulYqHZQ6e3G2XDKDX8DXpbCAwmI
nrXmQ6V1P7XK1l9G0pHN61FdZvKUJ9ieq23AAPdDNJlwR8UcpBTiw+jZ1QEtQnTN
TocEd7zZmKDabBVpq4SxWNIMVlDQ8JlxdjY2OCtq5fi4QU7hsreSmfRhVq3ujzYZ
I6GXC1RvT6O5OOowVxRRdxl9zkNoTT52g1Tx3b+V9racqbYhiMSCT/pMneXS0+9V
6UTvJEEkumP1/43q7gPAYrnqhY1gW6bmA9qgI7Sr2hvMwyA/x5kAXEYdDQaFkLUP
BssFyHBRQGylSVxm3UUJ89p+yy2hyxuzCTJSpbE6INY+C1oZgx9XB/8aNQTpsYra
izhoqMe/4nWiZTyRv3gZbKlRhnGI/T0fDoc1zMJfMjB8gU2vJsmDEKdJyDfB7Ulh
mniqeagsGWJGcFMbozo/xSmRiwwzdzPH7BAnh9r8BDRKbV0WYGy/sNM0xPwJmWJJ
A6CXQMWHeXMVEYWYQ+yG8xSqy8nl4u/MLYHl7CD/MQ51XDLOcp2E8RqXRw0Ntlpk
csOdAT+6IxhxErHOLpTlcTZEXwvHSpYdKFz2zxrgh7wzgpY+NVN1p33Z2kgorZ1X
FtNhRDX0V3yETGSGoq0qrJevQnimMUlkLYA8Cwrz6mBdRhcR/0OlH7JpUUoGXPkh
jEyA4Miq5sDl8CFfM4bOL0IXfNwVTQa9Nf6W74oNpo/b3mP8PIkYhXbrP++cSemQ
tZQkIaKKXpAe05rbun/IAb0P6CpOgJdVnKqe/OaO0DxVOPqz8kjGuzLQue5pzyEd
skT3ybViPydTaD+VVyTSFX45/Zti+ZWod54igOo6HXWUpUpJEQG9aHXzphf52W7s
BChDXk84rhmuMpVCXxaSlsOhmaDCVzTYZRXhR0uERee6Rts0W4DH0qoDLJKMLE4s
hVgqCh4ax2etsiVqGW3sLAj73F925sKLl7xPr2eaNgnm6F22BhM1x895eL4YL4l+
pOc4PuuxBrT3/oALj/dtgvuCHD+LOzumn0nDrw1EAz9OFzssiY8fu9mQ1x4SYm/O
LtozZw6xEEz2ZH1DeW6kcTRHHZzu2W6Rz/LtjWpf+GEpZw2+xdyu2+GtsW5ighe1
sb+YLe5TUwnxBQM+roMAyHEqMOPcStnEMMvtgVUmax+1g3kkQYkaZkCKHJW9ms/U
p3hOmFCRpmobhy/xKiS0H3i8HWikfEfjnobaWAVTAp6O/jYMd1W3+BDEDx3aFEvj
ygzeyhP/4/xpd2WSa01b5KDpsbU+LhRCba8PuOHLO6xGK8nF6Xmr/PdtfeCSmM02
SayBEEsa0GeiJ0dQeqsk7SdGaxBV0lpTxW6e0ktT5nSEszVcy9wbCnJkHVsIZDsC
oiEFe8WIvZ3LAKO+q5SNcROQ6yMHLiF5FVrdpMrIUKcjg/el+uP42LNyLeKCKj+7
PU6Ib1OjjjHHEgvckGWjhUgCR23cQfBBcsWVSL4d2GJi7+SKps6QWncyheKkkV2m
dS4SO3fleyf4epld41QKsaCGvGuCb1pi/YDP8iZscJpanNNwv/dM5B8pTqH+DuGT
FzXIX6SFZNqDI5Oa/DE8Tq9OkbcnsrV0NpeDt22vejkmD9pWI0WwE7PY2lC65azD
dxAPgzUiFIBqNtA6MIy8R4ni0SD0wocak4hbJ4HGnywuOVk8xM72HnkZyOstdtK2
qn4dzgKQlqL0eM0lRJCYF+8WgDsynvoLcaLXgorZ6oVQRAzKULCYdedZG5FOb/+m
huhwuhSIG2P99AaoMCvgzw/7XdsktRGl9MaiYl4ZfkB+XanTW3PK/9TOMphOJd+g
FAvDQREOc0+BiHPHwhQGz3l841nIBv0Kq6p+eDDPJvKIu8endu+W5nBG2tQCq7Oo
90O6pASBdIHb3z02tjuWPUhq9EbX0rYhlApab1XdWI7KR/wgCg5Y202NLKrtd09U
xko7OseV+NraNAjYZ7RJHy84dABU7A5IFBgDc3iXwbKKtmjY532J7o/9YhWj8R1F
ywx2fbyrWy+2FCvgkjO11d2zdcmik3Jfwdg/pIitndNEpkkjzNhdKQo88NImLPxl
Dzmaz4ZURXs7o0wRR2wBsjtEM1lX8DFA7DkP7QBLpI1npwd3AE/UHZ5gzSy7cW4h
Brp+omw/59o99QLpzvWgT71kLMiKewVkCiEw2PPx+5PEsIoq58KYm2PA/SVqZ/mf
QHHBRGgbMOPYd45h97y6WD17p7vsIk4S8mrM8nipzMnUz+gMsx0P9lZ2zDBDp7Vw
3RDqxtpX0ZZsfXT+Bi/lSeoGSEQWwbw4z8LOtPfA1jrNkGTKASMEr0sZzn3i5hwy
abddEMJiXcdJgSfAmjSqAJb9CLbzcoo6ZpCNvkzfgZCWToUhi44tVERcbpgwV33u
61EC1ye4Bn1fKNtCBdRjqxEKjzcKtXHMCZVzba2am8QJWLjwVsAczBxISg/k81IC
0AMGOCVcE4bdzw6xc9gWUKcSNWva0FpxLeJFZxffTflhbhwOHOePlFoloMB+XxC3
Awf+eJwUfntxwCbkrPVpLeYeJJOyDXgRUHuiniLTO8kKaHosXyOTyT5tsAVuqOtE
ig0V8UEB3OJEFYKdYEdwRuwV+65ywwva53wVYzFE+lh7xuADtMLmtRW16J4uxFWk
+KApzXp6JNo8gXngb5UR281cLI0JGzlR2zQhKgZzERj4SsH1c2jN8p9NIOHdUN1t
WBBFOtNwd5w6GCkC+r208IU6OvXVUppwqqeWuZhZwuUSOcBoUYeJjCUrazqj8Usy
+wEQJxIkx0UN0HYSJ1P+ciRfTqVfTEaC8277cs7AmF0pLCKeLlnE8xCy1XjlWPlo
EmruB0dbopj/QZUY4AIEz+d9RnzrFLxPQl9PB+NRW2Has72B7HQvoUPvstsYwa80
H3QMwl2hwM/06bFAV3b+6SOgfFxdjxvF5b2TVvIaT0Q7n9BHjcRa7VMFWaXONU5C
NfOpK1au0PfMnQPFrLZ/vlxC1u6OenfGUFnAWf1F8zArDEO0T9D+UTmjFFvvCt3h
EHPrbCwIWaEhgp9WLO7eRP1DbhwLRXraMISvNAlFAEfe1mPFFi8GTg2BqQqh07o3
k7vr/nLzMmqN0aQsEubUdf9rIFST9IvR3WpFYtpzA71bC1Ipc/3pWTTNUfGlgfEo
GU3Tz/OLe5Bxb1Wv8E3KzFJKBtCKj9nFP1H4J1Re0giCeTOlCCv/84ZEVPPwzTMB
GfovvKSKHYbDc9oMCswVrXLZrFnIa4GKyeaES7PqWtQOoPeDa57KFc5t/bnjoF+M
4xQnQ6J/2ZOsUoIOBRQPsN7AvMqXXbUaosCg+BjuBJnXVwN8I4f1wcxUjnwCxurY
cxItSib/bvTN5wMvp5jnWi9KKxFASIGbcTGi4IKMT5yydK7oxG5+pyJHAU56obk6
I56/qwBNIOKuN65xGNslvQT+VWhpjY5Lnht/iEtT/iLygsP+V0YFQloIs5khKnlV
3yohZgN8rdC9pDjaZrBjrjDfvMPx3Q0OC6SMuWsRF4zl7R9wmdeBMiL2slYeF0+z
GMVn1Qh779iZfJviVL55gpvlnEgRsbbwT2Pvh5jj+pzFzx52k++Nxurl9G3Ywh6r
emGWf6afiqyehm4QEa5aoOsvZ0gq3DVs3qqp0L3yXgkd3vTWYrzIgx9N99mS9VKv
ovuxiRBzEFeK2tmQj/b/TeoOmkNEIIPmXdFBOrfKg/UbzGP93K1Lxf1GLw9vp4zY
PrXKj9U4FPuj918jyBr+hKJxWqKA85J3sAbNSSDbiC8vyOdiQ9GvJTmbMQcf5c91
ZoEY1wVVmbi9Dz8RcqKQsydEkwXLZNptkwUJaQSiudWB5YaMhClNxh1eCJeiMzbN
zWLWTWYxJwQPFN/nyq5gEfZrP6gdrvCW9YGfTRwoAFhcBlP7msvmjt3qjViW+1By
XIZtBlghIidfBjquQiv5nKz+Vv0CJyLfsYqKpjJVAiveKU2vISR6rutqEnWNgGzV
3bvSrO6CNN1NY/Oux5PFWHPbf5FSo0onk6xHSm74KmTBG7gE+5fh3Xw2gtn/rycX
RhrrUm3K0plSSAAVbbOtLmGgxHZjODjQvNqU5NRP+ZE0nZiy99WTHoQvVNW6FFsc
KLYqJOB/nbRV//ScZJyf2PQmakFb4PoCMPTPNLzEbtQdDO8PVMa/xRHbqj9SGTyV
a3fWes73K0SyRtcM2VqsYiQp5OE/n3Dg97PVJtxwX2QptITbnDbOMaxOj1jVRrLm
mSeHl6FioHcx5ZFL62JzM30Cr4ISBLUDn8sekBfDKIFTjyCVmOEnLs3tHLx0rjLV
1HaePxqzHwnt9/KqC3rdUGPRTqpwmvNpB6j5RUFgmqmuLrJL687Vc/ax0RAyF6GM
EwvNiQs1c8MoowtW7DSJmzBKWBOEFpjx5XjMxfEWaE7hWgzmy/0oZSBOc907RK1N
MpxHZyJ95Y6m8s5/pbVPt4jFw/rVp9A/EfBfK/2QcZlTOVrv6qMtgbZm85xTkOQu
gTwdAIenizP3qL/q9X0R64FNgk+FAhKxZPdhZ4pVGVTNtph7pcyfRsmdn1XZlJFo
0y8JiTrbJKZLNPUR3Gbke8Z+tGhxt4C5E92MjJmAJKcWqzUg8H6PiYYCqjbof0Sr
/SLIXgGYaiZ0IIjovWhL9OheU2rsXNHDS31LTwgh2rvgwyXBGRa6fMIrfXeF9Q1P
Eg8VV3zwcakHhXu2T5BgM9vys8GZJD4B/ERPSX+uNfJy7gDEIB7KMsdtrsaozdDn
qU6gb7+C/wFXn7q9tJdlLccuKXW9LldWuW3qlSbMETSDaMS1Rr1vc3Y/NW22aleC
eTnw9VE6oReQONSV8/CmkVxrfVI2qSK5qBl6zlhZFQThSz+XRaGjPQzDpna0zZk5
7oDnY+c3nWbajtskZsL/6jswwkXYLRCWcNCdGacMbG627fG7z+2fsM7dT3q/w8pz
9054PRbRO+sohh9t0xeLkkOMN1XUaTxaZ2CN7b6jym0noLafMQxNVfDVL8Bxm72q
m2d1wVqiRyJ8D6mvTit98FGivtToXPnr83ocmSZyqiX9Ku/05lLYpR6VqQ8PSyBJ
8BRLZfK4dv7lAVhAvZepErmivtAy5UkvG0M87+biaRPKSlESJgY9DuRtVZIuo+hV
KaXJxgTnJs7a0L256cV7fDEJmTPdu3O2sOqPEOdCxrDxufOFDtmuLPw3OB2KGxUU
40dGwjyTIAGyYTdL3cDJ5xlBwEnSAYYmZFYi5NmdxzFMo/CPmrOaM09+EgSuVr2q
Y49k/q4iLS6/Pc2cyGXNUfIOkJoWj9LGWtGLZ6RmS6P7rOEUBZi6Nk1igrGQ+BpB
OLBlMgftLC5j9yfsRDGYEYKDsCnLuMUvaPg8KTk68Fkets1smMmzS3TbLP/Jw1z+
Ux2kljcKHWdrts1B6UD+1N3NcT0qjL1C+NsFnaq6gWgqBW2e7mrU+Ue/0rtbPV6l
SJ6FislLDdw8k5eEj6/MdVLJj7r0vZfuFwCrlv+iiX1Qzr4zfY7sXQl2XTMYpT2D
EWypEiStChXMlCNNWmkgo3jeqM36b5gd+Osnm9OcYxZho7BMF8G6WrjMqrnc8omE
/2Nif9THxATJrPJ/8Zv/NX9dUEMpoq8tC08ku9v0nWOGQFC213PpFsFT8GmKshI7
oYRDxpA2V1GbxDfUnn4TPriLroW9a2WetJrd0bqXWSzqdIB3WMy3IvSOrYul4wRg
6XutdDNL6yWurWpGj6srPtaWA88bj7Cu/i7YY0ZXJ3bBGzcsGADkN5fk2xOp4ls7
hGmGH2WyOi22m+CqzGYrCOqdAx77fWF6483oWPpedMJ92cN2rVPw8yx9VJVJOs46
00mg0Q0lNKd+WHGvpkyGecieyXMggWq8YYc1SNNnRj+Z9sjxAbWHHi1U4XbzI3/P
6n/u25Gyo1OvZfMef7eoCbohTMHCYrx4g571orKoq9RSKbbQ3N+mSaQd2TneBkdk
YJ8umkvaw2y/dz6bzVaITad4yOyA4lrp8DQiZ6sxu66VcdIbC6N4GCPVGAFTwKPw
DMVAMoAMlEdiAYOL1WvRpQJP4fbCiKuf8JRfFTUIgy1BGYZOc/ritHKA9o//0CiM
CoFMwbpmj8AHUZMFjWoBYtUQA0QKmCsxa2g9RLvWXugo5iUdTL5JKHcUlox7pdbe
OsH8CE8jeRSWjAND3HKCDrNUYmeCNRZ6bOFb8xor3ba5lB+fa8kdOJYdfjUt2Xs7
TItMdH8s+kvRYvhvtlB/ndl67GIQGN1BIxPiyLX3w/DotMWTU3XgiTuV7+PnMUwB
x0i16ZdJCB6s+1nBTucaYskX4jGHBljzvIs66h1QUs72BjKHt4BHH+NxroK3xG0b
x1WME2AXJKoNmZMUlrvsZjBTaLwfXZBmH/b+AvTqstmppGkv0BJn4DVkTG/J+sB0
mEMcRxQB/hZ8tmMH5LiF0OstpMGV3dFbESFBZP/f9a2Pjndm8/QbGFS5TTY2In9V
IT348vQ9gG/Ru8/EwhIGLxKtp6LsgenvxSSmeDw5d3JckmWNpSi4TM4mf0sNzpTJ
UpsFtHiSdZN8up20xAzHus1UcPDFipmp7h62vnc66gM5cwusXlwnJiEblW4M74Nu
O0SSeK7g8xZo3Z0hHnMm3iOo0nPVjESKIKCGb9K9cp3oJv+s5M9MY8qYYvZPfDtQ
G+h0SRNOsTh0X+Xumcjh+PuK7w4FKIyJ9GB7kJK04dm5fRbVCXI0gda6yretpLkN
gU8CQg8lru5/LQamvmid+0yspF+eELz7G4EVUy6ky5HTE96Z1Q1xvpwFELPAbRn8
fUgc5v+z7FB/Ct3qAEA1hosnxhlcGG91PHQfCVzt8jhcQV+dvhQJmeixMzGmQqp6
kJEDXaIrJ5q98HqP1JKpZetxTWGnzEwEj0PnyI0rqYp1msu7ND+jDEaNSjHkDfFF
xVep15ERoXHfUZe8NArInbL+OZxpSn0dqK4zMNDEMOuKcjCZKtFVMmAWFFJh4+MX
LuU/Wj/xmClMGTKdqbmZMWF9bch47bKp3jEGfLzoV3qMxL6XW4TVfFtUZCX9uBq3
RHUtAzi+VggrEmvKyPh8k+tmQRI4HN9S5sfbSDj/VuKOfLhDK5BZd2HKGN/y1xCy
IkMpbIOlpEYemPeDfCuSIzX3Ht3Erm+rsZLvIQf5VXiaJzc5i7WAz1t16CYYFK4d
7oUt9w58InIKBZgTVwB/v/i6MxIBApVFE0FJ9c9DvxxXNbJeTCQ7KWAYHdK+UNEg
NJt+X6qKNdIr+V6q6aF3N2K6RaFsrREXL9FRLjBtGZV8NmMBpX0TQykujR7MNzvP
yB0TPySBRsRJIuNEeE+q+b8uiqLspUuxBBfp8UaQmo525zePy77H4AiR828tFYZ5
sNO+9bzEvIDQ0oDZZBm4wH2DpBFA+mG3hlvApNRzXSwgXXlCx37/Dzq/AK9lLByL
JkFsbBbxlD09HTxMdBSXm3EcryJmXeOQ7zy77NTHvqnQqO6G3U5CZIDo3rPccCOb
EKOB/nMZyEKOdHq0aoFHk7Y82lJmZ7i8WBI2FflxKl0+uupKJBfWClCJHkPlXFzb
Y+C3E7CXadQ6EIWxsx4bnYbTxBETpxJjQpsOI//+kLBxnTDRC1DgxAi5HUsylIox
b5ZAEtOnbtft1xoCPCizylU8Z/T/wUgxsEbRyVHGgjMR1+fUyE5VFNIrWMOyiYth
A5ZvezgB5RA2FVeehgAzQuXKeoez8wxeGS+1AlcZ4XghxkAee+gKR8ApaxzoxVnd
4k69qJj4dfSg4TWQD79XGe9D89KnTBIqprDLyYetEvSh0b0oj0w7/au98XJq1IXl
C+fd1iXkEcc8Vs6Zv8c3fVLNFGPSpWrIlyJflMOxkkQgl8n2WGtBphYEyd6dN5Pn
btnJ9/1KhG9ZmFDGmIW3wTyOfvfen0qfhfY41KrSBuAz9hHoaBfou1IMpWeGU7Px
9Z8ILEoJ9ifWa8Fq7EoOZJXB4QuC6bgFCVxjvFfwyS8gbJxE7ys6pyHhSGpq18Zb
2Y07JSLguLXS/16SPJI+etfhMfnsDasC/C8BGJEKRnXS9PdzNCejbdBq4gBoyDEm
IyYkdojVX8IDdzEaEaRS35GIK+hVG4deSJ7j1b13Fbd7i1cwExLhDHvY3bkFsVs5
wuV5MZfZcqZyel4o8rfIzV9RJWL42viKr6es8l6lkJg4y8cFxduqmVmVc7HSmUcQ
9Brhu0uOxpPRsS6WvYFh8e3nwsAkkY6qIpd8pMXh+9U6Epi6dzaijS2wPl7MY3Np
G+t/2dKrRMqDFHQgIRC6DhqFfl7YEs5j0TEI7pb/gyCgvYFT6/C53fDgs0quSA5o
TQV0y/Zay3bb5F0gCbHfKBM94CqdecXa8Wj6FOdpiAjQ0vIoncFY8kBBtJhJjm5e
4r7xwTEDThUgT1tj6Vhfm5vJRDlGaGULw8NSi1N3cuFy4wcPA2xpJ/rb7lI+M0Jr
CISZc73Jyb6ctRQvMUIK3+DIZ/ByjhmnWcEKRU1DlqpZu8Yzv0dB5zP/nq+1TeMe
ge3HFCc6J4pLtc6WqZHQhixx+jRFhlr/+kz3qFEFqEx7B79wz12e1IwGXUWVIW5H
xjPO50h/HfOq0R3x7r88ZtaW40tXkdU5+j5ySeqrrNXDjWndVDMGHX7nnEBjg2MG
PFnzydxyYQnTgYOYe2R1BVu5CBPh6XPE03DccZjNpKEHDR+RWpt6G2zRVKX1ssl4
LXWOn3Y6Yp6L4NI8dbeKVCGq0wLOesMSfznBe7501WC5YqrVytQcmpqzAEtJVBCc
vhyQ8M3J3rhD1hAR+li1fAIIfJxNtzyCvPSGmkn64l1VCsZvn+xueIl4mM13HMxk
OLP+o0ccrns4FJI5RPAQJx+U5PAGhatk9cp3h/5eReGPX2Qj9gvGLB/pUqjN1i+e
r1zVH0H2ResdrwMGZ20KcYf+a4Fxt2eo2I7QjBP1JtrD4lhlF2s9tqOl3BXdBktg
4wPGJcdrayRNUM8HsnXylxY+pmbpHXhA4yTxHw//08XqVJIKmehG5dFHqDhJ7sM3
y0pTL/A+WahrS0b9xqkbiqiWNTOkXfPg67a9ggXw1a7BUCvws2cquAB0wos6fT8q
OjMtVhQ2fYiRw16nyc9hnviRWI4jVnrT+X0E8Sj+tMw=
`protect END_PROTECTED
