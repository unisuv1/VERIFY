`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qySqI0wJ88IkRK6aecE4Yd/EZAGUVoSFJ72w1eXU1cobx+EoKo4a4FkXiTZ4x/X4
5tMjKD3wgVzNoDNY2soA8BZLjgGXCqC74KyxPNIKjqTPyZq8aR7nBxir4be1K3Rq
M+q24PHYpjprJdpGwx3L0AIq+BrUfu/EusVc7ervn6PhO6TImxhUPtuA1ouj3CHl
/JeNShHh+R1CaNg4ThIrMTfYW9g3CbzYRwDUcQZNITGNguIEFLBT8siD07//qsix
MsTGEnmoGWSOcexEAxCHq4qEQzMsitsegVm3HkLSmjA3/d5chiibBI8WKw/dXSi2
IzALewLVQ7uUL3hZsFFf42Hql6xRXqlIzJz32jKqwWOwRMQmPtmAJZgAruKVFC9s
96YQi2tFqZiJ50hOZVgaWmTTvxOqDX8OMboyPNrnNkejz2dvokY84XcVetvJOLsv
vkPde3ogM2N4PfMrD+g3rOi/FSeoZFTZ9U/N2HgVzznLkVN/2quh2sBTJCmRPxfz
C8rQ3VhmiJxZ/WZ3nUq7tTJ3Tg4SbNpvmc7ZJ4zJwu8Jm2yKhwnp8y8qEQZj46P7
RwVnawyHfD9HacewCf5N0uXee+eHJpXNPYao1hft33xjthIem7NjOz0MDiOyx6k0
Set0MVcCdvq/zOFhAzIfAPgPi/gAWbvEOiznRSwn6g1C0a5bqTuqGJeEptjq4nDy
O7eItulyBAyrtzCb2uxuSeSQd3gvZuuRmnwxDqP7eq2EI1ybBPWGVZD9u7y44ybB
RtHjrkuNc4/OCoDBmNxU6IhgGqpjJw0Qq5kWdodjVxxt3anrMcL1nQ8Gjx5um4d6
0CCOMmMmlyc53t02l+r9ZUkIITnAw9imlL33HpHvZqV5SKGEvRxzQ3bDJd8hgdVW
CXzzXYqzoTq6s8GAeF/3EtxEn9BauF2KZGMD9i9zJwpdIJg6q+W9bm5/jmA1Xm3d
HJcQntiyqjNft0ZaQkFDLbDy3Iz2ehPLVCMHzUgbdOEJLElBeu/1RcNQ9vlgrwSG
TfhVGeMfaG+etaRUYeVB45vFMHe/YbjIPk1i/nqENiIo0QcDP4IzmewHsxvI9CRY
`protect END_PROTECTED
