`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jC6ynSDwLHwUxy5NcRy/LSxcEknjt2YmGtTL7GgHf+UrcSWas5lxsMj7Xqip4A1P
Wsh+bj1LKoSF4dHeo9trxGybaQ2My9KBmNFrODObkWGfEG40OZLvkU0VoEYS0wZd
FPFqV4ZNWT4iI+tau17KV9BZy5LWvDxAzL0reJ4e3rYeUH0QI8Y55/B2uJKXV+P5
oHWDkoQhyNzspjvgEkghiId+6EieDhv7nJiPjjLNPQ1VRWi504mEXNtCdeMuKJmv
GNdlYZQep9kH6kpxk6KRkkk2h34ELrWGYockd+Gfe+xzLUXscK6Qxe1KkdVrStxY
4/OiYRUBYnHX1pDgGrN5neBidX/Ppjgy7RF0+pHPaE4gOkAsqlQEZoTBKhDqvmzb
tkHNfspPNuvwQbhovb5Jn3IWDtyILYoE4RxBqdY8+DIKT59Gglmm8jbabMISVvPX
7riGOIu2vgIF2rUcSVJ/wlUxAjVCurxPaqzT/W9rbdrtkNtDGBEaDkphZowHs76F
9dxTlM7rVDTMLl+sDMtIJfynEpjUF6ASA198Kx+ZYbrFhBmflT9twi+KPq6oy/J0
fYgcja5GiGUI5lUCFwxzcyVQbnA81B3mNRNhlyqb/9te4hekt8f9NTkYFpNLCTlR
CEDuJok9AxI5UkalEbaYb83axOwARYKCI3B9JJ3mbYLuSJuwgwyjjNgnVGAmKc4Q
RxJAaYIk9YsAMX8iK6ISuGb/VIEGSKWAbh44FbnjoV/mTUvdOORC4GfpN/FvbNBt
qkr/oaWVwi/Znwfm/UBX0YlHoKphrtkXZFYislhZSj95xzSzmIxLa0Od8MCcQnih
WgyL0nTPDFU0gu18DhFPZkMGqVIJCC+OiujQZWkIvKM+xpK67Tm6dkz+u996Iz2p
rAzpglhxEvbbxoCssE1GuZZWg+WfuU6iVN/QnvJd91K9HdGxYMMooIPDzZWFvlMO
Gq4eHnJ/tJYG1rKF3T3X1ts1Pur/e3HNZRdIByx0I2szqlHUabvrQUCRZ5oKfG5J
CLTnJYtdVOXEXgNpLL1FvPTHyAORWl7FwCc7TvjhxqHkjzNSugEHNK8jJ6pqiLuV
fNkCukLvoV2fXSuFLG0Ham8kndKzVvKudlzWrnqHsyjwAxxKAdYiJj9o0Mi6YQHS
uaI9TdcA7dDKJxmx7jPZgSTfdEIKHzO81dOUPGtXvbksOJc3lXhHFQFSEWZqsskJ
eMNgHx+ojz7JkGhVR9EJJSW/GexQg884NJ2ShRRYR09VG4vTG7b7r+4FgaiU0CwI
mnjQw4PTF9wOsubNTUSV9O9aeoI8ig8d0FZEaDvyuLIsb+6WE/7PiJZAO+7wypVq
MhovAdm81Twt63tU+osb8rW8hfJ4fhY0J3esAqdGkXbIF+kfMFdU58qXLIr5vUK9
T7Fc7xCDxC7j00q/sVB4fV8gc5PdhYOT3SHs76MT8JBbPEX18AP5WmpN6+umrp7K
fM41f1GHnElP8CTGwCp+lEegXfV8uF4U/GcWIK0xrEQnugH8m8WjM88kkT7KC9VQ
ZgerTGEr2i71E1tJEBW1m81fr1zvI8e2pvYY0uagMsVOKFKw50it3iQWu7VYq5hQ
IvooLXamY2K4hTDrHizs+CG/6UD081f1pKIIuHDt/EvccP+8iB6WHprraSKC1UWM
t85271/0/NiUtIrtJ2UGZWHIF1Qi4+8uyDngMPoZnfiIu7OqNTLv0COD/3sCBnJ3
mXfCKksoUKLlHGGsFF64VwQKmQH2bmVhdIn/644lsgSCmt+8vEKQ8FMdeEJvfTOu
LHGr1hgcKE/W15e6O0SjrctzwReALvkjjmVeZKeWdJIO84QvMJQfTtv52SXVfvMi
ixI1C/8iOO90DrV2IWa0YvEOg4MTJeFNOcSMQki+uha7n7ZgnKnJr16gO85XfFzW
irfsye6QsOBHJu7wg9AGIqD99oPXevTUfUOGIu4JvVjWexkAzNFw+GBdNWB0oqWl
4+XDbfXhxDsmI/Al0rud1pX4gMxOhMW+I9vxsCx/FhBVFBVt8JUl/QX31+51kX6I
CTQlpV781XXbTnGDxR12Hs7MsMRa6s0g8km8IK7/ubKcFs9mVk3vfoxMpYoqNcIN
Bm9Xy4egk8tT/emyQMKV0kdLLobLvVyAzowUaVBbi72+PAWNAVvidYP9XmQBZQ4Y
w0aU79F21J+9Rg06xAg4jKdioFX+nE/d3M+lFFD+UQhhEWcwnnVNcJGqGzyxUJZh
RKMID61ehibNpS0EFu8bSDxHYzf1tGN1dUuQAqm07L3Yz9j3WGie7ffffJIFmheA
nzgg1iACjJ6KaBwy0iSGlp1elPMU/PB+duxlJ1O0TsgjnGlOXyXIV1rpDuirty5C
QPQI8Ex6+getYNXg8hGycQsLNqQTaCKCjAieKrBx1r+9u3J+gDRjxGq69In+Az5h
3lNhSnpapCOCTgxY1Kne06aYkfmRggZGzdqVjAwG/JlazRAXad8Wng1FhiwbMVPb
n1VcFSqPRlgDQ2M+wVpEpL3SpZ4mdqD0x5RVyo8ZFGPNIU5u98KUkf4WnL248eBQ
R/4HcSG6ixVJ/is8Pv+qG4or3QCsX/HUJ6jRUudirH/WMmc27CFJwdWivYaFbgPR
ptK/vjaIfN7C3sh89rrlJM7crF1Wfv9umkMWy2k6aUHduBxKmNRtCNThi0Fg28+w
tao/staMLXGxOeSDI1A9KZ6ADLajsnyhWZdgCkQDIcrOwu8B6VzT/HlYjUHBt1JV
dm57C8G8HudondXyNNDLl9t3o6ffeFbETqtRMeWkczZRoXNYDUhbvV93tnvZf2Y4
yek6qfIhgMHS9M+qI8McOY39tBMFqiD6HDG5XqPjSx1wvd+jTnF5KrzsvHoTlSQg
yRJfgTK1bNAd/3QOwCKr1P9M3Zz98tMFwbXnSvbfaI8HVlZa6yqgCUtnD7UQ8uNh
GbwR3BOhO8VngBDFfLMLWWOxiHFpqGZkDtDJkuuZ6cLMBjp5QNGSGyhSQxwun8rP
RqkCu30sZ3JXuhZU+RY2eUzh1mys16yNf7Lr2u4XWcJ6ccFxhZ01prbTIO9/uhnN
EKn8Llyxi3tM0lAARfYVufJpv4XSwZS6Z5kWTW5srzsOHQMfaCeSsWwevzRgcy3O
E/pV+UxtMOuHx6Xv9OIoC+iCvy9NkpCuSyBRwKQAVUCIwrMf2Fl6+gFPNdWw7YjN
KZ9MaNVkGwcn9zC7/tqhvwadw/4ySHa+6LA87rO0AbuybzgStB/0IZi7hWi4lLJA
wbEu42Pc6jj5JYy1h/sl9BKP/4hbxRTXSgdHGAHZDqGQJyJozozzXOQgoKg1Dca/
NtKdzGRpYSdfIqLELxxajKWX8/7NZe3y4Q7CVkQaQAOAyDPVR1c7LcqXqZ1WRt8Y
dcyoafrLnNOjiW0e37FTzxmPnNq8yt9xd9RlJchLtpfPjbsNEFDMuLewxyQedeEG
UTu1qy6CLpxIWoOECBX3XDB4v8u+bcMNNoVRjaeCZLjTF088oqSR0Wh1+1wRmh/a
/aCPQhVPdbDld+pnDaTOAFypbYGAOVYGddP8YSd7S4G8gdvzyM6tSZ7J2XLJHD0t
fkTevlPHPggqvHmHAM4FS+cINaGsohOdzUwISJwGKWqbPOQPEskO4FOlnozA9og9
TLryOPSeQnY8ozT0gPBg9Y+M4QLg7OBSj/rEtIDtFhAmYtoZYAWC8vhTVaZ9v5kf
oOl7p0aRqr752Kzo91/qhKIMEk0zgV3ybB719U4I82QFhQRpdF+o+/i98ng1xktv
QUs+HTOK/V9Rz54kn2NI1rM7nPRmvItWOO2FVMXGKrbBEgMsaaZHSlMe7FWfzv/e
Xh7xCRSOcdnfibqhhLii6m8rMrbkBjHMHDaV+u1JdFdtkac0Oi7zBCkDek+JZQrp
YgPqSb1KzJNsLaojUacYUhnPT6/L3vY3ia++CwCJqbPK3SwmAWuSwulumzBQMwz5
c6b3wZQRcQf/MuFhiCYwOzc2tUXUuL8aJ4huoDrggD0Xb0WeqnDAFNTMVr4wOxP5
g3jwJiPYYk6vW4DsPtrfvQSE2SoaouVADGNPjbh/8/joyTIPSFEaxZMVEy7VdBkF
dWNKtuFQdH/OM3VAzId7u1OyNuucUvuca/9BrdYhQCZw3T1GapGTDdRDzIPt/Zpv
WOkHMRzjbg6Z05Bt9cYx6eMyP+dZD0MvDug7T/6xI7qQNl7AbJw6C/AP+DcTvee2
er5mE0PZiZ6LEZkUjBJDRoe/gGfLTdYvSA56eclm95JNSJUccb4oPwB8pZzjz/OX
qAS8UANDDXw5hMXoDH61v03rAKLeRqmg5OHElk1WOGiEHhmbAsokakKsAq9ZQwjk
cHvmCtdi5GQtABOPjmJ24Zovk04TcY/RdtqF6y67h6PSRYhv8rvgV77bsJ/ZEdDk
G8/mVVWhgTQqJdMa1jPR43nAJwHh6Vjo+z5PNxLSzCsHb55kC9Q77YrLo057+2OE
8czIeVZXsVhKIep4orpdKns48Nym+LTBDpWwMmuw7ccc5cL4n58ipqS/QcV7WFty
6Xr0KqTWhx6v4k5Hd/irzfkKQFTJMvRj4QFDxWtmmCldho/mfQyKDbIm60pMZRe1
NOut5ShoFPIMsaQ5ISGy1TL766JYtPECuOYiJUSoNcCDI0GfdXXYOOPJvqiK6mYl
H15db2AQL1gyPj0FVX95DPr6LyxTYV2TYX1GeyPTN3Nta0MDcPTAVHEIAwdorF8p
gX52Woac3KlG7XvOpff+ja3fytL55fofAjCT2u/Q0TE8DL/OhWIcGJBQ7QZ4pEnI
lPq7sv0Ki+27tCbrmrC8N5kbLQRiA+cvguVD4+6GURbhgF1sYPEJ2Go0qmd8yM3g
urjvncexIB6FLvVzYk6eCUzX6l2AwYvbmKKuW4e/6yr/1oT+Rwolhz5B6Dmb4Alx
CqWNalypOw63ECApIq5Ff59fuLS5RnXwBbv6kmpWXJ8Nqv66+Ofm/+eMDom+ejFS
dd+ZjvX4En8smuTkam+DmovROvQZ2xLl6e4xnbW2Oqgnq7AbMNTb9NSumcfjreoH
ckezagv69bIZewatuYL5FdwbOn9hlko4tYlVFL/T99cmP6wGXN4cDpCdAC64dWQv
SPr00MF2snAUFB6XYWoaD4G2YF+JlPriGzdOmLdyK2V5Yjdmi51g++UGZ2pcvGdN
7EjIWg58jzWquksyhbf/I+G+BGcg/6vK526UBoQm07s6BSFB6GNlPDgsc8XNBZos
qRduSVXv1rRbP6h59Za9d9fHKAULgPVGkEVLxrNykfbPCU0e2JjYdf+OJzoJ35Qp
zxbultlQbxfA/yg6QB3VgqhuIcjtxPzur7SiltZIlu7mFWwXXu6Ew7naiQgVPSQe
ja1ptCytNwEyze3s/nY/rqchE5qmQfavsYnmZ87IKOn2VU+U1DBvA6AlLuk2Wga8
BtUcN7f5/IdDoFwK++XOosGDqhkiBAvTHDZ+WxLshmfYTAbo/7kv+xY0yffSWAXv
1AwNa0rW5ujCxe/PrMYuHi9+D6IJhrmB8E3QQZQRYpwMHk+9i9/iSUkJQG+fHqGX
zyDUUycpZnfbfo0Epig2Q6fvKnWTl3aifXUR8cviXyoOGLBlbPu0lhdE71Itg585
/GQe1N1zK3VXvaJvsZ5r/LXy3E8j+NWEiML5XecAIawrJaQgKWsW2iR/zZtfspi4
HW/1VKe6aYfQbyfDllIhxolzPiwXJ7jJB3SpbY0vjXEOUuowD5C7svPN9NzON3dL
8VzOPTOc4ZR986eUlsdPbXscOlowIOeTqX+8m86mWlUkvLF7QKrhaurJ+gCfqOXI
91My/2eGCE5nbHkUr7wxkKw/BfWGkcXAz8XWXA0JM+TR0qtigpmwWlwZ0yH/UQoD
k4UKF0xmEHOEW/xh8uu4CjZw1DQQ8vKRw/R3AT2HZkGRJBSo6pqtEXdicVqnGjGm
CFZno3g+dA6SmWtda8B9jeYFDEd2iFnbp1In30pyyBPVyAy8xjrS29fLBQGkxhPI
Cd9iEE6/OjxxZz9Z6+WdUmHVSm0bC2q7PUT2vZ1O9DYSmqMvr9qQxH4FAndmVhnL
UPTgDG2yLaon3t938cSosr2Mpbya2Vj07gQH+Id5QKqJ4sQKKE2DaLcChgYGrspS
sFA+wjLhlXX1NhoUTn8e8CBO865xbxldMba3PVy4ZFB8z2Omn7LKOxbdsyqbzaYl
7UUf4wMkikWC/sZ6ZoxXLxZCF+4JjBKakpTdWa0WpwUFv7QDqwo0FLzLqKbLxGAf
5eqSM7i882KKpGX8Z/h4gCP68ybASA+oM7tBtBvscu1xE1ERcCCOk7wY4O6jrssy
ACFO9EksNPCkWJ/yTknBAe2LXaKzUB6eL5qlsOsWGAo1NKXUTbTAfHQK5LA02b4Z
tLV5eR9bfd2JaZj/e3JQ0EfIW6mUxDew3fbMn9urNnMeJUXPyJ/BghoLAYspMFXF
4yzXGjsgyrhCwpKxExWEi7DVtG29vfDV5sYMzVq5Te7eXfMzhKbGHPU0ExqCmaLV
GbA6UsDYRCg12SmogX1QS/XphhcjuIDs+XmOOwon2RJoFCcmgZYaUHm1ow8VtIqF
fn0HZ5T9O6nrTxJpOefGzxaMgpf3vcJEW8O0mvLZeq9afw2VTI5vHcrmiq+JMYS0
xW0B7MsDxjqjlKQ/fGik0Hrc3NeHp6p2Xbhqx31Bkf3zwi4Mn2Wx48ZuHEF7QnMf
gecdomd+Hac2BvIg6P7RqV82BrfjIwGxoRgTZQgNG9HB55oiF1rgfkoVtxZPGF7n
srlKRo/dxQpMv8WISAW/34kL6SiwOUf9O254I/D7Xy52INLKYMMj5cbbVK8Y3/p3
N92pmPDYEJwaIuC9rZSdGA/X/hdQfSxc26XUefx8T2XzDF1JKJGL40xsSyGwbtdH
uRPWZZgPS2RuTe9O0mlr6m6iDQMJWkGQyyK+Fcy558UawW2j6o9uLAYYyPvQJPzt
pfTIUJ7vdWSxPHYcvA9fOXSXWxT4GF1SXijOSGzigUwqTJcH/J1FyFzemObuK1sT
Gzo5sUlOGx6jrQ5yditfZNfrAEe9dn6gBg/PMBmwdkOOLy5Mc8ur/0lsodSckFGb
HGTOPQaTO9z2evKfa32J8D1zsdACtkSL5sKpNuytxT4Q/0mfAwzcWwFsp71hTEDQ
8qf0jEZIMQH+ggtg3+umCRL7qlUhCUK26c8k7PKu4NH5W2wz1CylQNR/NI7n0Qg1
gHjNPWLakI5TcYMt2VlUoKmGYV8tHx7jMe9+xZ9qi157cmH6kX1VKH54Fy/N1gCS
0z4KJDwULwYP3bOf5sRrtg==
`protect END_PROTECTED
