`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LkcMCVIHLLg4lxhEsjlzOWXlIbHVIml9gTqsEIyisD5CcKem6yBA/mMxO1i/OUdz
9JLPZUcVBre3iSRDInHFAVbRZt2cPB6DK8/cGtc04f0ahPhorDTmKU+pqjXIF4uO
ZrkLFH1XXFImfkPia1GY+448txLkqIyXlrC1MllqKV09EClwt6JqM02O2/ZGKDR5
/z4HMsdtpP9b2R4gXB2X0BrlorEf9QeKsgV1iltJnzN8e1UqxAXwZI9XEr1RRuF3
K4Qx02VHrgWTofFJhfL4iQYR3d4EYl05+JadB1w3+HriN7RGKo0JoZeiKjAyVdpA
SwhsXHfNLU2G1rREsg0rMrj23/y3y18are6sjN+C+QpMJHdJh6Y8l48B3YCc45ch
`protect END_PROTECTED
