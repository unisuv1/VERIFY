`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
JOgeacq9e2dE37dYUn2+XZ2k6+EXIPnuJqzSZUx8fc/v+X66k4x/uUtFKro0AnB5
xlWyIkesEazMsFsgqFfIYwaEfGvpt7GaOQsNP0HaIRNc53RtFX7Lnwn07TmQrChq
4jg05wlL2y6eXQsusHYYBckLipb9wG3HjB2Unv2j9W1hiAXyNZ0T/PyoKK0QhSbb
wPrVt2lIYOrkYI+61bHY6Ebax+0xeb5aidPmtljzGPfq6ig1+0XTE0jLEVlTj4WZ
k2sP+4egrhPF6mMIj94dMMs8juDAd+6LknpOWPvCPOwLrzK/NScjS4pudP9Yvpnl
u/hdMpZIGutN5cpS53rGZUZM/FZNOmwLC7N1mJlZROMMvrzeLNrNGaODCpJYVm43
QmnLl43IuFhx7SDf3bdaSj/MxzJ/Afty3liofeE9WU4Kh8zYj0SxZM5rPH+J8/yz
qp2SMG0JxAqKt4/vS0ToYfBj95dMqFmWRC/Gabyn3GyCAaMpwKOpt+IZjmg3LqrG
CoOk2T6B1lsanTivK4i1wS8pKVKs9UHISj1WsZ7R2QBmSkUmhuJcZYfqyGZm8dZV
da/ox+PmoBPlH99nqpMjkZ7BjpzKFsRnLAVkS5PyQD467tLbqvUongeOnHyG3QUV
N8dlMDa5nH3Jp5wbPdEmYDRgaRIGImpogHBeBiZJHnyy1kOznjoO3+G/v+mOkh6c
HQ8JRL7t8PUVTCfkd/poOosrEebkz8iCXkvDDFkC7J0SET+MJhHWz4OsPVlhcYNC
WcsvPho5Dtv+k6n6imfXfSOVCuX0UIhO9YraQ5hUJe+G9Raed8+uUcsYAQadJXa8
z7bgig9zubKwDh+wgn+9jo6oXCcvTBL1+o9HuDdxjRHe43ku8xVneWl6W/3dOLyh
LkebhE3WE/uU4kDE5IpSMNU7rurO4tv36NW8ZcDKVdWoCuK8loj5w1lXAnv0iLYd
pBVBCsvJeteCh0VYpnr29MERs3bZvwDrEZOJ880aWBg2B9lievDSDObqH84DsW9C
nuETX5yXa4GlG+/4hSGbMHiKx5/gl9C3fcuOCZCigxloa5nL0fyJtRDrU1yZbKn5
KB2A9cyFOofn8+Cyn5iVztQkSL+2RUP4dh3ZEVx+KnNPHLD7SKsId9H0uWrwIxPD
bGWR1JvXBEiQTLn5V1obHkA6Th/Qen/UwSPaGKoZ/ZEx57OoIEvliNxgGSfHopbq
aXwPf4WbPIFyvsamboX1oNDwN7m7ZhnSCqZMyW9yB7X4qQxdSU4amGVt7CP4xRpI
MphStzcsjLca45AyJAEveP5uUKHHlVjQxRSHDcG0AThI2K2P1BWgY2yMNRTCDRAg
BoyqbsdmgossSCvnB98G+HVXzNl96k3fVDWQJeQOjW4wxRXKPY3zZGQ5OjRkQz47
LfAvwIUO0AJyOVwhYyJGVBqmFDLD2XDvcgG57AHEk9qY/UFapGkqEZGgsKFmn8uK
NgFAdf3tH7SzGu/VeRqW/WK3VJqSW1Yg+dJaSIUkoENkjlvtkRrmsv6RaMPtjIzr
iq/6LbMtXB3tSmdP5BoGCdk4MUUZ/NEHTFUjX7SomaZuNhGlT2XlIkfOlkzpKZrA
+F/tNsvaHuqOx/BDv6zekwo4hHAuP7L5XYZ/EzZzl2fK3RLGd1KWcLI5vC39q/Ix
t/jFRKaLnDvpNZZN+VWG8UKAIjW83nzXAsUhAeLB8nzFKV3LKHzisphnd2bI49WM
uBomHAP+Wynelpd2J8FrUalbp9BpmWPTbJ/pa2DWF+/rpk7mvSpEmORlSz6zOxNg
BSPOb68/HkWsgtJ72O1+YXEPPQ+QP5k+m6G/buXAzfxbijUxEkc78biHOKSFAVWm
gVyFvFeB4tdCe1xi1v8tUIPG2AKpkOF6GnRzxgj2O6zxUaTLoQwIRDqICZ6Y2GLZ
4q7MnE5ft4K/sUmyOuTIXVNpkdWDdj1ujgfp7oJa285JAQSxLRCafI696FRbaD+9
xJZjZ92ylZw0YqRQZepyikyM9wh4biuY4Qq20fMFmxRu70PQfQMuEoITS9HjHGla
HojcxUu/eTMOrRCGr9nXBX2zgUVBVRE0MKJSjxaD5zqnrZ7vLHSFBelBthXz1T34
77Mz7Y4tn5mBndEABaa4JCNl1nNQr6beFT2rk6WanA7gXQ12bEOSSCO8xvLaGqCs
KzcYxMk8LFNCrRUtSE9lwANjwO5jpi44UnWGV9F5OPExviJvLXF5vLOPVy+dviOI
kcKgW6Sc+VAAyFjUBVa1ODYoM0Td9KxrIaVMMQGDrtsIqtu6Bh6ymcVPSYTq4ZkV
JDLmJU49jwVVkhZos6UedJBVmGfoFRXQfQ/UJmtTABkUxcMjJSPdMI/wiIVopaM5
6nKaN7Z+CcJVyJraWOYKKEH6KmoJf2T+k3jjEhrk4URoc6W8dsP1LCN7OyU865YX
PQFOxvnm5pANPB7S//F/KqiOwcMVCgSwnHm8+QPP239vqjCEhCGCcqQNIT71LTtN
SOF46kYb/1An9657YTCe1Q1ejF40lISajWAhGfmjh+fbicWzsHr/9itkE0gycrbm
05g3kxbj8IlmD+7wOD7dVF6xlqfOIqwZzsr+Zda0CQM3oZkmTLsuX70rG7iZaBjj
LOlAxLN+8bKLl5u0OF2jyYudYlpmhFc1p33ztr0g6B0fPVqsjfAkLlHWHL0lQfFV
eqncvokGKIKSL5taz0e0UYo1hiemYJz42aptgxWhOZ00RRh7djVb5MPw0VI01A3t
eCjM1ljvMesLYvp2lB6V1BFQnvA77T4aoV3slTYrzYT3eZijuStpZ+0QE6InRO4R
koh+pkf05MEzLMPd8pNqMrWXYrjLUsJpcu0zrJJCSErvuP0zaBQ4ynEeuLXYamA5
fUC1xLTq1r1VU4jvEg4piny/n54tsiy6HmH9NRTisnOGUJGG+8XJntzw+dqCmcfK
Jm2qe9Og66Kvnjc1LQvegoaV++77jPpn7CGNhADtmjSfiHf0N0DMMaw/kHujR0gk
Au1biu0StwrPTlHO9R4Fpx2ArdTIu1piDpebUsBXMliP2Pv8q4cuu7Q3c82+wN9O
URKn7z6D1TaLcwULYEVCIOwLq6/ezycE88ibB2ncl4NCP8czkGfKwDsRpUzozVaL
pE2Z2RUL7h9krU1eW6uDGNFGt5bIHMbefJwAyx7gg6jUEW9xMyeGy44sGoJhtWSt
5JenbyHcLW7DsCErd8sm3Rqbs75I5y/54Mn5RNfvJfN5gSBEEUwGPCijiJpClr8z
Ua/xRrNnGs1QASN4dgzMkdFYzkcG0xIrtghr1BIxzVLrZBpL//TM1xm+YHrUk5+4
2SR86YCCcOMsiz2gAjLsLJU5nYfB5YhtltMhbPIKvePmzJ6YUjTqWQBNSV5cm1no
bRru/MHJN7lkzzS2YyusPtAfcGxvBA9qY6ssWF0Ir7Qg6mVG1GbRi5juWKTQI38M
zWF0Zche91j6LaKlGHxBHUtKD0MLKMTh2Fv0QzyBFyIeUjfmj/1tlKLBK0X6YPJf
wzYKMxS7wDo+MWSSOywTKtju1OfKXObuylSoDMKVb+ThQmEXru+1o74UAaYKOOLr
ICCc47vGP9kz7Bz+IoWVytu/taluHGxKLPJU1z0rCDHrQqDvRM7+uFkMTN1JAIFi
bxnvF7q6oyUvXSbISxa5FPjK0Q1GJA7eUlOquYgfaR8qljAUh5WUikONulu6m/Uo
TCoTklB1pjFFOnWXgQiUkQWKAFbRtLERgzrp9VRlrVCzKLx//wQr9U957gOX8+ME
W3Wk8D87Erv7YPToVJJxUs8I6Wxotiedzl8/a6QIrx8M8HCko5zDj7pnAih8emCH
B69CIPV1aHYB44zSf288rhueWjTUdkg6G5BAuR02CFtR8lm5xE16q92ZUadzKLkd
gAye+sh2B8owk0rUJDt5STwjw2lnMTh3E9f/Z29DEWVHGH/k393e/sKXPxhwhges
6eVtVCs/WTI3oc8YaFoRyPvU2Qr81SVAgcDOYNkfSYLujVGweKfDqcOkdF2m7jM2
JpKKieSsdqAopdoLcnuUPN1I6BD3Z42s63SsRMeVJB1mggjzyINhnCdFdNnZwRvr
Bfa1kJgAZAb6qvcohRdYHwtfaiG3mZRo/MqXrGnZqyARVKhiyWM+LfT9019Me4c0
rkkPsyPwWSehyvUE3+kOz3+OOBGzbeB/J6/sviz0702k/c/iziX/JWXEkfjU6lIN
HH1hO2f7JifccwKq4oYvd4WqzPzoLPC3vblKjtvNgq+k6ySt2KXHybclOfR4rbj9
N16uMgHsyuLhoSQYG3OJFscMLyCUvnYNfLSiA/PDCjSTNoaHYrZQvc41XTVaXpk2
8cxjkW81KChqNyOmfy4VSCDy2SW1n6VnRCstoqNkiRb4a4QMRBWpCxnP1Bvup0/b
cnFupC2P3eqUXANnWAPQku5rYyk6TiZCq/9WFjTT8+fpMVDJgkthjFrNGon0MhVY
3peRCDrQ1Z+DTV4wh60tndxEve2lN30AY5sJrSPYBYjyPk//iP/bEe0v9imWZLYW
lanJB411iSEAtWuC0zk40gd9FiiBtkJmlPRDtiqre/usbKKBOFWV1d5S3BH0HdsL
Jm32roHlc4HRhfW3PRh+WrpAOTRxLE4iWMxZ60RZko3JOZ2U51IX/qlBOirjcr1F
MxG+lef6LR3M4wg4QmQphmPju+QnPD14mPzYxPr6R80svOO56xMqa8vhdm++4asY
fzoT0JuegyfdOtetnhXJYZrzGyabnnSdeqObqA/8kzPy8PP/50jKfZ4pDszX1piu
2bmXqe3tKMK6b0aorhEZbgHbFqch8pHLgzN1tWGFh++0kZOF+/ov79vototYXnD8
XiDwwyXOizDGUhaaHwULH2jCSEwHN9uwGab5IX1hRyp2JNL+wShNsSJhXuMSpIew
acsZIOuENP4JWX/iulbnXg==
`protect END_PROTECTED
