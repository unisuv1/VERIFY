`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Z9HybGv9OQSx9aJO4XTtYAjlluGlogwJ64N2GH13MaKdgGtyRLwGNwU4DKzC9TLr
/9BW9H5ipwFKxDNlKeZjvzsWTqj62nW6+1QmcfBOticgU6lJyaeU88VK08wsm5+H
kpANXHH271nn4S7BTzckVIfXFIzVriUth6xpyPmCSe76ZWOALxwJfYp9GAf1jUNY
l6O0uUDv6DHtFcj1pMWOVcjS4JtZFqTw5rEntU8ud3JuZvYOmRmchYcsOVhDHSi3
nYbac26f/oBqmzsQ2mriWthAm+9DP7OchKsu55QdXVURYlfUaO/CaQ5t6QTpYZn6
kv81ztA12gDsJU0dLHXDsXx+stYa7q+pyCTMvms8Wm3WTWETZEYHqxyFn3vgQp5E
gaF1rYhsWC8IBoghf65FaYBwKhEm4TJJWSACBFs/8MNpDg6bhzqrVDHrxZ36Yzi2
UnhCPbrq1fAl9ZYJrpnq3iI3+zItJp1HxyisKbnao/B8PcJ6rtBHTI8E4A7xcIRK
Nm7IS90rJab8PP30VRjqnIBJNYcpVUufuol/NqfHV+bVGjN6UzKbZCbKM+V0hosi
YEyUf2QY4M1JaAJ0ykd3Ao5qQZoTjeMpHmk8wmq3GqIsx8I2p1AM3Zz0saREI+lp
lDczpf4Y99QCrNn+U4GcWM6y+FO8YKKGFQswplHeV+qZpsEaC/9TbAExiuGw+iA3
R0dbfIrnynkNHC0JtY3NejJD1Z4deyMxnwZwgpKMvglFfiED/EgDGy8ttsANJSqB
J4lMXClt4bU8WL0IAmqYn580d28qoVhqdqMUk2OtYRKH1QNnDmZqcoNcSpJTYzzw
zlZ7zEd0XGoCUm8aJRQFN5loLRQ8eIrLH8/EVOTb40k=
`protect END_PROTECTED
