`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1Ixcbi+DkfVLaBIfHTlkQ9Rx9KzL7JSfrTlYy6gYpg22PWeW7zaLnCqZ2to46cJw
T5pzocLQipUVZkZfHGdzqL6YEEhrRiVrk8m52UtxpNArwbv4us6Wau8OrYN9wz4Q
S5p6jA/LhSXbdVHgyNizxJF/XLy7G5xlRapTYkkX7JYv+gQWET4D1JObvLagmPQK
ygoqX/JKzjKzvabdM79N1GSxYTHwFiCYGezz0VlcV3XkiLX5CHhpZBJCNN/JqNMc
bp9/+6QdY8O3h71FIYSu7tocznrbOGGvuy5YhTvGs69lkm0hDbKegZkakRPTGf8i
zbQ++tjtr/Hx5eROmHuYyrLiWMSJ8g+WKbo49QbPZmLk7OQgrTcXOhQx7VQgP3B9
`protect END_PROTECTED
