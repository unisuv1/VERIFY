`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wVWS9Do2R+IxWMA4TnKT5YKDF/QAIZF1MSH7uwm65FyMfMz5/vijiY/b88RiDPWq
sxL3DAfjo53mVmE+ur4Q7WpV4mArkihp/B8LljFkrUr8PVaI0ybd5UsQBBaDk9Cg
m9JerxqElBeoIaXioSvXIw0/nn6/qJcrqVo3ov/BwnwZub9hjZ84w9+lF7VW+o8E
hbCiJgj5p7vVwczIulAOls1bfz0wN6W13z3HrmsmmXpO4AyScA2kUyPuVS5/3Bsj
q3OUFgfd1v9ZSo5dY0dREGl/HTPWdxgRBlf+WUFcOV5aAEZSLaIUkdK6TiFotpAo
Ij9ADzjZQ8h0fSqlzPX/6pCsyFlDuWg2IBh8KnDS0dX6OS6cWJH4we/wR4rPmT6W
9d0nLY0S0b9oCA740dagkBQrMyYcFN3lEwGcxYAGtD2LhoPs5jG/9AyvU7eqwMKc
51SwiEMAepbttBdi/8tlFnbqMu17W8fS9nCmQTByCqJyAC8NyWZLzz1gio8iZ9E4
ilG5gFBnJ+XP/i+nCjA8fAWMhrOI6p5nFc2uub5aq98Rj8JbSr5Jyh1OcJJXNZDE
32I32v4Etzp6QN8WbwQRXaT4yNJdgS7Vjd9Wh9hjMipOW85K+acCgbOFDUNzPyom
Io6OxYEBtjkxToRkWlKkELo8hrJy5qth4In/wiTClEp3rcMZHysmUv+DwOnA5391
3KEJRBqenQgpE4v2fRV+lZWr/nqiKDhUFTJ2jZC4dhetlJ6zF443QIPv13wLDNp2
Mglrubc+FXW8bobt0AX2aRj+lE+UIvU4l8EO8SpfMPyKqcisvbxtrjTpSs9rjT+m
C3O97bfnj82bEmUQLQVquhUz+rNP4Hb+QE/6pAnWUAEIkdYYS9ZQubIK/bOC8KDQ
qsYrcvqUyaupKbeWrrOL5bFL6LTwNOZyGP04Y3cKivwwKz98r3wED7HE6XG35bcD
bT80UL0Hgsk0cKoBsLZgN7skqcjYDG5lJbzu6ko42z7mklGlfbl3jDv3N3XdIlM5
aIM3z5dgNimL6vhb1ILcO1MgOUEONuAoC7pE/p/QBrIG5LIydUzb1AxA+WoYKBgY
+cBdlvzfyEHoZ61InTO9luZdjqpLKIGlqEiIVyKD041cG+CW8qyu5Y435tXBbb1F
buCFqByYY01+GxkB6Oj5io+Z/4SYlCC3RVakMfV+ORFCPthbsB0x+GYJ5K1BslZK
S//wcawZOhJYRdARrjP9nq/xuEr/I5UAvH+5fYn3hkgDRudSlvBejq4u96to8oO4
fIrmkXlt3QkMeTUZ9pOseMecr01W7uKcUSviaWL7F7c+I5pBaaHiCimSScZABgSD
JbNDNrPuMaMMkzvEKg0Rm9nD5YwUfVY32ODMj7RNpRD//5K9egNgYH901x+HLlmn
MsJcVGkbb2/pZlaRoeDYmkMWNBygAhq0C0N69Uc0XGmCpqVw/x7fSAeM6KoVkelA
Efld58DddmJjjfg/Q6YoSPsGk+1DFNFZo8yv98hb89qyDeg9q+iMvepfo9lTtkrH
hMq7CBGoQ4Bpm9IX9N8TBlqyrbMzo9P0vW8g5b95GOdmSwC+xIYWwVASTHZaa4kI
OZoCaRUcxOfJPC2UkzXkjSKEnMJhVNuNBgYMv1gm/USbdP3i4B4939dokSbggJ3L
5LAoTFrRvsc3pm4H6ydYr5VHxgVcpWFhkl80wuozDJDtXua2lhqOJYjjBAUOwFuY
Q8MOA/zMDUOdLX1+cOcFqxVQWQP/OT387r98jleW7eb/Af97hZn5xWu1a7ISiZb9
2oEflTpxdUHyl57fkE3u4547Pj5XxQPueYMm3b7eXCPO2DRRLt/6rMqKrR2xpuZL
FTFrkvDKGV+LNCThKYPT1obXOJNw7XlLmAxpRzxq1A75UYFq3aZLAXEPoJkEjJgr
8INvGlxh+LtjZbVH4VpuAY6upe7UcJsiK/pKcofKzq2DxpFX50U6mUemBtpQBZtV
SGMel1WmDLkeb8lN7XdERbavf1MWcACJl8doFD7YDhNE4wm8w19h1UkMOFazQb4O
y/2TviDC8jASg7Fo04ilgOPsSm6GbGkfZkygylkT9DaiZt80XRSfNefow3/MPvuV
4M6Hyu3iHF90s/8DmxFsqyA/e0+kykk40UyZyQQpvkrJjvO3GgGM48WtM9uGupbZ
oRUoz6RPuiD9NOzJJns1OeR/QcvS2ve3ejek7HUmwCcf/FGeNN1f7qkyTqlzfDoj
W2P3mcmmG63gQGKcL/mEkqM7bY2WEHY+Gac/lKXmHiCPffcHo6J6Wh+zwbKif7Uz
SYRGbMTGdzum/NA9W5Dat3p0vhxgp/l8ffqyqIS0gJUBh/NZx4RlVdBUKTOgJXe8
+Yv1gCy1/ROr+Rzy57IEVnXCEaDT9ESjevoGCwDtjITFkKCtRvBtkeEZqK4rGpmz
WOcALDWqCt5vRtTb9/e5GIqTXPFKDi1QGRzf5V74UM3DEyJUxZ75H1t374v0VHku
jTcpZsJaA5tfsqiK01dWXQDePaLhr0EDTpu8KRZ3P6M3WODFhm4f9VJeVXa7XIc4
3jeeIfhdkSqifORz6WnY3DG6imcMjnMmrGNk192YbWbRJSfcaJNjuguKNZ6VROlb
v16zmO9sMIA23dRifyQwr1hxTS533j6vd0JVfRS6MDbCNy2m5tmAYaNydZAouFg0
Yh6ULKrwO3ggOafVbpnAJUo4OXyzNwo4o3fnHmJBzYGuLTqhrn/JA4vUSPtNlxlz
EQdF4mGR0G/LEgJk2cNzRpC2c9dBtsFJOIIDkQW3W5dlzvMERnEi6CZNX7gUL5PL
KD/3gFos+kuiq8jE56kwAFx7E10mrCsdcIvGT0uKpn49Ysk11lkKxi0GGsBE288+
diSe4dC9rJib9hxlRNW2ftfCkCcli+H3gcMemukZGe+LrUtob+Xzd7utHFx2vOe2
t5EOy09qXgMpU1uWQv6n91hYhV0Gyfg3/yO+xfncfEunBHEiJWxnV9aAj2bFxiT8
PfP8KQXwGS/jGJARTJ4EvAl8hF/D2sIbFevCPNfHoM6eOK/eKCLLnjlYp7YP5ltK
BftLl/E3TM6A1WNpv06x3e4308XNFGDK4ZPS+OyuiLV5DXbAQdCmc2ieVc+Rsg6z
Kz4YlmMY7dfaoVqZUTO0qMc0iKp/lbqdTB1HrsQ/rBpzkzVBnxWybrtAXA4guxy4
MsUs9EHlfrGmJL0WDHFZlG4/N0nmiHpwjhwsUi1tX+Ajn6kKQ6uv+l8KmGzvsEEy
eSoT8RZdBzwiKb3rp6KKc1whQRD/ZeofMq1uLo3JRv1FWvzNfrnjwDLIg5U4ngTk
NmcATFaaqH1zKRLsdW406/vrtXWbNvYl2dFpSiAtH1OzOsteREiLKntepDKBfvs5
AqfkLnPkwReeXLTuQ52SkYxj6S4WPN0IwITU7aw5mdyStEsUycSRBDOXxQbIyXKR
9y1ezAf1MMD/CufMLxkRyy6J/R4O6FOAOkaM4N4Us+Yyn7TAWPCCfI1nfwx0w+B0
/EeYrWIP1DPNjfJStLf/RvQb2EaTKdggEEzF2r/PJYPaHXyCjaKE3tQZZE7+n3gC
c5fjYH2TBonasjLeuVbpZApIVaWnY8O3Oc+1yOUdCgTKPA3aU8Qj5l6QH0NSRxBj
tFah9ASlHMMLonZ183shoNY8PUXWNBngZ8n8RmDBmt2v6HHu6772wjzPtl+NlArz
CXimBwODewaSTEqKnn0XUkQ/2L+tw1bl/+MxtkfNvoObdjcWa2YolKzp69GMjCxk
/RokCGVYiapbUioM745z1NUMVIN/92cgtUALMDdrYvH5OT78/PSKZtjm5qjPqvno
toRPYXXI11uznMuO+DH2+SJsVSI4mOM7g/DsxKtCb/bJZgv4dBmAHsgB/imZjpzZ
efwA/WzHz82zJV9Pd9zxRQswRLuMxHWT0IICpUcSdx3r8i73kzuYoJgqYDkINjKs
GYpfwoIOL8b50oT4cx3Bom+8Nu+2i0pGjoUnVrJ8uUqmotVA9UstCXHJypd9WnWf
rHv0aa2bw5XMh0oUNBQBIDHJ9MprojA/DBgZVQvwhdbU6x3xwioIUID5xpig/yj6
2SpzQFytguFGoCOdIJPk4CPeIZMXQLZ1tQR7Z1MaMKrwyEUWIzVXq3ut963MGwHl
8RpJQihPmvH5H+I7exvZKP215dyN5YXOtWPkz1nSaCNMld1wdGOsdWEY8YqgCNP/
r+7mMeQf6fiHLRz4JrOQR0ou92PvvAUWxi79nipVSHAo9g2tUaR8beZ2y+2cfxbt
yDGT/1H4dFtDXAO8I+6xVNusYw7Cr9gxU48ASxJem+SZCQpLYXMwzqsYSnwdKkxg
ZorerYgsGZDnRMyzEIR48RwpL5ZRlQiKzHZd+W55ZF/XUa7Fzfs7speuk+HFgwqJ
k9t1eZdR8iBj0fEP9xggvL8hJZaMVXY6jYPK9KczpwO36uexpQP80ELXrmx1uryt
Ve7FkH6otnEXc04mgwimmFzQ7QbUTwC4cxcHe/dTMJy6GbJu2dhU85aBnzwStxog
CV4qLqinSiYsAiLrXuCyVbiw4XaLT48eUlX38+g7K1MC0+sIIV2PHNSCKNtfafiH
EQe2yGn2QHa4z8aGS1LeKi3zIap1qnGCrDbPJUCsNvQbLDoOVwI+2geELsgB37tF
HqWIu71nibXEphR20k2C9hK5bBVdf7bLyAAJcKL1B/QVC19inMBgzIiGeE07Tmka
PpnWU1tzLXmbFYi4ZCaWKiNjATnNl88XedAqSyZvP+EctB9k8Kon7ms4NZSbf+ff
BCr9w5BT9+1H9GhgW9ElSk8B3NvouwysGp0s/pZM66Qi+xkquyyiC5hDufOc2K/9
jF3JEp57sHjjgLu+m0zNhf4Yx4u9R85pA1uHDckgDqOZL3dn/xsgrlfqv7nGeNQa
RO5eJHD0YKsUJMfDe6X6kvyXlILHEpQzOMjuD6dH/7L2WbvEnh7+Q0s7wEkZSUli
dBlMO9fv3XOBTmUCHRvGbZPq+nkY4PjDntVUBjXJREfEg1pmgFHJlNHXEY/l3EQ5
EBrbIyL9mKAuo8/05EExo6q9bgGOCEED/4zZpcQQYI2e1LyzivibfJ7lXAFCtx2s
gKPbqC1ps1UbDSABBs9vOWzrrO/xA22nKKXgOE+LmYvFb3B7Andp7LZF1dia1qXk
SvBlAKLjCiXwK0SZnRBd6+1hcmZl1bpSBAlbv4vrfJ70xpFSuKFCPDs7/4V7CF6n
QAj27r36CA3XRa3Q/zL0GSCkba28haFW69WApPaymQcxZskM2oHvBidK2FmaXfLY
85ojo3kVI+Y4Oldqnygng5Ba201I0xDTRyx/qWB400jYraDgU+BGjCK+TwmVmQBy
jviP/527uk214kw28Isxms2mr8L3QAV1WObs8PZWcWZ90I3B+H77ey6zsrRbq4BM
ZtbeKuMDxsnklvpAkjqaFWhZuXV927Kb8LsQXMcWZIFR3JBQJ1WAML7saEWhBnDr
+LNuBPiExqaMx3smx+gIoaeGlRpK6QOX565ve2C9e1BWHgcsP2hCPQcoqo7Vy8fs
3uY1kIgnIMGQZR85ABp/Sq5wwiiJuhohPzTdyJQULFmRgyvYTlXd/ychmf9CmbIW
ROzsmAtd0rt6/6cMcGfLUcQRgiCU3SQjKfZECuNpQb33rGrmIwM2xjQo+KXbF/4p
Df7ox7vs66fiKiWQQhsura9cZl32fh1oUwV3JgVS3FGUIRFPFfuYJ2pHXXTcnH0R
a22C3sgrYRs2EyLGUDorCqZK69KS8M2lkoZo7zWs3BEhzx+8AmI3+UuCW2sPpX2f
XKD6z2q2DLQFUbfHCIDEONb8s7Al9/5T7lkyB0eBwxZgQ7C3cZJyLKBK/BoVku29
SzUCdzNuQSa5aIZw0jeeTs35jPHPrjLSJyBK2VXyzA5HhYrFt5AAXH7t3I1++Dpa
UdXhHgW+7eWWk2THGXHT650oFKvfGrEF6ec3GrTm+odY6m45iDxRHbMXa7DGlxv+
/oUagqGkkLlm4V1ppYb441KKGbIwNx/9VF0JJqK3Ty6UxkyeuOntg0UYa3RAD57d
Td5R9oheNKz1diqSEjEahGMT80yfVCgaQQjXtdWnxIsnkFCBc3E8ts2hzr56aB2O
FYqvYiKpFOHR+91MhsTUaxN7AYTvDwDt8OdSuO1M6KO4FitGCjd5zxP30GIRe9qI
IdVNZJ4poq5i36LgBxZqXJa4EYsnKqQwXRhzz4CM0RDlBxIP/dTnTIVRMdfo3NUS
Yd1ziYs6OR/lEWt60WCbqUQ10a/PV4VTCZjiJ95P+plwDN8X9+2JpLJxOt6q7Aup
xV2jCkyAl66PE9aXKkpMF2/0NSPUIzacRtYHNEdp3fTzUpmdIvQNu00uv8hS6215
W17Yl/376jdeK4qVI7/XevAT86X/y5QM7KIXBmKWoYIK29eMMACqOvAcIBsfNkzb
DJfFAeNzAxJteao2IsbtBoPudPlG8UYzzrzzoL79VdvEzHlUtula0jTGUjDasv4e
k+CHwpWrE87WBPycuMcTWJA1E4o/fjKyv/NjUd/oIVq6mLx5uNQb4lMG1tJarq0W
sjbLSrCi8SVTY7a+bLVnEPQGeiP/HMtVZL1H1njZoPxNS/Ay9tuJJxTg6kWP0yU2
ZJsKpGYS3cde3wx07lCOVzqeZ0xLoOjdJQ3eaytmFo8fBR+QNpVeXU3H6jSfeSgU
V+IoAl1lNnmQVO1J0bOJo6geSQ9XXtnDT+KseEvwkANNHsOc7VNNPaC4t6jNJujF
zIugcq5Xjfz5rNYpatjB6GSIzfnrNKH2Kxd/ku7Z73oqQ9Gl4QzaNV68ehP8+IM1
+PDYhtvYoQc37Qydk6axCDzQl9xR+W5+swmy86tTqwZXCLzZW7ASA2rtBDpnx6AU
EVL5wdIDThdDrdrlAPBWLvqsBCy7Qf02GR+VDwRTQb/M+tnDq67xDhdlxtxSw2IA
yuqoelEcn5SDDxy8lzGoz6eyvKbVaYqVSV85jAIrwMuAxqqFmfYeLoCZDALkrOK+
daVzAjU7skK6Im66ZUQu2k9XwmriLMbEetML6YuAUAw728bzCUUWD6YFY32Jvv5W
4CsPQ3GWMH3J1wt4kKKK6dtIKbXYwqVlTJ8ca5xSV/Ihc8SmCo4a+BZrZoaiSrUz
fzb9b7OgjbOxXkAEZ8dVmbSUYK3LGyNkT7uaDv/ife0OTXiYG28NBA/4G3PUCb3j
j6DWEw8rI4Rw0d9wzqsLH65rVywKQhu/z878y1877IykWgSM2I/j8t/SzQpBkztE
QW3PUblvZ1eQevqV7jSic0LinKwR06d56jghCS4ENqNKrBGLDK7V5ALlKn3+5ALR
dv4jtCJoGUX2iFH9OTj/KN/psc3ypKY4XeinkGCxr2Fo4t5WgtyMWPZg6YHhqnQs
I30ho8YK5GH2Te/3fOZUtYUFEDiP7EDtZLvmozOX8aGJ5AzatNVSKQ+td3Aequh0
NgfzyS3mdF1LQ74NIxuIZixDMQ5aGs2GDwJbpvNH1y6drglMetvOYXQuVbgQr3xr
8DG3OZ/Pe6m4K+t12mXgycQ480k3+wVuzECPjRSadbxnkwVDuShMrH/okFnrir3z
6dUlKXtchal3KgTqYnHESXVZul8X4AI94j4PpWLEQzg5BbbT6yxQ/tMrgz/K2PYQ
HZ+gwo1cvcJzWwVqylsuovVjsXDgqcyk9fD3l6vr97Ztf8oOvGbYht8E4EOreARc
h95LI2n0IVx/Apw9NjaOnQ/98K1I1c14MptwpIcT7b7E3szKnb6lhOVcq2XOpFKe
MMBpb1Tx5tEphc0B8dc0/j1QjDui6iV2n/AF+2NhTZ3L51vz0hi1qUoCbbIZrDjT
NGuZ427bFn7VPuZ6YAyb9l/64grTyeY4b0OILTKloj5HDvGDB+zSQmGo6xniNde5
M0MDc22ODN5KrSTfR+/kyp0MSmMCLflEesXoIEQ3ftywbdc+TRjtiiTT/2hcWBP8
t1KU8E96HFFE+csMBNgfxsCWXRddvdStXZy42ES8YAg7dnI/gNZBIHxdDHNTMZ40
wZYKyF/hrWDYwCMfnIxSHYY/BvuRpuMGxph33KlymeIINTv+wouH8HgkFMVu5GdK
Cb3wgBuqXCXJbwi90vPnzBI6vkJ+pnOWGtFwUsqlUnS9HMaW8JDhRlwz0rTlmHZC
hgKN7cN2gQ0irpV5/H1LPE4DmlOqA6DsU0seDgA1GajR3hdigHBiXoBIOkzFFs+f
O5dRlfRxd2BKXp+WhQF5BG3MlThCaEmkC73J4FTGX6MSM0CeYcNzT8XpR39nntvj
dV/Sz0nF7Dy+PhKmZogPXUVfqB3/ppsqehfEoUNoEj4EJYHqyi3vC5R3LE+bvnUR
R2BhqOaL6TZAXeGaYOD43DTGYQ+KWb6Ty7BojnmErQJ2wKwuW1TPFXtJUR5zD+fl
DAIpenu8zKNeD86eVEGUR2aBQKou3aSxSYPo0FLAw6TgW/uF7189qI+JpMCjcbFV
2i9uQyDR4MXr2Fe5mQIUXspSCL5ZmjmMGLrT/myx9ND4KKehZO0HiPCnZjqLFSi+
+AcQCgQfgqK7ry6ppB8nLzTVQ8XRsJEIt7fKv8Ta3tjFhWbIifd809cbxNpqbhZT
VnZi6ANp1poiUsh7sE23Cw5Fn9NEGchxoyrSTQLYsuxiJPyDBFfRXMxMO5g9ddLv
SA7tWhCRosz9bLs2f1jCLQN/Y+kLfb8bvH6GJCPLzsRGFOHMRoXt/7/DJaWpK+VK
FKxGHnkQZuduuY3RW/ajjeJabZ30kHAuZzkyegN5GKzDCyGyev4FUf1/085Krg3j
0wNlEJIgAtkVkgvRvFUhwF5x4SoPupRG82IpFgJnXQO4nZH2foCmLzEWMx3FUlDe
m4eoa0KU85Sa84Zvz6CtM9lB8EC8pLLklZWeUUHAAQm7ZMc5idz9yKSS9z6wxlbA
v7T9LnpJg12KS2M+KIJxQPw8G8RZh9YAG/7CvBOAezj3sADWTCGLDp+bj5a7GUIh
FGEjvft5iOQam/hWy594ybPG9NzEDNZD8r1fOft8+rqsFfFk6pOy/GXmdptRtsuL
tWldtBIRlMUmIEngXuYFiHOSSEKwrV03qtEkVNll8zzOwmTsQKGWFQTDlpY8A2i/
hxiFyqY+FYldiV1lzF8k+RC3xXZjOHdpXZhqGsDw8CTE94kxy3xV6Tycx0JTb53s
qmax0AnkPJSWGulxw85wMnsjc2b1RCS/f/f3POgGBIydm44mdUeIualoKGIwxx/l
ueoZWM4ZBKOxBXllE5kCe6tg3O7SpyoG3FakKYk988u2imxGdvlL3e3q3/JRjgjO
r9CXhZV/Bp0389uuMz8h65Md0kwcpmSDg025dj8PL6jjLjdTo/OH7bYBOej/wEMl
S5Fo3d2CG9D8KKLhgBQEIKLH36p6/8pJwrGWHoGVc8TFlzu338JxdgS73lHvTFol
ZINY875lQd15K1IeoN+KD6vrkvJgXjG9dc8/+RYh09E1+Db6B3KjOF6Oc40EjkIt
WnNSb4QAYNQHKDN647NWPMDQWTaMuvEcdoIeTCNrxYm7Mz/JvrkIMIi/fXBgPeFr
8MaVqzeW96QbA+TKLEKUcb3Qan2nm1p6l6WP6nmPjQQ7vQQNdk9NwNtExvmRpBZo
JiguoUAg1BBoDdZgV0YDhcD5Wr23CG0HrZp39Cr1hUMSJmiCwyg52v1EHAZhZxTw
hNz1E5zrPvDFpZjOYbRfXwusJ9xQg6mvXh9vqvOZURkK3Kk6Lyl+cJM0f74mI9bT
ZQJOju/lOLwlK3NUhbM9EcE2bffu8MdklhK8MSof82kvwOuj/o4VfAYNM5tOl5+N
TPJ2KRaeZ9RxNPy9R4Jx+68qz53aAdd6YWE8VOIhy932LrnGqzlsDyAo+49ga0OG
MfKXDSlFsrVnucfZWtqv8H2XXIT3Vsp7HO024UAmJ2eKmpuxcQsMymQP0BpbgF0O
5s4dQg71p249WoXS+m9uHIs0Hq93GtItJdCLn3/Pxf3IF/Q1m0EmF/UZqVzBnArQ
tvgypQxZ/rwvZ1v+P9msYPsK6WcK/LLv1+vD/J3YY5YIK8gh+/VhpS59O25t9XMn
QwKJzAyTJ1C4zk9V2Oldx2pJz4SSSnoevgtYyuTfipFRgrmC4VoOa5HjdASe+tXe
y///NiH+NnVQdQXHrukgwNz7RzVHoIW6ulmKi1FZc2/cVlXYneyROynS8iSJefhb
VOVMg12QWqrAudyZKy96mN4S6LyC492QOwRTik9uBttlk5ClCPZTGvhM4roNRAKA
QpnKRVb+VhYA6WUKJDm2NrGT5SrLknlle9pKX8K6OaGxNtBHc4pqPxIFGQR1adkD
PYcTRuSVMvtJCZTtOOz6lcKc1d2AiJuFgJjHw4/wTh8SO1keUyLpuMHvh6u3ipTf
CvRhsv/NP67lgh+aPs+Ih8ag587L0mz8h+0fnv9anNQlSR74L2Ac7zwlIdg5rVUp
yavgFD6cIH/6DyV2wNCKES+Y5yD8knzjO/Ab7LpaGBPMXJB4Lt+WMK8leWSN3DEZ
pRs0Q0SCzeLqNKEPU54+FW/lS8xHo+TanfFS3OihUGemFPFsbqh7owZ59XKWrdq2
5clg3CmfN68uixc529BpX4OO+6yiGgyoT99TAunIoTeiOxarFiyL7oIeAKOA9WoH
B2aJ/hUDWYdMCPGKE5e39oD32fMuK0ph/n2MKOBqpz8HASMRZ/wv7mdD/eh2tPvo
Xwfpgh+tsgIK5P6LqmGJNMQneelobEJWo5YOhppBmexpggpldl9MrTeLA6XNuYqv
6ieetb7AFaxCzGHGoIe33dNysPAAtRiKETbl+jJGaOMtvffsYtNCADM2hGgcgwYl
+7gcl3kQTI03MjK3sKUTRxcH6D69qr9sgXE6fm0V240Ng3ywJeyFqMJbDfve8gAf
+9/SPKXuil/MQGHKiaXSAwILAACRWoWtQJlJoQJhcNQX43+fYMvmR0HDflQMrUGt
aYFW3Vr/42iqXgT/qU6ZGk+Z6XJi+OE6Y8MmDP+mELzGIMIgxdOa95XZZ5/VWMpV
52FJJy0yA780n+jW7/Nbm116rg1oxoq7hllhTimZS9ceDlaFknsj4dfZa7mdo1MQ
yRw2a7WGUKsrSvlkHsdrsGkfkWLWzRsDX5bqd/Ygc/0H64NG6gXz40qvi2b+ErYz
88nS0c8YlKGULGQ1vfAGUSS90MMHja6DLRVTTxvlzCn2wEK8ggx+f2s5Q6or1RvB
JNvc2wlYiKHnTSmbk/ZY7F3wUt7YoKC66TFfim3Fp2pQzsLlm0UsYqOR73ufZj4X
sR9uJslf2G2gQBulaEBUbuwB43saCZdWE7dF+hqZEjvjfNU1JSzCenNIWsjvUbMr
G+JDhGgDx+V+5mxXa8Nrt329p+wcB0Ip2tF+jFE6kQ1yrvNlMkXQTzBDGP3CcnQt
1Odh92gGCoyD3uQLOHQCCOHFyaxp4jJ/OW77pBYdScsuwn0JBolG0zm+QsQGI6DN
mBi8/spo8dWZVVChMR1VIuPi4YmEsLi+rbEBnXh5RmJ2SgG37gYM+ruiQlA0LpQI
nLNAw5EQjQc1xzgFReMuLsQXiGe0HK3NSmmiRu65U1PpFOcSWbOZ+o6Ahb4vdePP
xNf+BR+28Y58FROC5ch3Y2HcDm6ARLETOMh/kHZpX6VKDZ4nDdTFOdsRbAPfDB36
kU6ouyx/Z2eGTXWD/H5+rR7iyCCBKN9TN5oPfYYeoZKTadXVZfV8AJ00szXbFD7t
niEo6eRVJC6WJT7dK6n6+DZzKYYx9Zkr3Br8fTrL14vmu2OUPfzWRmrLacmlPI3e
yXVgW87ZiXOc7gQkiW+5IikZCJP9VB7L3S5lOSKBZnZQArFgUGsblo0yo5MKIVPs
TrZquUMCTRKjpcAx/TSoEjTAcidZ/YMX3WVm74JY2xRkcHzGMm/BSHrYvJGqjT3Z
c9XG8+z+GQbNvijmOBXOojZ5yeNCRONaCyM9dyHid3DcByR3/MQMfndrePw5z7Q1
sSpIv8UAAAIKLloP6mWT7zU9j+/L7JjFpZEjAm4NSXNwGxcDoBJYgNpy5BeDJquY
qIz5hywlJytOE4eC7D4XxrfjQVX2S7hQBbmRkBFUGVwMe77aTkjz6tWKSOlMTvdZ
JZOjEcYJBQqgtkp3GdJYspDsZ/UuorQbz9+pAcCOa/UiRC8Du15ie8JHDVYrITWb
sZEkkmxtufyyeXVjkFhjwzV3WUPxSYg6tSIhEjQr9pNxQggOXUW/aEDBgbatA5uo
ETWtQ1uNBL+V+7yfJxGhQ+2mg5M3gAaFPi7FmArJ12/G6rGQulbXJZSp0Vy0O7e/
Bkq02fsMhYVutje6UOxwAX0ki2oOGRohQ3096pY5TfediAoXwlVAcGljxqBehhON
gcQojua1cG2veN1BJ67EvphZxfDvZDIq4BaETcUuIPNmGfkMZ9kJYaD/f8jlXohJ
lFmjo0Um7iIzHchU7I7FdA6dPGZjv3YZcZ93W7/ijDgoP0VKD+DanFxjRmCEQqqD
xF1DS/5vS5eDsUmNZ3xQg5feCsxCSeiIg2IWXnytzGlW/8hb7sZz9GyDly5dfouS
u/JZF0fXrcM29JDJLcdaQX/cFU9zoYz4UUJu/TPaqUE3nC4REcNrLYNopPM99l0C
lk/p8+oToFHiNawDlYE9PL3IeYsYAtpqL/KcSr74tg4aAJDymhSi6lSuy7RabfDJ
5hY7u9903ovWnpvD2iuNL+/DjsIW4CCOzP5eeKwt0pmlBhIkEFUo9Ib/HU+cl9AF
L8giy4hDRDWap/DoPJOU4cjHobcXcp6KAguxQNFLWW50rI9aOB6faAEREkWgswtD
FDoikTCs7ErqBzvoxjo2Wa4DcaqWJoLM51/fnva5zByGgjRhREfNuCRxKZLpRJD6
R5BOgPpwr0wydMPJPzg2n+WSrfGnoSho37z2ukWADcxzyFJxlvWNimauymgMoUe0
zpbqXElznBASMoqYa+OziH1KqJCc77MedsTm7/SUZKNLeYzP168NiYwsblscmU/N
fJc3TQZfYP5o0R/zXgfE7FcIjt9lWRv2fwZSoiynT2Rk0MyMrXKKJQt+JRKvwwqm
dPPKCOVeTFcLK/0s/lXyswxSJZ2JdEB0vaWsEHMj1LP6wHEdg82rt6DUXz71Q0W5
us6OaQ+KvIENqLL9aipbXwZ2J4aauWhntEkVsuMhZLsZtmXOZndi6Xxm6u5Oye56
HCnTGPNtkQWU7qVMKcA4rZdDC9INrgNn9O3H9JW3MVFeAQ7DZ3lKg3OyeXT/jhMh
hCEkJ87GdP3tV8ea32ykMZqdnygRk1rytEF1137bgXjzbHfhKAbyQftmJsJvlOgk
7HAgOMBYq+A/yK5BMiXw7EIllmuuA/wQcOx5uR5TmKvSC9JnV0oE91pCebgiDVtD
ddZyOa1VHgV75f6V0E/qgJFMwKbAn05R6TH6j7OrN8WVZjwWZvrfPkz/DSG92D3Z
ybFFnnyQ5TufhM7dVBh02oHk1SsbvSPuawPspE9i0s3NmbM3Y6h5Q7SsWEVy99Bf
ekXvURJdN2wIAfEkwgqDvgX34dSldwaBUcFkicM7+BP/h4DjtL2gmAfNjgKHAEkX
x/btplHdJDyxj2AgBoz9/7tsCMtf5hBj1Cvs81itbsW6xxvPpLzluq6KC/TAhcYR
wGP/kd6fgV92gT7TUGioD0zPkYZCt6GSuIWntPBRZyV2hG6I0i3gmkJRJzqZaxtn
YWWZR8EyXJ8Z9IdKX2IYNXzkcInzBjRMrfSYK0VGyXDQ+HOme6JWPODrrrLtLVqR
qtndkz/ggKkRlIcVOGKvLQ3nTjSSDRv3zaYqSpdPhPBTTnDokEQ6hLXY1ueKcvmO
RANwD4qLY9eTM1RRYjk+293eYtqgGT7oYpE11C5sa5P7O21IQEUJetUebRoo+yK8
ZY79x51iDG9jgsVv1MJv7gu1fH66w5VvzJqow38jYmTE5duqECfMZBZz3YEGfYbZ
1ECLIzWQu9uuXl2IRaRBVAmmyWC86NqbN2rpW+qZtnHTBAK5hZQ3VZyALBrqV8UU
M09dCOCDH5cdWDfqDt/pSTzY/1Oppy2wPr1l3gHbHqDZP0nf/sDZTQgq3fE/KQnZ
Iooq75PqRqwDa6go22N/oADNzNdPTfrgoBi6MQLajtw2tniFR8RZUWMZmSP2losL
K3ZehG257Rt00D3tZuX3NRcWTR3qg3PVI/qXldExQ1qilstHsUsbX5LhQ1VOEKHd
wcFVixCIGiGUhfkvaCaKNrzysxqjKxnhFqZHkqTaqcM1y/hXBbB1URsBWcg8Dq3q
9iCdTKjQFeKtUPJqkFSFOjED1k84rNjVfaSCaFdRuLmA7c4WRmpWNcL5Rj4O9Cbs
XnPN/839hYFi2tHuV35nMaQfpvHN6Qbp4MF2VkvjcTkGE1u7R6bK3qxInC3GFoNG
h++CJWb/xIIdkAv2YadmM3kiB7G9bfnSi+yVemC+me11XCuYBhSze7ibPUc27N9v
5d++xaVzgjUdoOMUHcrjiqyS2fb+jVRgQrQaHrTwTbog4JNeAGjiwH+l6wBBNJ5L
11QWSW1zI1ugo8PAINLFBOpAVPDhavrFo89dD3CjFoEK7+9KkB9uBU7yJIUNt+fg
fen5HC61qXN40JlRNX8sG87MzwV+K2oSVa0yxv7jjIA55Ua7qXTm5KbEufAHed0P
eEFHfBByXUIYNVJv1q3JtMmMNxKAe6LfrPz5Tsqaw9lHavB4hOYw2CHFq0Diyu9D
dzhBeNJg7ZNliTPMPEuwN/233q5aOn/aACQ9ZZOtdqOIk4PFHxzo55CLJtjSySD4
118+OaIp9js4h29VOQ60egBmrvkoBZAyyjFjMXszh6RqxBACuw3bdEZhNxfKCTND
pEn3P+G2shpoN/OcubKd60mJm8GWVzTPZ3KxiZ5E5pSSl19EB56V1yRwPcs7DPQa
7IRdEuqC1apctDb5Bzyu3lX2+4h53quzQDnXVFiKN2lMpiGJZuwlk1q5hwMKOTcq
TQQBpDabAcugG3j8mV5fs7rhbOuIL288MiprLOinEQtwh/26OqYWeAhfJlMEkWQz
MXYQRrMjXy/motCeWJaqY+EuWXVersc6PFwTr8I7/bg/Ckca1WuLujCTXxwxyC5l
WeGGiBb+T73YXUbcqZ6lrIsF7xklqedKd4Xo9CrWTwH95xOUVScyD4Mo8y4m2pOn
Y2aQ2NjAs5p6KY8xksZVMIH68hoHRE5VrYG+8W59aHKJRfVVtvfEdv9g5FNDcb/f
O3N9Bw7xuDdY20qBo8wnqeXHJOmSGMx9OhZY7I7xRIqHaENF8aJavg4HoSP+qeIs
l5NpXp2UltS26TKxN7YQjTY5EhJhLef6FIbPMyIaAvTjccKJxtUHwOcrPoWLchbg
CHGndKfsUQD1bcQiXZFS06+lJMWZNtEbrrhELgWni/g0zM/WGiDbEO9w6SLa8a0B
KfdqkB/AxKEDWjBeIuhR8hvufrK4bS/oJxkEWliTlCJWVEKL9pO0Z0E7bAVq6u6d
j24lLzzbBR1o2tdfJjxo0VzVMhcDjwcyqCvmA7Kf4WD1iW96w6OJdFhxfvAHtfgy
lu8pzLr2iAsfqj0keNlSfihABLL8OzuA83knGWdk42vvcp/IcqghTpy1EjbFdr9V
xQ1h8nHxM/VMPqPaxYAy6umDRXT+1j0bQhep4sQcxd5xn7KSf42+OniUw2Tzlfd6
E0UqzgZ6m+CaOH3X8WTv9a0NzHPER9u4gzUea7RbF5YQCuJ50hf61LBLm/Ln0rMo
TGty0XE/f2bGPp8s5dwfSXyGgZDz/52R3TFXkH7N9nO2B8I5HM5FIdn7y09+6YUq
iGGOYAQHqkrfT4n2VW8edZPltZh0VlM/qYq67N4A1Nfp4yFu/o2mIKx6hHKJ9e3j
xqykIUcnDbqrvCQ7sAaws7sdUvirgOszvlnPZH66KhCCZFlN987q9yg/5ucwZeoK
UdlchA18ZmHuo3095xU9K6T8eayMMIYpa+Kl2vZBEIjS8RD2BqdybqQtaOyv0+AI
T7TLS3G1XaV+InzFBfqgxke9eZF8MAZKnvDT1qb5KDF4cZnMHOueGmIdjrhkqZt3
VGvJIyf3jmUmoQuU0ISfPVz8dVK3hOPKjcdq5R6W6p89qCAdxty+qDci36pz4cQm
ZAi1LPpV8Z3j7k5lm8FLMli7PsrQa50w4ZhcGGNMHZNYiUAbHkJDgUmeQHovrY0/
8VlNpQU7a9OEQAL2K9Ij1a8ft315+eygaypA0Qf5zsaIZitY23sEpaP2ObatxTsH
dnrRAQcBVX+ETR2TTlRnr/uBmlJ7Pr6aKO90sg/TXuuQC0yfcQX7FNfzje6wO30a
67f/Qj2liqwhZou+AGnw16vDcY5peLqoqXAPVvG+f5716rLle1IE5dL6tp3WvtNy
GixN0ugABCI8Ai29xux1mREb9wjGB0UUkM8iev0q5QnuuZThORH6Dcx47wq+Tj2x
qdT6U80ZffJL5KLuE4uCfVQLvqyNIEVHVhJXHSl/2m7I4H6W44n4+1E3jFIg+GZC
sD3nfeIqMPd5iCJiGbb6+N8llSwLY1J8M4W6/CqK2oJMqTXbpCljKjvyU3Pf4ijt
imkL6/16vWKU4xMAX0nKa0IP9cXzbVvkLgfo/x5wQwGufM7HDiYuMVavX4KMwwaq
6B2A2alSB1agMevPZ4b3w3LvIwra6iqy1nnpOYSC64ULXpp4iQ37kKQcPyfYmf+y
bNRhWpMqQMXuanvCOi5rxMPwDKV7UtNmeu3soHBjkhqbbfnSetE7VShyT257LRRF
uEApy05F9ekYirlQ4EXU+7WZevgDgb9UsLxA7YWCG7MUwPbrIT2xanWx80sCbW56
PAATWagWCZwzaazhVYiUFNKFGTl4SEW8LjlRg2a+zNKJNa49s8fKajxSawlR8iQQ
9t6bkuMhW3R5G+iAP9r4LSvhZK/tUG6FX2j+Dcju/ipR0EK/Z6J2vplqzX8FGjwS
ekjZqELZTA9MeESb7Ig6UW2L8tcV1q0cZnVS6NtZVMHP/QU/j9tQSyL90Oysz8CM
tiW384k0lw1mSfBCqC0OUZvItgcZZoVu1nH1GRW16FJivk9/RDfNONWpljoikPyS
fldXzZyn3qeqDXPYWZqGii7JYgL2fR4CQ2oQ3Ekm2l3WKkWUkw1YQcGbuIofuCq9
JCnFccOpIYZKWe+18hOIONTxK2HiVToH7f8wfOGS0/rjXRHZRawI7OoV+MM+G9Dq
6XRnnKWcIJ9V8ahYWEkW4r5ROuuew+TgIOb7TNzzFw2zVFKaKfrvAEcfu50zxiIb
fAFaQa3l1FnX875sQ6ABBRL66w9f70WVDIuCNUz3FLALFfaP2RDQwIy6yJPxlRBH
uWNf+bVZGKMK442hh8j8ZiFfGunInnXquQoGq03MAB4tvRIR1ph/axgnF6bvfwnp
5ID9A07aO54C9xjjZimBXIGEKNCKHmY7y8dkGsjcPZ63XYFam6QS6E4wXndao7qf
xzz+quCMaOVfslx8DudlJx8ijx5JXW962pI4OlF9HnyHJzC+U7TYn/ozbdVupL6g
+U5ix0FOQEa7lynqN0krPHjv80LIL244vIVauLI3J2chsqxLqJYF9NDwWQqVb6m0
kbDuNnuDbOWL2Id2LM4SokeBUSpezoURYUBOgXB/NNTkLOefBOH2++/+Md5/50W1
nJImOQcSWN+MWqMg1P8QdqdnEaA634oTigpY0G7Gt64xoOVFAmpw8qTsCARnbFv0
SvUXdAcaVJjuKajR1pa0wRl63qfrvfDnWSll6u7KENS1t2lFc7SwUH8Ta2raLUNi
7LZp0b7ZEiIFr/IVgp3zOIySd/CzAm3+Wav0uVwFShMoQXEU/+72thyBcBFYTi8R
37PM9sc/Tf5oqQvAQ5FLc6vc+65f92SC8S4V3CN+DjtjlgKvigUyda6AsKNzSA8I
3MdV7xYmT5G1Co/ZAQqEwDm94ZEpefEvNp7Jnr+WLy7XMMmP3FQFM8pfzx2jqDpV
mkH6j+LZDCd/mU280Uo9tK31LBSBYulXE50Th2RHU5rWxewKQbaFN04qh+5ToJj4
54AUV/fVvD4nUCH2vmawNzbTtEOv5HAGtQUDunIs4kNB1TBlWQcB65Wbptc7KTqo
skbc+rHB6Rj7tIjA/PNkrJpKQp1+iSkoD+UdzEhsN2+p/oKwUt0iUNxcYLAoyFEt
tRUNY/jUvXQJ7elgF+U3UGF1fkmJ6+TMfBOc2Q7juaDnNdOrwZw2pyAiYiA54MSa
O0SwAh96Sw24yF8KnyflDaGwizjbuAIBaD4zYlOQHZOEnUxi1FwR4jjwvWKRQKMM
187CWKSf8OXfOuK0vbZQ4PhHcZlcF07ouQijMqoqWfwucHJ+KjWpcSUfoJ5ZYTd8
vpZLKGhUDmdVioeMwNSXGCMFV2BXFUcummGYhBiO5Y/6oU0n5AqbWRuLfPG7jUA+
Zh/eWb/LhoveLdDFvsAMBOKEIUbi5u2AHMYV/yBWforo0i6riPBVrdaXInvLWqTb
3+SoRvXzZcJeSMDGLWav6dgaIlL8pagiPBWYhGKf9DWfrkyLOOWFvHGm3+quYgdr
pRu5SE//hGLNDxCr/Xmq5lCFGhi3KgPieS9LM2G42kMFIq38vFF2RDY4hIWriv3Q
iEzemwp5RKEzvw53XoaNC8VQtZa5iWJrLCq2Ko6iFBy4PU8q6YKMxQaLFULLPKhg
yCru7CrNFJQArNo5+OSEATN1klx7vIJuBsTTWVLoC8mofhYGimJ/UGYRZsbLPdMY
xL7ada+gHbXZrQBx0aFgDaSQwVUoFIUMbesUIcyLhYFCP+V3mAVjZtZKvo0iRGvQ
dq0Z5eXR0C/0u00k1YjCvQ32ttlHiLycmWKFRJc1plQeV5yP/8zJwC0k7BAFNvaw
KqpQ+CLmcB4T971p/+4AqE8v/oVuiNRJyMTT5xo7dGKjZsifuTyUVmtlSuonpCsh
xrr7FcA6ggoR4UzYA3dIXfkGRZhogdt1PikHPwLWS0usCDuXK/UJIVT86YMX3BxG
RqzyDFgdxx7AADSEyP3MZZ5PQp6Qf80NlyicJb4pVivL+yl8RIQ8CMSZKy63N8Y2
GVc61zQpjDkzBdMJkVkJYEeumq5DAs6UvWP+GHPm0P2X643GKleAGX7fxHHYmvH+
EP4UPbybs+6XgguhiLWW7gCxjwSR5j535VXqFsR/8ho48hOKP3nFMPnn1bHTWKQM
T/SFhNN+dtWYkkSmD0aAl/bib2oNPlCIY0270X7tcgaP6EEkIlVIpqY9KRoAmq/b
mCiDNEusD/bS/TzvejQ5g5CeVEer5D2XVXO0HJis3pdd8HtXAiaN/GYARBpOk1Is
H3QGN0j3aNY0FmPCTy2nMCbZHZ2ZeQ9T19ldhXBu4ELEi7kXSeJIDRpvQ5bPCi14
/VT21Nn3s727dMKmPYgeJdbme2T/KwbcbPjmhEZZH73Wx33LqcoD32MkSqHWBuf0
K80m0UUqjE6ZtNTdtLAwHp+1jwW6N5eX8B3ToRLOT58TYSG7dWX2UcE5ZxFF6ZHN
dO03gg2A6amlmmFvQ/4QGUVlLmvw8SyRHnyP1ApoAUwwPOKl1CUT89QB+Ll/87E7
ZZOtkBxoGNrHVXpRarruHn82d4ckcA6Nh2izYxgwcKMe3QmLWLAcP4rEM3oP8+PB
jpfWxWJl/D3cfNpZcsLG34La3A3pJRTyMOhPjMEoGHO1BgGwL2XPzoa0uIKKZ3fx
EoEynZx2Iv6/gpqBGtrJF/SzibeD8Qc+ePVccLWnjklYbwHcKjyxCUzIFExYgMTo
hJdApS3IDmZY09PtpEH82c42bHB8HVhWBzKmMwlrsVgC0OGbdsFaYuZLJBegZLuk
cd/Mm0KItEENWglaVaM/fsKarNiCu/pcKDh/DwJJu8ymJXPhuKie/3IY8gL0FDN/
pxnDaHKu3fU9ItxWBlHYFLWp+qCaFmXsc+D+xHajmj9OQBQVsh3H/UUH1x7CfeVB
foYSbxGUJT4FQmbgJP+lUBN1b2U8fntsjSYdLSbjNjrujj8XbfEdX39fMVBsl9cH
nDb1PercCmD7fGuH1y2A9wjlL88oekyKzq5kbWWiV0ut9tIyTAPpYsIRCtjMqBuU
1J4f9KBjiXEODVQq3h5CPm+5vT/60yFYHA0XtWX7eZlimNKZIZzqd1n13SmjRhxc
z90FzigULqVG0nyv/YM7a/BeOYk9c83tltuy5GBT4SG84nglte1c0g/qdlTLlAKl
lROFrpFv4VTT/u1fzb59hDwDvc5hJxU1luTgeBGit1QMamu96x0K2fyc9I/Nwm5E
lUX3zl7K1KnuVf12L/gS6MDtj8S1OFLiV9zze08ogf0m6ighVxPYxKsAsp4uDLa+
ttvjTwGEwp3ZOXRxTEPsIr0WjuykHHFBeNm3NZn8ufx/SxYlElyrJrYC5Ci6CaZz
OTAmoNrifpfsRnGZMuzZhek5rwo2ZBrnUw7lCNHAJ6lUajbUBHxEyqGMmZonHFGG
tYa6xtGVfJqyqHTXwk7BSkVDjw1TJ2rP2ObjkQGYqqfaluQgrw3L6KhquAqupHqj
+l2fHNoWKDLFh5XTvMdAK4hdqzBAVZ9DSpy62pk0cnfbSP1R2Yga/pT0dWFzmer+
nLyfKvxAvISamm2hNNR1An0r6AD5Vh1KhzLpiNrOOdkc0qtKzZBjOpYzyBO8Hw7D
5Mz+8yab2IcmJucK0mIiJDZvONDGdB5BAx5BF3S2aAQsV7o3hkadj6b4UdHvAtTV
WBKxRD9Z0LhF6jp93N/EWRDfVTYwn2ZGGsD/EBq3CVVBQBVYhy+Vsea341ZAm+ow
28+zoafrHcwX95LOAAq3gMAWdEJq0IkxSHULjc1/pbWFsGxdr2fD6oWfcq+UHbsE
wvT/yhpBF2/5XyEAl7IvjfXD+wsKmlIkObpsINDzd7bV0U/lopsFhILPgMEt87E9
vKEeMweuUfG920Jt3NZZg2eEyyoZvXtrimyCeY0NOpbfzq518zkkUi7IWLtNoCcR
KYKk6tsUj+jvHpHvYdqjfx6gV/VCQAFpKylaQqci4lnLXM6GrpYw1EI8qhVZ/nxv
WjxWlOkVbAWa8jbkmOE69jAkkWvr+2AimXoOCO7D2xbYJIWcy7O3xsTanf3Mn9eT
gMQFTBEo9R7FqFZujsE2TzwqnEhN62Fw+qlR11YhpSxURQ/Iq9HfQZThZzTlAv2a
JkKiOlgCcE6rfJeq5PmZGQDg5jrYbCjM6h1LA/DVahHWbabmqld6TlEfu1wOqFRO
kwycmG1yGD98BtuPzJlxmeVlm1RquDpYzSLyNOrBVcNlU5DJGCmrrtt1UZjlwBgw
NWhU45gGe9ltg+uXjZfZSCqizjMv51ldo9QjpMqf5Oz6XdvokeqZN29ZtidBZfX0
ymFr6DX0eNWmdhKUS9k7HHUqfuyOARyErbbn0JTLuMTHr0DQk/RdpYI60LFQSL2A
Yyix8Szw5wJH6m5zgraKd5SfXVBH2mL4WQgMHywOwr/O6hZz42WDUNjLmbCdORAO
DrczxAMcdSCCbMcf3na7ykbbV3YUX+xUR6fdgw4G4is5UNDwu2TL8cDG3sAvEVrP
RRQBlNS10FKMcfwfY6v8bpOynlfK098tDmgUlXhICzYyuT9MO22gh0C3pjJrwA7j
21QOPLD7KCx9X7uYS9M/UZ55N973hwVr6eoKlRptYagnWs4h82iqldjt5A8iMe9s
1L/1G0fwP6349T5EQadOqF6WchJGer5GO0C4zrOv6fgZkHcUxrQliCCqfrxzd+la
XDxayIooek1kq63tznufQTIFP53L2SiQBCyXpfGtaP+C6ZCIxO/Qaxt7z44Wn0B5
MZO6RITaCFVin+3YCmSbMJTxivG4GxwkcdHE5fdibVl8SpdBLlyHnZO0G6eri9TI
QSBLWgi4ObZuXza2C4KQQPNFDlfTwrtDKXZah+1efhbs5Gn57JI2Ddr18Eqf7Lfe
UwBCeHZreM4G5iwI/3KocgR1p7kKyXKVffV7jCH+wm5LImudivE6bUt7cBPEfFCS
45JyrtQAMiVk9e+G7sPbZMXs9UfZabKCwd0H1SfnKR6b1ZEqzhfNIEL6jXSfJqLB
Z/D4pBCh2/UlVp8mkFrd9OPb65cQ/fa7jA+adELKmpo7EJKML8dfIp4Mr5TL+H0P
QrBBR9Djfj3HngeO2sgLFJFcJz6n7kLXT6rRG60PoILXJJljFU9p7YYEycZ/kWw3
nvcQlaDkVLdRBzjbDoA6aUlf9qyuTO5hS4f5ZoQIVijgRvtPgTo0KxNp9crwRKj/
wVX1qVbEkyiexV31Up9hpHzsG8gbP8n0LOGC5ImUVgOZBp246OVqbn6WHVZVeC7V
H6Zp09dr2GGJlWDmjlrNmmJPayF5VcjL4QIlNzLtN7kC8XuNTx2Ym+WdYuARpsEu
dFSd4lCJHWDlsy/IBIs+L9pNLkjbkcdSmiEIKVQ9L1Pv/nXLKeA6D6oTkkVKQntF
smJ3Zndo7ql+fKFVFA13fzQyWPDtbW3Qfuiva41SMKjNUXgOdJI+SMhN4pqlgZEe
1cpL8h4S/SG9b9jmB+Q7gZXKWjIJjIw5JIa/05y6gi3bZDeItwj6OCGs/E8K8cq0
4QL8NyWcvAUsnJMRkDySXiFlz76ZTiQ0nf2g/cjX6/xW/qEERNcB4oSEwyFzX+pX
iSMe17UFZy19MOw0D1bMwYQlpJK6+gfgxMhYOyeTsQXgCgGP2odasBO4FJ0CwuSu
oLoAMIjfNLMcCvV+QrP3gelgd/K/g1AjjWHr2TX6Kh5dni4FY0H962T3TQRmMWMn
nxQILqzKr8XpR9CB9rtRXxbK+F+txOPhNCYVcOhs3VZqCmT3RXAMbb1NYvJCGk+s
Kj6LFp1PLjn59QKmc4JlFNklJUnIg8qfttA1fT6BXCYndzqKe3QvOA4pjBzuRb3N
iONOFIXAevHmHZglD1Ye/wR/5daem4A3i0xcOGF4KQ76hng/tX2h9fXrqwnz8kFy
+K5aSNLYhk5mYJDZfy8k5foRDGKRvlG90B1uSQ4/yxrCkmMarQkqzVhAvcArGfd8
AS253j7kqxrB8yUifij0NxO2D0/Qv5EkiaT9JSh+7PAdpk1QNFevnbo2flyBaEF6
pUDd37EgE5KKqLpHvJcUyNny8E+u88EeeQZeM4goLKfi6MYkWcR4qH5m35Kjnf4c
rlxpCPvpCG1ZYZiWdmA8YY1Cq0MCsX/5lc3gdbEJme/dL6EmW1dC/AcJoviPwNt5
HZARf5Ip3JwYFEv8K9n3YM5/uFmxFT+zR8mD5JF4zLbM9YlvNHENJVyScOptWhBM
ZsPZAD72qkIZvHxfbaMYbV9yHwBsn9ytZaJhcq7jLo08r0mujGZftO3P29hOJZqb
QAalzmFBx6W9AP1ZajM1NCJ9jupqMF54zjdEzHrfivgz4eY58Zw+c0eo2xS3hczS
d3+KbjH/wc1JokhjPUtSN4bzXCNxulWQ1XaAy/BMHJ4tpz2/izhftalayZqVQos8
afNU0IEkbQDSWrP9+j3jWY1Re10GbS60jEFpxm4z88egCvanmtvx2oWQSM6P8sE0
b864hTB1r2dFvnDK1+496gqcjq3D1MS4fMRCGOxkgZnJ1Sln3vGM/MZeNVLLjXz+
xTemi5pppJ0fGKBFxZGnQXGEG+tQoFR7W9HilJNOxehh7o35zWDO2PdxpL2pymfD
0FaPKHrREWY1J8nXREH8GZFbSoGo3+C8YG4DU+wXCGzFs9uzxf/VYBWQQWYQ88We
x1+JAECGJeBv+DnQq+WbUxQH5iKCgnEXnc/jMafEp0Bw5aBIdMxSus0/Ncy1pZn6
RSDIDopstIbEhzkY7XNMnES1JYKbn/hUIhmDmbOMN1mRbr408dP9OY69s+PuL0xR
spfJ7XxL2AVB9oR3v+Zq9Ylz4yU1mhJFfDDmHR+d48CZ4en/secNlc2r5x4Q11Yt
ekeKf4WE8cjDPr9YlYwx47RHZnHhf6UVMfMxEkCqKGjLD45ZLMPF4KWFoN5KZHwn
4JrATftLLOMoyBFkZUFuxBTGeCmU20eEOUuE9Sk7jRyniurln1v1g1U++BonQMgc
H5t76TBz2OMicyvshMphBJzuUX6EYgXgCUAJ4InH0uvGAa6jvQWE6twMopIe+oSy
GKZAi/ZeUitKV7J0Nns4wsWBaDneBty9Udm5Pvmi0QNZ/7eZA1EObLbUUihAkAv9
HyfnDREGD6Ony4au/23PQazuGrbdk77FvWkAT3lnCB6aUYFYC71maVyCESN/2oyV
35Ty/lETADbOJ1EU6sr24I/xzYAWqsibwJvvT8TOmWITHd0aW1Cj3SFt2hv09tHY
a5Sitgpxl5wIO3zkL/Ag/b9OC4YE7Pc5HJvbnLyHSC6CtaeBCpJHe7arNExjbLys
oZEfpHRmNa89duXHIPO0XXRcLRVQIuQi+gPXTvZGLa6qPGBcC+xmW9vKMOsOOAJp
L+d2rRWATxeejswSWlITVXSZHn7ob2FoGPrC2xOL1daieBqG6ean7Q4YxDYaNfL7
nO8sGhsDNb25k9aGwdLJa3yDo0avmW5BCHGbJjjxqd9sKAHVkIiPrHOf41+VgWAc
9+piCcaogYJLtDDXGEwvVyt9kB0dv6LWHovvjgR4FypJtN/W2vm+KePYuHK/NxAe
VElRkBqTIfZHWWOq7q/jNUSa+vxR9xywAzdiRtPfoFFLJG6ymFNTSHK5Atfi4HDY
6eVRlBzPCAFif0lzDPxF9xlIM69VzmhmDKFOWPbnHubHqm/CrXOhYCHWSWRttG4n
2ngeECh5O9lovTfu+Qx0ygM0FYb+ZRZd2c7qUWIzImk88XMMOlBQoN2P6chC1p2K
34aP80S9HZBV1at899GiriABwPwabRW5VFrYDT8SdDfVj/nwLmvPSaaImedsw0C9
r7iqwOUcvHJIDUUdAFm50rf0wUrz8euo15BNLkufMvTWO8db261Bf3tMcyVwRcJm
54/22DpcmISLK72Foz8VuiEUE3M4WnAjy3F962A1UsV6FiQocwzqEXC2RnvEWK4+
Hm2FuNLNifEH/ZmHdtiAK9z9ikXGB7mF+L3Exd0VYTijqUQ5cq4UT5S72F22dVPs
BDqThNwb6rNPCgb0suuVIB9a2sm6gXyQ957MEokyS5NJWWLavCdgwLwp88qE4or2
otvU7RBFlNeDMdCPbfqt+CHfBVfC6JnqOQ/I6Ye1xzN25cXJ90Jy9o8ywOj1qccO
JuyK2zjmaVmA6gNmH+tXW/4aPF1MlNrvyJNXgjMqtHWNLipD8TfcbKOxYgYOs2IZ
KmqgKJvCxS+GIpC3QkUNcZGemPWYRlS9lh7pk1YLkOtFQ0utAUzD7K48o6a6SwYY
KkKhuSuRX8piNaFdGOm+y3W48VAIkC15zmCKpbFNy0jYmFMh96DzA8x62IUHOHin
oTyDFqoN06n6BZD62S9pR5x3JGWIKlmfFa/J340lRFwIgxvgv5otuuPB4vb/wYuJ
MxpmoW1E2D+qjGDwHLtwwlDdq/appczreqFBIMgGA8UXPtWjZReZjD1UOeVwNNuM
QoT3Xie+JqyI8AqZHSi3h/u2qFqjthQUvUeh1LABbKzNzq7ssEtE7JLUkj2xl4cE
CztG9ViMqAkc1khLM2eFKwyn2qrgltc6M9KSOr51RCkd/NT9m4Br6h5WpRwr5LpC
nmGIIE1H8+f0aIHbfVYJ/uEw67hXNwM6z9s13kiximwd9lw5TNlTc/WAPa53+N/D
29SGCdX38PNQ/q5om5gMV45Vk5s5Rrv0yLkJ/o58tU8M+3KTYKegMVsUOku1cEnp
3ImL+T4B+s51V1f2TLfFe6AuAiZXlMMIUtVLk2XIQB5qAgoJF0MWxD4vXTJ+Cwg6
vXH+vqMO3m2CgGxztwnZZUX0djNDLskzXoDfBgORMLoqj1fCjHT5wNgU41smQxWY
ToUqFnB2gN59IuzRvVDInILYj5tbGHmDssmISNmUwNJ27/e7741a9d5rN2O99XGN
Vy1pwuLekJ7r8VpAhyE0jwpemVLvdgfWj5JnSSEqrQQJS4c8raUCoTTCLm7muN1c
QHhW/k54qzZmXdSQHzlvxTZCCC/H9VubPs/GAf0lrBPq9aY7UaWXVC06MMZzLhlQ
sbqssJB4M7nkfgSc2DxRaC5oRquI0gM2a4HNTIRTLYsG7Qmwu5bV06JRPHbs8tHE
Dz1uawflzn1vo7EGdrQTs00DEmTuKyAj/WOfcJMJb77AYxh5z+1gl5jS0Ectd081
b8HHfpS1mozu5fxKBCSLhckrw7mKLh+Mu709JCsWv631bIbKCxRJIKyL7qbGbR2i
dTalAFjGaAA02ZZnuBvaCfWubDchYiRN08GW6X3M3v3SQBMliyVR0ItNW6eFozxk
loVHQAezYuXRFm1yIukrF8pEVjRx/bMmFJr2de86ZnXV5Xy4sqlRmBnj0UJAkbrM
aNP6Zz8JXyKbH6U9en+B22Va+GF0BzU0+NQnaROz4Ixk2XqAG2e/GR6P6GaLijwi
dUGsQVHQpsGbbw/w+VojHdu6yflLgWo+V/80bxaRmVJprTQIXSci0tUHDfjJzNI9
qYD7xD0LCb2AwntbcRqAAH2LBcFYSI4wH4eCZi+lSEnKTQmmYZQoMrpgCdjxMGeq
0gKl38wasV1pbaD6d2IJ7KgXhXGavb0JGYM5iCU0ktHopsgTkceQApQ1vQK6Kul9
W11e24NJXmb5odAQBBFahppXbdD/xHN3KQQSH6gIs+xtXs2jYmqiXpoaWEggfYuJ
ZJEDTAllvZ5l2HHtF3qR3/p5cyiM5FBcuVelDSN4KFZD83jznTpK1HSIqr42lqmf
Au5DEW98+ua4C0AC6LLgsdqsdnV7uf/GiHsvi7WkdVHIa/FzmSaylqc+Aplh9gSk
hPG1dJkPHl42A1zVImFnN2MDOy007FV2ZOU3Ty/q/5rD6lTo6Lq04OqQ4qHBXd9r
zdiiafxp2RI092TqwiYwafm3Bu3vlaq7tutgVMv/EqOEFxOxap2/RpQeygUI25XC
4r6QZcNq+Y+b8h9B2I2/Dzo03bgLMArv33FsNS59/aZ73HR0/PeH/rhu8Lz0Wytk
BhTUgmPyVkwrj26k6fa3DC9ZkdK8dGTF9OHZnOKnuSVNDVYBd6Ql7TbuFODIHpfJ
Fh7Ao49V08k+Jn2/yEVb0q6PxorQnSUVj6vvSeCCdel5CA25NPUJszsWiS35w/qb
2iy92pYGbtgC2S9Fgf5amrxiCGMSWlR0MJCYDHwUJAavlBi9v03WDZ5TGM8qTjup
H3NRVmxRU467sgAPNP2aA3VHkCKTnAoI5IStC6fmDfpagkA3r3F5AnUP99miYzGq
etxnmhMvgNrWkOa+0NimjyT2D0i9jd2AqfHIhJGC6qh8VkrrHneIyNKb2ERH4+Ks
dp53qvufdY7QQMpX3rso6DFtYJu1dMggkCgq99jxoKgU+vRGZQAcN0/+GZgaLwBj
GN7TcJOCjHlNNV2b1xUhCuqIqWRpY9V9B+umxO+BsHK61+C1fAYOSaZb5dZQLcTn
gojFCMn8RWhkt24ebqgqAwY5Y2DiQqBLXMjEKQHhcKefh/fet/PEdPISgWhyR8jo
/DJUXnMb1byAEtfXfboghHXNnX5A4QWundJKiPpQucl7KlXTTxsqm7W7wHEYjW1g
uDa8/pMcmOL34DepF5L9lJRQNNIGFSW5X5UChatN1RwtX3G8h2Mf8a6Jwlv8j+it
jrOV0A5ci1if4xtjL8Ri6I8WgWvEUZy691WkJQ1eqQa+kL5S+090rU6pk6Q+6hKy
ydN+UELpu9Q7aKS3chDCn3rZV3bVg2Vr7Th9H81c54Wg60ogj9uVx2jHU9ZR5xG4
leSARbviikeIixuIJ54SZiXHsRe1snhqWQizV3ktVJ6iIF8D8+UsiRkCTptIU3f3
3QwBJPSWxacr9rHdHUZlgsaVkeCdYFDy5dim6sDd2a+QDCrxlhTSYINz3sQCE90j
Ce6piFoTmvdoGmHF5VsqrZ/JVEFEhP7O4Lh+HOPVbo2ou06ExJUGackVPjkwApuj
J338LofQwbEJjnNQDVcZ/RKJHEVYd2pR+BJvAfwc+9BS+ka/rVWZ144pXCxIfuwq
7TDKIPJ1a46KMJK5XP75jTEm/oymj6eI/cpR+NNYCcViNQhVNU873uF1BiHkPmks
9CkrxLEuXMlfBnKTZytws8EsKr5DFJ1ir5vVNCFhxgl6G/XWOvobNZD8V2W/9DBA
pJGzHk2iTmELUBe5G0iT2wZSrmwLpmxaQsrWZP1io78V8E/hcrYh+SXybCCY0XGH
DXsqJW1BPw9qKoJukJbc6264/xWwRAgoJyBpruhT2vZ3FP7PQduX9ci3OhZPN4QW
EEm7zYvInZEnOtDLjbRYyyE7cPdZZcO/r2ERGv0F+AHSWTxvqYtzahSeIAIRvv1X
/1R/ikPB0DUSqQaznPDV+btGTrd/WMFGoP7T0it6MNQY1xLxbpCg/7rYSVbtUYPR
0KqaHD7grKyWHwOs2C1IlzKTEnjoMg5HDL3bfIw6RtvCpObEpLg592WaOyYJdUT5
0eOzBScDXpF/x4kx8nuxbbn8ZJhpirxDStRLRTKZavrMDyM1zHmJPk/h/MAaF7z+
+CwDniv0me5nigc1KACChKUMhR/8AlRY9Bl0kE8k7QjR378e6IvMUG+pFfLg7bBc
eYOhsVuZhfJHjse+B0LXnN+mW5t8x6dDOPAPuVwWr7ytDLi+oPogN/poJrq3VJeg
VdU1a+Z29MWIkUs48AEZU6IoCTWPs1UjhU4PtyllHD7H1QMTQ1jl05yEkBG6oZlm
wycZKT9DVNEmLI/VmyJM3eUj36LOAtQk0wRiXo7qLaWWOOW8Nmz+LDA/eAaYjO6s
c7od12B1H0R6isptef5Vae7PiD1Gh3EBERC9UdkzlqFsWieUwZRZo/b771fUfnfH
bm8+BOnlfscSiVirY8AtnCzSwkOlih35SUlIOBe1t96NA8wLADzt6IWdj/inr5EO
RgKjLPl0cEqR9a5OlWcYDLPYiLKURvrhPeYlFgGjjd7R1mbGTwrieN7fol1j60pG
s2zIIfQa6H30DUq+K8aCN5tJ77Adf44k6ACE8eX57nqg154B+42dVTr3Zv2GpY/s
xw4s6MX/rcwY0seIPmaqz5xkHPP6zdNthJwjJD/T/DSwSqGZgZ6LGBFdabBfs1MP
zterSmfIy0XgyPKpuGVmZe2MckVQy4ryVglsFssYxoVxVYggedMsnKMkwdxUIU8P
sewZGDSYg3YB5KYvG4cxk+c5iEHoCVYMsw8UdlrHk3s1Vk7rhLVStgsLDZB62C1j
y7HOWaXW2ELSCOZJnRBiaSSqX6NQMoFwF042HHP9IYp5coF3vOZN546rUpgzchx+
YMHUhp5nD9S6419KTzsBb3uxsgHLf//DVOuTIyBSZXX8z6jblPw1Os2jru/GM/5J
JXsgeU60C2koaoP08ax3I3kd0MWpuCuIfOdW/ewrovEVVXIWYDCYm9m7i9XRwr0s
axIiYPeqRU7f/YXSk7zUGP8p/jmqHNyov2MaB7sXoSyUd54K9ekIq9zrN5bEth5w
qHXOzrGvDxzEApCPhlxhzHr+RU8ptPTlz3kV2IdZeoGJcQMg9LRzLwDqxhlOwt8K
RsKVbIlAWNZp91D0bIBHwhliWmo08/A6tiRC7DzTiOO69M7KGkyaBoXZjGiHBtpy
2TKhcKdkP02Oc8zTjdK9w+pdU8wKxPAhaq28Dou68Q6PYxfv8+lKddvQcTpvE2yX
ZLedaF1ASbyKJCgseS+ZM7XYrsJDOx02n6PL+KBrU1fBcLP18atSbTLaxYyMsf3l
5LA9JSA2im/sA3K4adUc8OnQexTMXVIQ44HYJL3JoY6WAQIY+jDZxzZE8gTbOvt2
UL2Gtbj1qwv5YGRfUbOzU+QYcJZNr9dnwWk4Jt6sABrocnTQiPN67ncTctQjvQg8
xBzcXc+Mq7Vwf1t3BEitO7ebPLIG0RngHR8WinssMVQnVmFUHLLEl5iSik95plPk
RreoZp5Lb3MMoab/Rpl2emI5bcQ/rKs02n6GSxDIqiebGoYVXipfvc8VhqHwE/H5
l7NhbwvZssHtXlHd0GM6etHTWPmTWnnC1IUd0oxW/0IJSL/5raWRVh1nMFEHBbUC
JNLs+ZNDI2sSYN1KxdXhDKxp8gSMtc0pByi/wNoQ5NmR5PxBg5OeLYpY2CK/sE46
iUBlAjt4SXg+SiGZlvLkOYM9dmO8CkHFb+s8rJtRdu/GbH6e3cNcHdPH67Mn7V0x
30uUlqmt64eL1zW1lxp3EeNno1R1t01rmv6JjcvijRkQL6T0rEg9laC2VhkXXnSH
pWakeD4t3H+UDF/yIzm2o/Hjy4+nIMBYxOZSTRkaG83bSwETSJMAplr1qh9cdSzS
hHe1+2SQcgNRpL0YYN+ieyPVe3RXx8h32+cLZonDUcKy4I/UrN/Bu769tJ5fnU9e
ZXpIUJu8IxpoUfNNj5YLYOsFR8e0jUk/rWB8wh7Yj8+8O9F52g4PK925bRlpebM0
l+G+MVY7aoCPUQl1+jGZ+yKZSAfv/5fUmCJLBhM45vX+51cn6o4AdBxj+Q/WVUSO
H1Wg8zAsiXpRezoDY4YY4xUBaVF9F6brmMgwXejX1lZUCUo53vBhSWhw3eVMFlqz
wgIK+8xGNRAQNqFmUIIqUKmlsWVc0ggIemseNM+fD+I9FwahW1rbQzmpxlYx/wcY
isStKdqZObcj5XpfCZ8egQ9sc29+2kgxEA6G9lpTR5vXoCTYssgIclBKYY/q/ZrS
oeAAgkuWQtyDW3oKq9O6EwuH1rcB9CIiNzQc7VhILwM8ne3QZ10ir5QweQyZxeCY
yHp58zx8EA2Zrd+xayq3a6xXBl96x+flYRF/K/8IUpr52jtWaPTkkvivrn3CpafP
HVxlYMuaVlSCbXqY8/ZtRSRZhySeU0BIVt0e1KqYiq6/oUaf7tDSmgGBp0Yrrr3H
5h0fDJt4drv4UxkPl2olHPeQJdRPdOYwd8sisKR34Z00ub2lIvrO5jC4ODKv1NCK
uV1H2LXero5b+3iQ4rXABPFc3j9EfXyHPsbU8TkGxezuA/KJxtNhP202YkFRt9k+
bF7XICh9W9FJSA6MqZ+nh3hi2Yb3Y2JxhDMoD2PLCA0xXPUTrNsw0EHyyBf19wuS
S9JGBLOkGr+jau2Miw4dB5ZuvHf4qcTKt+PRqbXAPAmUf2AD5IX+03J3a+UxHQdz
pOV8u0jjUs6FY+yHJSeozjBcnjaM5xTrVeoEhwkCVoWG6I1zp5DA2kXKYc4qp2Gy
UYGa1aN6LLwJ5xTnyaUUHBFQreAeIDN7r8Ug9rG9w7xL82u2THIipQoFPx57INQ9
ZdxYCWR/uOfS9/iCdImU0FejS3KeAUux6KBxyJGOoTM8kkfbCbftpHA0QcXbqkOC
k+ERNZNQckBLxd8yupmTOL5K5bLFm3d3t4zDJidPXAZQFxVSf/w4vbYHR0tXke//
ZNYtM3ra8GTyC6JCQ+dQmOrPfMpodJ+BX7ZeDntXL4z/WsQMR4Do5pdri5P/KzRL
1GKilcdmVT3R6R2W1EzU3JTaDqx3kOL8/ZlUOwDmmqynPCR7j5V8+fvTfPWNO8CN
INV4AvhSVUX6jLmJlfD9R6crfzqv6OVsQlIllbvz6mwCQfrL4JeSECd9J0oH6w7m
EdEKT81hkl6W2E6DBRe9LWghPDz2kmPxkmrXymOr/wJttJH4LEKcsWDyGFP2tt40
sNbETW7a4OxtrJp+3V843i8Jawl/VuB/wZb7p3h9MlAZqx/jZvyPay6EaBZUowql
rkWRVGbmv5OV8A74m7LycelkhWYnEeT9E8mdewuxUlWtUfqpHt01nEtM2k7UQb2L
4Ltz+3i0aIxEkIBTDENLDAk7sF6UQRseGzvuiT3F7lcw4YMJzuxVZwGp3LKAvz+T
FW4sRg0e8z/b1I29EV0yTZD+PCjG7XYuLwEY+vntUlM/9k795j8jThnZueyfbgWW
Gf5lMyLMa6cItdRIqmghpiCtYMvazjC11ROKne+8P1rK4ufl7CqLFe72Zh3qDXuf
E3wLN00F+fZB091f8uCic7KXs23ReD7KHlVSiRA6sQxoQ+LEUfQ/EmfFvEc1LfCV
n/uPOKnjw54AjBnX4Fr2VUoQPuP2HWCxfdgQnoOHQ3CxI9k+ZRIsw5MdLUjndfUr
GlR2Hlv8Rh3pnIrnlmlAyBQjZBVxsNASPP5ccM2TpLGCF/tnHAMM8lDL6m5Q8Cs/
uHBHHgh7M6u9pi2xrqvnb3z+7F/DzJzZ1N0VTY4tmEW5AyOFU1KwDBVrL/z/7z6a
drLpUXchK3krf/nkMhOQtaKE2aLCDJywifPf3QDRdSfZfAh1Zk0wP6GeCiYT90zp
lBo6yrJvC6iiIKVWkh2wrdqmyfQpmeHJmm/jAZc+/RqMRjgaa+6K+I/K+cA0XOaR
QLKjRu9sDFpGMw36ofbBgE/eFu/3US34EWOFAmydsRxZI9im0oorAlflJr2qdfJS
+qN/NTMyaTu0s6HEtE3XW2x6K2NQpiAsFd/3ZnjlJ3SBY0FA3fcf62yaSGiPJHl3
nRzU0yjoSWHA/E03HfH43uusFiuGMMVbRQ/pMqWesMlgc1SulDnIs8Dt7G3qE4+d
gF4MBexRqrsujbdBUE+nHbEFq+2J1fBo7xNSdSpr7PNimwucGaUaDjJvWmETS2qQ
2KyE32ZFJ7aDV3mRRkxwJ62z7GL1+kUPPYRD/oZRtndlLv8I5R95FhtVfq38prsn
SBtZz0+EBLusVcRO/cNBdQ5NRfrPfyohDOPmdj3yIaEQKfquM274BiAPwGyLE204
EaISrtFT3lNdjUawqGMw+NQ8d4pd7GOL/T2/CIV4VBeNJQ8lC429GHMxwbMJOpk+
RVZ75r1TLuK+9PRj+BpZZtBKoBQ6DNTiLry/HyR5txBAU9lBe/UzmNFm3+f3LxGM
bR2ZbUlL7giGXER2vdJCuF4vDyKpGYXd3tIed2WoPbvKXTGZQXd3YXp4ZneNOw4H
np8UvFI32G6bX7kKITIETu2fUBLWsv/Yt+v4MLRe7D5bjDzdwGkyIQv8uuoVY8iN
lrlTwvhfDipraLQDujJcqwEw6Yxda/aj3bIpnxJ5YwkFe6woWiqIHbUKPDq7eOkC
1S6JlMVyxu7oOkXFOi0WK4gxqrGLXcTAcYjxGEE+3fcmOXP9E+8ef8iQxW2S36AQ
wmKuRh3S0cAec+bveR/KzDNXRC0c1MpVWqeqKKawmK9SDgvmdQphHlgUAfcG6rr/
GPfF7DHt6Xg43dASXltl8HlKyN1UUIsRz5SkDjiP1THcZRaXSc6h92EzcRhI99vK
1bdk3taZgD0FkgffLvdfvJYTgP2TmD0Kl0PF9HA67OFdMwwZdJpoAs0EgoddzM3P
NL1Av8yLJX3nURkSGmhRL7di6cSdoYA0W0nRGmvzVyRh0dJgNp/TORIe4mvpcYMg
3FhG4YYlqQKO/ksudQX/Bjh0rUb3CPc6dIt02iUOqsWy2fZzPo01cs/vq/42qWrT
BGwjAxKvQf3NjQXoh4tvJQH/MQCa7aUmEpx35DRWrdvXDEHF81dm8dPhOLSfbqTr
q1Did2KAyZbEQcorSd1z6D4U1nK+ZM52PlvH1slRgalA29YQpyudCOSLKMskY8l4
gqJ05OnWqdP0e/BpU8H6bt9tPZRjC6JAsiD6WEljC2Q7f60kiq6BgqIVTuZ8dkwk
9AnuVZDY/c2zic8q2C8jeoRlWzbKietSGcXCleI/nDqKfCeP3TkTs83Kdjzc0OuX
VVm9ZlBk9FapoY6SCFg7PjQnnljWZ8VmDxL2qpUZirXYfZcfL6tTDCdLeHRLJt17
hfJ1QuSvlyr4eK2bXnmsio/F1Ut+mq2uFYZOFO/mefHY0oq+xkDHzZZ8vekEyDK1
I/xJIXKuYbwq+uhBrIaE61PwvhTofH4ThC/vMvMVvRV4oLceyYldSogfkDDh1jNt
itF6CdnhNwr9Ys6P3muL9d/VHyFYN6r6Nf4KkuULxGDUP3GL0N6N2apJ2NvpMBTa
jVq980H6zfU1ZaIDTbnGYZQA3fPy+dfi/WY2v018AG/OKsU+gpK/b2NubtVI+Hkb
ira6gBh88XlSKctXAqnWZAbjxOOrHKNtjfxteM+MN/i36/MJVpm9soM3j7bYYFuq
sX+s+XhynOu76SOzv7amus05Fj5gsQnK7OGDXj1thJamejpnNSAbPkRcYz+PNJXL
HuwJGETN4qGiLbOZCxnLNl55A8hzPHRE/NBfC6oAdW34S7giXq0vj3iS32Vc14Cw
xsfK74RchrGLbn9vpMWi44d4P6SdBmo65Z9Ff5RmDCMVhOf3lUk2+7zooSv1EUBF
RmngUlrOjmPLb0UhDzrIPHNqH6uxrbEHho83MTOgWl9LILFWZqsk6lfQDbxn0Ufh
fpwocRH1ck/aYyfdsFVWcN1DrciOyIrdkM9Cjig4Vg7vTUXHkGhtrkjSfyPyp7qb
VuZcA8lEOPEBBxPgPnnFIyfea/Y1WufV2wbVOHD9x3qVf7oxqqLE2YXVT0PjIrWz
vLBHuJ78bbfi8fatDNpWHJnGlHAS7V+IF1zSBO3uTz/sRRJNQHSxxE03IUaWdp76
pRvm23qjQcCZHYjn5Rrwj6ueSoegqpVC75W+RwBXpEFfHayWSlE9YU2zxSmXJdfa
85R3whkMVivAE5ZLy8iDTUgCof+bCopj7AQi23Sfoi0Y83k/NST963GOPPED3lxM
sbVUZfktfo6UgQH55aEYNClKR0baDJM2gx3I5QQNkPUogGQ0jHW2YPUZszEo75Gk
OcgGqk4CIbpayxSs+xJHAwyHW/NrAhZDeYo61UqeVdNyv4eeg/94+y7cqjfF+CP2
tJR5WL3MudXMPpyCcbwOOh0jbMlNuOKzF9U5ft2ajVzgC4rzMr8zSttM2DO1/5lx
5Eqo320P8XfSha3Or3HxvMvu4KkZVONsdokURfUAXJMX1C+jrSvlL1EHVVKsi+AX
hzlF5ED8xPAd2ld1URD723QBomHPWcDw9MUYLirA6oTBy8zVr4ZSjijZTvXHAJUo
sag4yPV5G44YbFUmd0gV/AjfIci6VkzUEELGDHK1xs82+8UoCuZ5mlk/vUOX+oie
eiLmcN0eF6CAls4xPRojPyG5OHCxFnKyXwgR3QDDM7P9vyJJE18cIp4LoWlYXttQ
ZqnfdYrxft/rF5qFWK0w1vxeAXQ3YltqtfJPTkyB/aqgmDm208cF/AsCytAOOs6a
9Ef/MH06db9BehzjvPMh0WGGMw9tIgVFkxW1OFua6hQyE45YVgPGQjslZRVAXKtu
y1YPbw3SLHfNfdWZmMgpEpho6LoPHMsuMX4Cpxp4wDyIAbgGMHra+Th/ebKeC67S
v9aDjnVxkosk02OAzqhgxgx+jQvkJ7vj1eEPqRUtu7RmNeGMmaNWuspP3Ty3tWvV
ZDRczXyEymty2Rki2pP3xpIp6ph5RqGguvHjhLUJXXKd1NaTmu/iO/7m4Wn24rMp
qoz0caYmBzsETk+M3qSLSU9BR4ypHVMbQ0u7OG2IkZUJqXHqky6g2Nq0tIthGK4v
v9+/u4u9LZ7HW5hxSPKqqLbeCdARaiywP1AnvSfJK242W4ny4J92GENtVdJ621LB
8Q2pQtfA8wD15GxJgUuDoVPmbC+UeW+ryFLhx8jlJNJjWsWojAWXC09pbjobH+BI
wJV+A2j7korvyqIdZs5Mg0DznTQnJWO4GG9zy3nmVjwejGx4kr4/vQjCgNs9/uPp
pGH+QUqUp5MPrlIB5L4HlSNsvn72BFtKI13JNT4w33guPhHINYOIzmCl9L9/W6cL
qPzuArIsaAvNMIVNVjW0D9TJohU6QskU3AfWrytcgxztNINiDTm6cAEJCKq1qP3N
TefnRKVLLjIu9WguuRNfb4swQkQgA4FcmQe0vdIU921ybPeevIUid8S9jarwDVXG
aKc+f8XSTiNpBZgQa30kAk25CZXMx1BD9B2jQGcRuxYp01waRrv6+ENjVRgiI8yR
YoTPjCjsRlvfkYeBwgx2f4ME36DcIz8JPbIhXr0FTs7nzRajkLnzbDGDaJ1I26TC
OCUI8UwpIuSYAwr0s+RKI3CqWhW9KWq1couj/PFZRU3d1CwQEEOZaGg5Bc78AfQG
cqPhT0rU4UOSikEAjSdPQjZypjxpOfQDuuBs1+Lnl/zQbE3mXpZFvk9ktTQuRADY
cEDaT+3JHGbxx7Vf77IiI76vTqfyNV1/a2bAielgzj/F69JtXuq72IGXgL7sJPKl
xoolb47of55P1vbDvJ87uEG8kyUTTNaVhnjbYOv9c1ddangIRStAa0jJYGYX6K2M
I29e66AWx4EbFeqGWkG0JyboH9+ZQBwepVwiX1MWGx7zkj0ouOasptsMoHg/3PYD
JOJkeEkPnjGRtZIZEKKtJZp/QsgiQukmGf/LiD7355onIFTzSJUELNxMiyifm8CU
lS4IVu+9ZHTza7C5DpIgjWV8zoVE7Rm9hF7poDSII+CEZvsgHPKVYVro7mYLxcdT
usn2e92dd16GHjBjCWvSYThOl1Y5ytLZnAIMTuj9tG80TR5/ecGGLdGWGTrBcK1A
zH/sgPHthJYiHVxmwDRSCo0Hofa1Z+OoeDUO1j2pqDnbLBp7VivmYBS2e7cscDCR
FWBqgGJjEAVBSMfJiz+9Us6A0c8Q8NudKe3WrsYCnI6GJ0hBekJb2dYA0Y4b7NgJ
Cc/q+csO307Xmie5D7lOCdBGs7RXJuzKlsSzcSfQ98NoX4Y+1D8sMAoaQ1OHfOKp
bDy24RSyWQngznd2cum6Sfox7iy97luUwJV1iXh0pVymgVjaVDc1nUhE/RmnWeoa
Vt502gbqbsawbbNbn7csnoTavWDuSfGZUnwWa+DjXoKUrGCQ7CXSF4pYjm/JbPvc
5CATksyc1qmEHRSA1FA4UpCbD7ceRExoPHLbKmocWsGzSWZ6FZlVNR/AepKDquYk
vuBZUNrsc0qHPE/f/DLnBMlJs58skmBeT9OmGzB3+JfZwjmUdSC5539o8tFdi1zo
9fMQH6r7ilSzvBcLu1f4Kvi6MO8OyV9CTjjIdiDCsB3ZeDF2rXTnYFz9kKV9oIvY
UL1IKPIaC21awboL0r4X8u5rhgZUqPqQg9zmx1Ss36JyCACQNpsXP/G/FmGUZ75F
DshGYkRA1moZdTySnsNAU9Hjmln6RizdV5boaXy7rpeqJpoEHMsZMs5QV2CU6cuP
l6tOUDbXyZHCu6wVO9KnFubk2raQH4FZn6ByP/eh7OsH81pcUx6sIHmr76KDlwvk
NYe0tIsvrB1WWy/qZR+En+jboAneyhBBqqjLFdiwmheOVD3xBVFYdTZGmkG4w81y
kgto2JmXG3/YhoYNxOk5JfNp5Yl2v8mJcuNVOuAzvnpq7rRM16K7H5arpP+XPpoS
a8AYRlwyjfgSPqT6kgo4V1BIlSjYaBsWYS9+WLiw0S/4zlAT9oSSrg1XBU4RTGl8
Qdm4ZA1YrHeaF+wZlcpGRcBpj7VUnIKQMBq+V9lcx/bm6lgmt+4AdO/xWntKuwpl
fDMHHtvtPevfencNjeEeEaepiHfTLluZqGthePHhb5N2OkKPzPXrj0e7TSawAdUr
qoGafUwvUJIsP4ev7eDlrVSTCleXTcFVkA6LYoo6d/831PjvuhFOflqoewYDbKoX
k022NCzR3oJp31EDGKWiHOm6KP+jr8UO8vQoA1/VE2yHjYwBCYun6BRDp5QLUtgV
nuGvZrPSGCURDMCb+G4eDsqItt2lhIkS3e86ILOZ/DHkWd9XXHnAjtwfJDh7UjW5
CyJ3u0gRtQ2Mv/H+KGpbPOKXJ+10XIeP6gfVUYOZVgJBPyjv9Pdb07T2xIwtSOIe
3O4BhMWfZ1SDfI4/8PT96hYObzupK9lyXD8z3DnCbWfbrfM/LMOajkddvRsN7v8Z
PPMVn8gQffb3rAa3dhBaQIf/j4bbzeKTjsECJBzr/kp47HqMxiMWBSNTmgUt8bqw
Wy5HqePqLfD1P1AWWBEaMX7tGgmWprr+9z4R0+3Kle1LDwk7zz/i6xXeGgo7CoNf
JEaseIJY54VaVqtXMZk30wZv6M/MntPyZCtNW8+rKUT6i3t0GLBSVoUZ/5pQ/Tm5
lL2QLUIqDpZ4LucHar+aw9+Wpdi7Yiwpm5DkrzgXBecLUufx+MfinhEwDlijAC2s
cqLRiHfQry5wgUmkL4Iw94KjunIhiMhegjkvqnLzI2wqxKaFznvxQbGGxksHeFZk
Ui5oEPgwXEc8ofg6sdRXIbE86jqZxx39RyROy63q/PehT2pIYlZyFfypPQCa23rA
tgFj8NIFEAUndzzV8th5oZMYWW2HsFa+sy7Yz8kHhYDpAGrpUCNYybdK5e41Gu0/
4jkRZh1PrX7EFwkhsVfBMfEsA8PsvV8w/crwDkuP+0dQBG/tMt1by96CpG+xvGKX
x19yVdTa6S82gRGwKQOGxb5WggkjsR0EFOeBKZMD24e0tJz/hsSMx7musrgqkM98
qhrHE/2k2xPTTh48zbDmLMuIdoCfGa8W3wmYSpc7CAnppC6k6sq+8YU5jITEjKAg
lggW/6IT6WB1WTBuJ/vTSTgbwEmeM4iuUvT+E7GC8dwIF0OJr6ueJyF3wU2428Fw
sVlDLP/LjEtxlZNaH/cyqeyCkReNZKgLVm6Bs+jkz5dSEucNhVV/E9VF6/c/J04M
u/2UWLyl6R2jLq+iIaMlzDiCesFuYj0dZ7T18u4A7vqCSxyKl1LHWA0Yf0AOiTCO
MBYBa2q1989OOYClMH7l28ZpunKyrHxnm9hA4C6Pf24lYMri85FaTBDV6shrSndn
wl3RW28yld3P9qyRX0NmHQuCsdG9jjL4Ot7RaCucDDYG18tsZR4etVISEAGerrex
D1ddWX8izWkbe3OI6p4H8qcCJBVClhugiOIrRYeiJYLXNvZT/F+plLbTUfpysJbl
T+MtKZ5eyTT81hj2x5CgNHM2TdPtIItMMZIYYS+iUZiHyw6FK21SvV+TvZfOBZ0G
eXnX+ryqsqpN6Aihzs34+VXqJOdynk796jiTfBGogXZ52MFwyTyanieKsUXItoYD
qJucl5qCz5UNHWuve6l4ZMcPSE3QPJbwzikgiCJMH99P2WkZry2Qez/PLrq2lQtc
MdYr8FRVj612vSuFY4YCr6krmEfVE++B1BnrUiZoMARb9bBEY97exj1OVJiApg4g
EJzZLFJV1+rN+pJ0LU2EuS1lgZkXCniPytjOPQsXltJ4qGrT93IbNhF/vApM7v+8
9GbL53CICip2skx4tO7WhIUcNHGnpt6X+G6TuQ+6tTctZIS5vrFFMGzt5tRnKe6q
HbEMnVO1VDzI4N59pGM5BUPkHrUx0U/mKsZD0X1EqJNgQ/zfrMiSfSumT8J57wAf
wh8fgQ2aRUxgRte93Gjzbo2c3kbRf5dL4NUX/Zdzdfn4tmAHk9DT/Xiq2FA9kOEg
mx0ALsJVauzF+HlkX3s0uplHNNCc0z4EM9gszOsBhz2Ph5qt5V68PAEJvaR138j9
Gco2A3BLjcZH9b28gQEdV9jYL4aRT3wHULSFpYFcAQAlwY1ry0yCQ1zBTb/LTXRE
QXtRbYVBKrNEAumzuY1//CEjGe4ihTa3via71btISLDdIXaKDcjcQmrwo7Jf1BaI
juOeqzNS6f7DuQ6LqHNCPsezEnQzs7AGlxVaFZ/lUyi2XCvrgZEj5iojCLmD1LDk
Pkrrk2b3BpTIgqj4WkIkZZr2ZGK6d5I2Gb+igGhAJ8vkz109H+Lfx2Y3Y3gjY2at
5bRTLP3Mpx+H5FEm9c/PeoPaEAbazNBodIm2lIGJ8Az4DIWcKhvn+pCeIIbnf/Go
UbvYV8WcQHBcwbdePqOOG5d7VT85+5+fyiSjx778rTltBhvntu5GANeoQf/LIuG2
uKBjJ/q2eNd7mkdXF5xFkYASGrb30LZxUHBwDcLketYycVIyGSeYUW8O5eD2h5rE
cgxd39Q3NPIGTpW+NPOBTC6BesKyqPdHX5UBeibOyGq0KhWLQnhgERrlOwF7yVoh
q9MEQTO3EqRfD76qiLut7JI9PmNnXicyaOKdEqEio3Ol6wqJmlco6kXNkyd7wMaT
ejtfSJTXmBmTlDmG1YZ2MGluqRPSk9Hg1U1mgxysYaHH1ooFDppxt4jcgAQR5G5Q
9ODECh+1WzNk3h2kO73MHr8U99ZWFmbQJJSnF/NjuAOQYNa55nbVqzCdgc8jfzoM
Cg6fG81AxvjXdfr9lTF+sEuBaYUtFuLVr5rQg44/GKbTb34Y+bo4vmafaeqFGUWe
FrR0NXBZVxkMCT/6Yo/y/9j38Hu6yx4A2QctdBbfV5KlG5yH/L/7L50qB6Dknriy
djfV8xfeh3mvVrwOoBQvWeeY4aidgkcvPht2Th1BgapDdxyXwLXaJ2HGn9fkRRWX
QnPzwWAc1pDP1qp1PuJwkqAo1GFnrzNTuTozlJGViyCyvdHaAYQj3ns/pi2EpxVK
P/oRvS4zxqeTPGudNufmDWoIeF8p9V5nYXryscqNTbe96s1aATR84GMj/DiutxOz
dSvfIDPK8rm0J4q+a1PmCMau3X/yi2COrwdMGhDOWFF3KgHitHN2JZzgXbgG+aMm
vvNnCgXRzgMk5Zf+gMcvNQW2ETnnJLP/OypmFRPgr78E/BuYTSMtqbfscZoC9TxM
4lZBGvK/t9e3zyTVUIeuU1zt/2vUIWzopx90ZtSKZ7K9apliD31OtjfMvX6Ntl1e
qp0/z+7wyPxDfQRRc4IcOg47AI4tcE8oDkynkn9OIitZpv5+iNhdmp1YpWXV7NNo
RmgvPYk0eO66vR0jJM/1Cew2dFKYcXuQmx2klrdmTYgSn/iiuyB6xonqIvLeAs+a
Nveqk/A4qopwjZlRJ91EevDjyfhNeS9Pl2/eNPODlBfFVqkjsZBaZsVhAsoJsVho
ni/MYNHSguzCbCJaqNdMCjSrhM7OiaN/TAk7pBRdEDuf0xhUqVCB+fgY9jVj9vj2
aRAeiHtAHEPx/OCTRJTjyxPqFu4rtxv97Q5dwC1V6NScEEfr0K7SqTw7nve2TAZ7
xpmSRxgqJtQfT5ZHgZcZAV9smEz/pfa6z9HFLQz1zJTL2bIOnLNz8pKqdYXyII3m
CHdREmWI2t7qvl0ujoGxREwiwt8mR2ZEOVbx9Lr+VMrN4o6cQ6dCEQT6cS/xUOKx
UOTS2jPEiSPUV7fiTaSOujd7lRAu/W+l7kLv8/OESeXM5hnEEVn4wvyemwQeGZbB
j2waAMxCd4DOzcT6tQ0y7rKMhlmEHmcJXx0utTtcVSWO94BBXS78SZ0XBbVxhruP
G6Tzi730WecEDHEofOd7jAQzNxqD2TglA1mRJmeKVngqXVNHT8lqb+7sN7OdKU3e
5RJ8WRx3/nK+a0aou87qsjuu6hYxgI3cVYaRGoZ9tURP/pu2AQeKg6Qoo0QWSDBk
WpLC5Xf0By3uKVBKpj2rISlA0LG+sDYWBg5MERMwoknYMCfsAq6RABhUlSSuQHZL
8dmErsdHpfEmcFm+94PhNAbx3+6UB7GRS2c8qpX6iiUuoT3x+apX+Pq0CqFDE18D
9bV7uQGjXfGoD+lOAzSDCm2WwmLphUEjMFtQyF9K4fhJRy3Y7h08+8677UfhHTf+
AxkC+DkeRNNGg6Tdk/1SVbLFuQs16gAm2cpzrAdCAM0Doj5jfIYM6n1R5Um0GkXh
ofaM/yjabfsW7Ip0SBdn5upUIjnVHh+FOuLrYslIdvT66OPdHLSYAB9cxziRLuQS
62+48LHcWVYzVEP1/eF/anQ0+0O/nKqlHUSBU87zJx6sBS9Q5avTz2Ep58p+HsZz
FJV0WAJ5JZ70xg5dn+rZz2zwt6IRP6CYOKoeoEAdfhpUpPTvpKN4xdbFOq1vyw/n
er7kcrzb4Yi24RQMV1p+POBk0XX/5x5/CStCpOfHqTj1ykt/+Bv//OFu+zqud6Dn
+iY3iJwvpA22yUmdUTi3iWAe+t3hnCdeGhTScSECgOgcaHs6TrLAza3iiEN/rASa
uj7KPnIYCGuisWM5JuoYsVyjDuOzvHOoV0HNs6giR27DeMuvXPZ6iJSy8Qxghed9
4qUBapXAJ91zhiJbmPbQPjdqUkuU/COOAfGNh5i1su7AxyI74f/MAlS2+ON5uzNB
cql8IDDvHa22HTGVEOp6SbWlvbconhtlcOXbhiHYlR20nhLcNFXJg+Fjq0WzdV1C
tF8qjL+bPhEMgOhsyKh9ASLifumrBaTC8QEADMJiBp7vr1lk/3W9xr55nwSiltAE
N+48k3IktlCCY9sQOSYkP8+OQlAYrTMzbOZKCPBHBDuI5r94YSU1wop2LJxK6b+i
OAD2FWk2b/Hiud9OXDex8NRbCC9jacH6//AUGM2exiau+kVF/hkQV9mDNBZVZ3cW
luWqkX//Cm95JVBMKfnp9144RV2TBXIUtOGbgTkQz0C8bKq/CbO0GLP0zynMQYnF
kpm3hJJws84vWkB3/Xz167F12SgKQiN71cvKbXqQKfV9WiwmHkVWWeU3kk6Dm3pq
w19zO07+eaDVj+7o5GxC5DiniFFkbh5zYxu94nqAxeudjE7e9+4yUUnb6x9tVMr7
4MNUPCXHWKe4eo7T7BOklIHuObrK2A8YZaB9idEBNebCpL7mJ265LuuA3kP7Sn/i
JuPAuMiej8EDMxw0IDec2KSIsSLcby55705Ta4SrOlw1go1Lwk1fy49T7D8Tg7hj
dJO803DcFRxCYiqniO8+bjD9kAMZnZFnUti3QVS0N4gfWXtQhVy4MciblXulZ5BB
Lwvphr1Y8hjEliwVYRQ9HZzub5OC0s+1HgVC7yICGoHPmJ0/khu91eN5dk7g6cgX
b5RDXo9a7/liAd1vtUkS5jIF+W8NLm+4RWDVl4LLr2ibrSAOLhyZY37WobSoHbek
bfn7PUCBkhBiWjOlNbD1LGfHkL9aA4lWPSgrMcWeBL4MKpngpGWi7PZ33H9roSsX
HDohvOdZYOd9k1aI26RH+5Ob13KahsxwAjAhMklLhpLKkwvYe+Qa92JTzGAuoMAH
pj43sXzTXiTqgjI+Y8BaEyhB5EbrSrAe8OoqrD96gQ9VpzvmXLo2WThvidCAb+wM
xxJxDl2KbeEF2CkWgKIL6/NEyOBtZFJbhJVZSqukLCgyOZYtXJG0tsjYcfH6B9Ry
87DlvHkkCX6XpbeOiKIsCmpO7TNvVo1hTroytfbrlAvwywWYGz+h0Iwz4bZC167N
/AU30lzf4ERXwZ2c8CTVUwsWnjaEn7uoYXb82A8on1mKH7Fo4CWT9MOt8GY7YbMB
F7ene8e7kBImP7ZWYgLLscgWfThwuqCrRvO9QL5D6kbWhYRisHXA1ko6hfRpUj18
Z1s5GwuO7AIRbjiRc0mAKfnTG+8D22WRBPsUSD3K+QyhGU1DTge7SfMuPWu8J8R0
E22TG6VLuQd2cz8/d6M++wJMP7H2ieGpGlyrxCiAnNT9AuxZdUO7bccddriLqAps
+Y3rkW764MilhCXuRnhMCQ4xhZGFtCSay5Le7Dk5UNEaSr2fwiEW5+0xl/tptTQ8
NNq3HG9S2HHlMFHt28OuLLyZln0k9+3Ldc8X4hxghxFEZXMv9Exr7rynGiXL79Mk
uarOfHzEinayQdXjQc1u2D3zW0TL4cy8nQ/QWwN3V/3mANNTyLq1PufMvRnjyTeb
SbIP20KrOHxBBQV82Kp1gub7LxJljWyKY9XoexnOYJCt9am+ZTXXWTIoMIBmv4mh
CeAcdL7uavvuVnJ642c0GsIJB9YmJj+qwAwszK+NLhLL3/7LLMk/bWzOQQw3NiAS
vMJksM11z2DwixhRX9oUKWM26wMCoq3OyDl5Q6l8MT6Hbz1R8iU7ZVdJ3YFnbDgd
4UBLVSiCbeBAWTCLcRFi9mxSiNIPwfk6ysevDZvDK2xMEDPIBk0KISpOckpUEvV+
UyCpTgvVGkyyY3Pb4pQ5Rdv8bAcYyP7YaD0WR40fOgMtB3dDuvn7pNL1PFVoy3pU
e8+V3y2LSOKsGvX3hl4s02YYhkPEN3mhAHcisJRN8u++ko4tvOadvK5W9HFqa2Fw
K3t74D0lGgZF5y9NamMu7KseHJvL97BUSnoptnGQxrBZQr3ACDpFn5ySjh7pzO7n
IU7CAZtp/4Ze5J+4Iu4Qbfv0cdqTi1AhwM1Jc0lgYNajUgBTfn8dBu2v2PlBucr1
MYF6tehUzEz/0kC76TifEgyBh9omgiC0eYs9AiMXw29QTLSN9IsGElp/YGCtCVcv
aK6aIT6Iq0M3CYegUrSait7e8BSqjyc6Vavnwnw8wVpQsGD/wBMhlR20gjFiExdQ
zh0VluVEvHvIoSUzpFA83x13w655SjIGL/wjFzrV/8NJoYunjI0mfVzw3I1hBAHT
75oIQf+iWDCzYt38kl7falmq0Uk9y206u5uWxlxev9WmveIRxhqRHwF4THj6rZKc
u9yeWO3oLU95UWolJyl37m9M0RE4wT9Cwbnwq0e3viM9r1sPdJ/nGsT3Ue4LgSvL
JDehd5vcmfYFqJ7vjCHGgyCIgxTBW/nkxmI7lxtk/EUMLVGfdd4+lNAyMi+NrAWe
z5UrTEqd6afaMIYVvB+Zd6jhyB1etjiaq7YIgSK7DeFZfET1J2tlvwRm4tRcpjsv
UnOs45EA9RKRgaP0HTLYm6JP7VpbXMGAGIn/KEYRCvdTsED0EvtCWHYDmkRWudZS
degH6T39e2PISSM5sA0hREPV0dttJnU86Y+hOgWgbFT92QkngJScjDYaxh8kYS4+
m952iNKz7XlgHBAWFncNMcMCXbFu6Adhp75T10qaCUwKJivZBPZxBUhG1X6PmFqR
ZvTBMRBz4H5GLRDMBN1gt1vG+rduu5zGHRevaHTsQ8ITs5QUroZNwS/57W4m4HG4
P+1DBcPfoZrXUe50P4jiIOrRwxZrjNFUpxxxcxKQz+EcMGlxfrNRBhYqqdyzY/wm
a0gx3EwzQrOma0Xa9koGWb45i5o2v+bscx4WjPjGkTnXXy7Fyw7ERCGP/lCkPvuy
32DWHOxgx2wBsbJdLzQe3q6FZcFsIbTkvasB2Yk6HXTwhUfPZumayxWvmh3sOJQi
eG3WIjfWsNQAWUa3XpjEUk07+Aohj1xIKx2Tit8jPMUIQu5xrqt/HMjVU3p/r+QA
yCCsLJ+hrg74OQZqSbGPnW7yoM5UDYLAIQ6/YSG3oqlq2eV1hlQ6ZXWAgEAWhfTx
Kqo6/O+Xi43yl6jesiZ6++yYRP3wKANE4d4x7ZQLM8wpa8hmuKhPSAAgnOB31usN
xBwG4Rapl7xqdB+9F5/u6QisxPZ+jPn5DxBQn7EDF5BxgQmuyETb/EPdHu7smmXV
Lp/iBaKsST+NsR12a6/uWzAKzdUsWtT/KHT88MQFAuzCiMMVm89KY5C9BwW2hCJG
Ct/4gVQnsqmNrlfGzlE0goceuZX9Ibucke6iI1k92VmLZGkqdYjLGU3ObEShTQvJ
jKSvdRXFeT9e5NH7Y3gCHDXYmwTKlekmQFmAIaZgEEqyD9FbFlFdJTM64eh1mGX8
QTEfb4WYPd2IonWlM6PC4jMfKhNwtPZaKEh1Rw9f70iNpVLtszl81wLJbaagCXxK
Prv3awu5KNTJ+GEmcUNxvn4Ld45VRnxETSukMt6IgBfkmTKxJHB1SznuJYEfbLi+
2/jAloD/RckGMczkmqwCedofFkx5TyUWZfV+rfQaveSP/U0K+VBestbhnemqCxNe
583QrZrglBG1mdLyigRksbPSNOAP1yTrkHNPlM+C/hwBxgHZorGLNNjuxguLE40O
Jh5addHFtsmTmXAj7Pa0VSsx19/jmmLsKkbHkbWyrrwOLedLKACIFkub2sRCRyga
hLG95Y1RGeYM3MHfm1JwtS4NU59cDkXroT1273DLa9QVRTyvJ+GPImp1HUJSG1HN
vAO9Grc2Zy3c4bcPhePdk40ybK3J6j8RCXoNyDo9ILdKt9eE6YWf5bYUshRiDVH1
j+IBSSBdiioBJlTmgekDXqTSeBkPCBAFsofzZfLie+1kA2H+dauXzTUv1Hk1CTKr
POJ0TLKw/lFm55l/Znh1n46q/Fl2ijYtac9mGuk04IeoCnwGx9cjZQUK4baH9XB1
Jwop1NIjqNdsCroBsIpCAEDLAFRNR50fyzv1CV7FbgLsVtMZbITdtjuGeovAva6Q
2N/aoOnpsRtKYX08fFP+qfuOIC/zaE7tA+YYp1gbWkwA/nIHef6kCDorpuxgVAKz
nyocPNdT4bmxsfXh4xDGWney/em0XsGXbmfFRXaMd7DwT+tAFwYyvNPmmgQmNahN
ASgCv2MnWxPIlKIthXWF96u2F/V67Q4u8lnmo6MA9QqMnMSshNc9gwBJW9areAMI
3P5pdWFg1+iMEXQ2TSzwbDZ/M172N3BFCSKwzEa56QNCiIiubERGdO6Pwfm5PU0a
LTzG/mWbtF+K6ds7Ryz4fddv5Hco2kjvy9LozqnsXtMp6BydPfnES2zlG7vDnOZD
RQxzjxDsM+8/RNmZTROyRYtKx93eG9rVVytC2UNVI1+Ahm3HBedKUQxss6hymK2X
OiTTN0zr4q5Q0Rco2Et0vT+blW7REf9/SjO9VJIOCgMZjg1KzLVkG58J40XA8Kwy
Xy9FvGxks1KhoJuIhvTiHLurROMsW0P5xcIkulXJs24R7cJKckhHJZXoLmD/ACsq
UKDkvBAju4iPwlXHS7KZb8r1tCp8feHpIYrZcRzCfCDo9UIbRCLcZ+hXXKjSiuFZ
zzuxsFLPWQII2LrTrom+cETpeHXdoxAgaoDZvVixxcCXLI7w3wQ9L46S3SsH6LVN
jD50S5JCszcxvxwU4/aH0WPi9EgWVvXSWp1QM/JlYNGHdO0+UDXQJzIouWT4+bCR
lobM5yZwpM1cImfSoFUsUVvOBGzexckY12l5jCukgUkv5PRySrFR1jic0KlBDBar
BsHZEFJ+V5d/AEuFfwgguidN395Oyty6qTcwPt5M9bMG/ceBbw6AHB+SEQSwtlJK
1UwU0YdkuOz3VcH5DIirtm2qs7qlZ5Hd3XpE6htpE7KPL9ATkkRVQ9rkjncb2BiI
DeGvXvSRhuXAYag30PjACsZx0mNgkXZMtXJ7CMUFNieQclJmYQ1BxaM7n92XJkt6
QoH5HqYVbU69Hyd8Ah67BcuqtKYVxb94vdxl0aq0N1DraYZAa1pGvx02pPcTARXG
vNuAHhVTzA+boxzfkdXLCPqy3q8zUx+LXfb08iI/6EgUns7rutuH3Mmyk8YHqqz7
yUAXbTiz/b7U+uvE0alBbIWLCp4cMxv8Q1nlkWdZ03Fdvq9BsHz9eM7CRFlmvVvq
FMtfoD+YTyxbveRwUXGaISC/FSenH060LRP58Xhd+m3HDKY4PW0YwxGIsoRcQ0bh
/zrnHrIUfkJfYyqzY/zfGRiZg1RvOvF+IEp8ob5xLwWoX/IDDvF7ZO23d1yJyeME
fy+ixdmfqFJugIDRIUv0dp45thBgUYlp+aLkqZGSbPuB6EK4ON8PCL98X6q/EETv
ANqf8YCGsxxg/iWL2O8TrdJR/veFCNHGp4yDuadH9Y65aFbX8iXLbBr8flcHXW0n
oY2Hm5O2vBPPR3JsIstZLWaGK4xupcMP8Zw7JDn/TwNXjVRjKdyJKFeyW7v+8ehT
Fi/ABULtYX0UM2mn8Qyvoch3Xc9udSlPDLumsX0oOoTKmmtprBCbYaVEUtl22E06
OM2WIq3PGzVZdKDHQe9THo7sqEPJjpnNOZ6CHm8xNwD+/CDXtorHcPReZAOUY0Fc
AFFon6ld7JcFrqejCMokqHQGbI1vT9nEw8adbEt06DVL6i+sa6VfDwgfmF2ANj6x
zvujiVl/4TbRii/z/7lE6dpbyInbgqyKIGPpIsknfQLVcWURPiU9IHUK2MwOHUmy
pR3FThbbi6+C60gb0sgh8jGiFtTGnjAJ79+/32A0JTKy1AtzTp1wsI+tbu54zohu
DfeDWe7ZUnT2mKw4OddrO5JRGH7fslFnFMAKg3wIPA+WYKXJcP1XsAKJe+5oMqrp
v7I2YMrI/vYt/Md6VwG+5sxLZv725+8pGCvGjCeJ28fDnJ2Yb0LaKGDg9uoQoCnc
Ol8Oz/YzYewjban2xD9KqA77WR90VtuDFYOXPxQJzcg6/tW+VRGC1MCrEmKdGcqj
t2Q+WJczKriO7N/EkvzeiAPZ1yMzvzfsXgVv8DR5vxQ73TlJGfKrbNy/vFk1Yca3
HaNcysS0bANg0wTvt+B8IHHvscM5xl6fLN4gi7TVi7u1USFRmUVSykn+WARFteNk
2uGCPd+uwVFhq+0einN3V788aH3ENve2NMvGt29XS2gX2tiXC0IGwVBfHRzZhize
awg/vJw3ETXtvY2HEkqkoLiIwd3a3C9uQgUPFIqYDEtKfOGZphm3WPXm8pKsoKU7
tGRuxUqz8f4pk+GyE0eV1qmAnDaf3HZBO7i12vZBe7WIYB5Lj3VyHSIezb4rG2Mv
GRWhH38lXdHq2R1U2WoRaOK4HuJdSttG/r7oNTshdhfOahAJ2PkdZwVoQIz7E5LJ
LM4jQJ1XwcdXxPxUoSLqdVyoQULGleWLQih6cBQGjthrDPxPoasjDO+Eg8mRBuH7
9+4A2hLxKsMdIHQRyO07kpNRWs8QegG0CvO2YfBV4oWiHsMVXN8vyi4Zqs3fhUUW
9bvNdPUMwzSj0ipXZGAoZAtbTfHf4nj/yvQZ2f7qpFuia+nTcKyJ931n4nJ5RHRS
akuw/JOE4eDz2zb4JOliP/GTqFYgheJFfcEzn7fbgCjuJ/ngOGci15FKwg4kB6Bb
R9MqksFbsa7xMRk3/JvOd+teiz2qUT9/NBYd6z5rhWwhGmpWhjKZaSE5pvfzoDZ+
CfBhurtUM4E5MDgVxZeN7srshtGS+p52iFJlTXmbVbxtiUAm3hA6x/QeHsO3HG3d
8vDMmkL2hpc57nOd8e9xZh4FynsCPlJ6DDMQ2F6mdn8KAZvevPFZynFFyhFIsezo
7xu/CaBnryg8sDrR9sNqrQZ6FbC7J34SMvs0+fMvXFegnqQ5zHaf2x21X9D6+Smj
EAnw5IzZrpLPmMiKbplgpIEKfw3SzKZEJ51jjZb3TguCvNjt6cc/21Cz5OUldM8R
bxNKyXH/RpTx+Qi5kJi27ahnBUWcBmu7uFIi3RmeydssTe2l5oPTxA3ixq1lRZGq
vc0Sc8lLEwzQXhIfmL4AGtULge3M03x4STAY+FaDSEqDEvv8EVMALh1xIoqbhe/5
M53CkwhN3pGXzHIdqbyCHxcOPtceNE4wc1rWh25l0WgLNuXqPqHfVgJg+OWz8nIR
6bhkQrfElsk0djwXxzUUIrWiXujYpktJlPiiy/CAkwYokL0eDP6zI8AlSnnAytt+
7XaN+0NMILbYgKIDrvEJt5GSvsTsDQX8qtJAUYdUaixtjawrswj7O3n0eR9XWs9+
SVBiEW+Lrqq5/vpwWwvdd1+w46ZRyb1WrIdXHmXapapOaZ+WozQHZov4RPTeEnfx
9NcEihYdGOpkDm4qe8Yi/9fOSAN2SyUGvywXV2EgC9WqsGf4MQYDuM5eGHTioi3T
lHeXHDRkpM4/d7TsE0VmC88Mo9wh4f7SkoIx4Zia4p4Xtk1sPnP6RO+I+Z5VsTBy
ZSHX33rq6s3UusWkMxw8izj8QayzN6B/ib7mgXsAmCpa4AFpVcWyRn72Cz3ipaGt
3tgocxrgPhnHHvjagjHlvexExczakmbGPJ+zopNeeNkUhqUMjTyswiqNxp+ozRi1
aan4iP+XvdWJs4HHsVwsb0wq8KRuEktujfnJDC/RL/oSnQZGkCpGIfgCzDxr9F2s
xv4dk9ykUC52wAe4C3D/U03TDFRKIrsVeHoI4zoyTlRqUs+wKlKtustwm92eEmz5
MARTJtyg7+U+S10rdORBmnnF4HBBqcU6/NrrivAdNXunXmpUEMPQLnPb7SSHtuAL
maGN9H3LEy3gI7323i6flrw3UWa05mw0i+1YMimbbp/lOVfb4hNbzWHh2j282VfP
xmRk5ljqAMXapw5m66LJBCO7BQTRvBeTM2CCfGV2pw/WAVyKeoMOqrXgZeXGxM3e
VFnJtweesF9Ol8JYNQ2gneoirx0jMlSBiLZrLnf/a2sb/oKja9ZiQq4Fa3T3Y57Q
fAWJFwq3k0JuTytJfaBVrmyoDsQ8X1LY1o6I+a9ABPnEuoCeWOKPLYIphD9n3ERK
BGpvdgO4qxXLioFQlt+5gQwn960Rgi39M7eHAF5Plo+CZR5ybDadQXxv1aqUHzvE
Uy3F1EhFCgFukcwBh13wF+BPgDE77pj8xlC3EEUzZWzdZXGzRJWYe5BP8XJJkPH+
OZ0mIcby/Wt5LfB9KEJE2isA1+9LT9dvcM2SVSQEEoiyync3HMYVWOZ5bnfywaTT
QWxyeYjhInXF4SoV1lkiZgHrYR1gaqm5Wi+HrgQYHLVIZFGdh9nDuJBweCD4lEjP
oic+uvkupixbCcrbhuNdFB2vOPXSlnlInuIESNESfEUtLlibfvxTxopZClpBD8yo
9t8Y1HcQ7e3c4t+Mgr5exNTKszI0GqN5S/w36YcXYMvweej4pqdrI5BqbQcd81Oh
1XaFWYL4jHQt2I4VtBGNhhu6KLRk9mWOyhxzDxI/QOqfoR0oK6alCJrua5ioXYCy
lM9jUAITXzLb8Z2Flcby5sLDx/PhoBZsqGV3Jk360caOpMkuppohYo00j1JDWXQq
uHpxCoQRy9uv2ApbjWAUQqeBkcsR9fbgECDUByFaAUErviWNSfuHsx6mGfE19fWw
GaWEG6kL2k55AMxPvhRmtY8ki2D3nJhoKGJNp52dE4cF9MfuDATVA/S2IvFpywWg
cyrgym1OVsnv4MmGl4dbc8eAn013zUp14+hmnuVmrP9bRLhY8nJforpYHFLcBYVw
cA1NrYVooZTc8kcylOHVa3YffABNRbvCqXa671ufN2pNqehRj/LQLA4x2zlKCoSc
p77/0elBdo/YHYyRqIFNmzNfHUuJ06pp+aTh7dhWYAoDyLnI65fLMlA6g+oO31Yo
3rRaHNjBsd7SSCK2s0DcmeF3PerMvuGpugTZg1b4aDmLvLHzswrehTVSICJNtLgA
PaOUfyVyxhd/2YZ61vvjMfglaIJSIU7MXlREFetGhyMSC/dI4EEXnUcwH2AYcexi
mxk+8CEHp2y4BmaWH0iOop8BgodjukrNg1E5qYheMQ19zXKGl7oJxU6ja/xx6rp/
xcg9xdlnSqbLKZ+xZiPhGOpH/DdLKoFfb/5eXB/+Q9zemZZR6Ck/unIf5ozsnZDk
vCXcwdX2fq9GK4Ia/czSI6Dta6RZSgs1SOT2M1pR41J4q0h+30QSjRTbxkQ5TUp7
dTlgwBa70KJevWJtklEN+M5T+5dnc0Na4ZP15Bw5JL2s0BArzslsFwzwfOq2VPAB
924tFqCeWsk3TvX/cERHMty9AhI1+9UNYQO2J+wMk7wmfXufSE+y/ltZ8KIJVYx1
2Rvj9P66qddaa+nHKn94ussNUzqab23Cqdbmjoq4PDpBRwvnD0vtNm/Gw8yDlKGZ
GlGTB+kngp36vf5zYX9S1qvG7j39bxy8bLjIiEEQRjvq1wbgkphWd0PRCSfh9l5Z
0yYH1UVMyyuSkz+53gS2WNa+7M0xvKEh5VdaUOPHCen/XZOKGsTfWxoEKCnEVRuD
2E9qwIJX5o1VBUmN0tZrbttnWUX3sIxNIm4wqHZuZz7+v6KvE6YWonuW1w/kPmU6
ITScIEE2cQg/pxSInk7HCiY7y4f7F3mn4pkBLgTYz+aFIb+IHjZn5omSboLKFygp
ODuoQiVbhgjnpdk3skx5n8fYvzVbbdUqNzIgBi3GnR2goKsl9c/cPiOCBhivyCt5
O1/rTXOIZhMTPEOa7xNkjqcIVOU7d08zdqshfVIp4cAVpJINN6+AjXq5892OZWLm
uNHs9+SmCeu3vkKVmrDyYaS+5SiFcGm2OxX+UmMq8YW9fWgPK+CSK94Y39Tc/s7p
TlOmbtx15ngRN5Rxz5xfS6nZ4Plfog485cD9VYvf9OE6m/ajaZ7/f6iMgS2gvIbG
qfixaz9Ton/hU7mt/U+J3kjpQhkqTgh6NX4U/JJZ9pZdfLLxG/EqgBDUYLZi4LT+
IaQZhpqMtzXJBi+UyX2x6TSSx56m1uB2ASws3V8NSSRcVygwB2mkDVbalgB2iTh1
zbSpGN1PtK6CzdZ+uYKNDUEe0ZvXUbNHPbobxooRrruEeFn+aR/9Wk6CNDXhG8fp
Ol0aR6uO0+i1UFjjgdbnVyq1c2ORHTt50AVJyYSXxNdeSbpgv03MHAprIesgeFhW
OaruzRWDgnmByzzfEp+n8uDJrBsqzOwdbSB1XAySMrh+OHFos2Jafo0el3eUd8QM
zmTuo/+vraiKc5Nb5+ttIQH9cnxdpUn/HThWq9L7C0lXXEyPGlfBxUScZn6/hguP
UXDflSfQcg8IEqjpR+AmqPY3phzoT/FHeDxjWYj6+aGegp8HB3/0SYNnNcAIdPmW
Wbiq/GQrGN7P5q/HXxVFQ0X3LU0sspJeaoLwVborA31Yp4L5XLZvorWwRsUy/sfo
CmYLfF5JnK7AnyzNyF3wHkv0KOFU4pIf1EsonHzGI2OI9vsMlWV8BMn/vNtovtYk
cYIVzFUW6woKgjDq/ZS3r/UFU3PsZJHaS/pBZnyKnzQIhU5gWuqOFDtHOp25TZt3
+QBNeJYdbezkhiyoLbx7yCbQsjTAMhKHj6f20kO0z0vSSBAO147Yua1kOdX1r2HY
J5V+Lp7pDi1Mer2orUXYqT8DMOYMnshdJLo8wl6xmktZAENQielzbqnymMM6K1CE
qJPdFSmOGPgzjGKckBzRr48OvuW/A/4yP/WqEwOztHG52VydQRsjNDY82/3LgUhQ
8DNQyJZcaNab6f7W4+/2BwX5uFlmRL89OrNlmAK71C6EKriJJ0w1fMe3CY5hSZQ1
yKA5Tze6EXlA9TUBgGU3sj2OztwztXZHtHYuU8F5Y4a3pZyQ9FH2ILl/r8BxdErK
Jr9UNLtHPHx824qgedBu6zt2AlAwbHvIBaC/dhxrHOUnBVMJwwnAI1fJi1HLd660
l0iGWN1FnZFOGEAKQfTcBVDeOFCJRP7UMb2jcAeb34tMYRT2t9wsyKJV2Q3/XyUj
3vgiJDf7VWDjHguO6BJunWbYmioRj0hmlsPLZXjo+DxWGoFQzNyC2D1Z6J30GN7a
JoH+diE+zVUPKWxIslPXc3cdo+MQLE9Ok5xHjEDQjFHQKQWH3tTNtKb6baB1cdpX
qyvrmL4TWusl6JK/Gz7OALqsO8wvapYP276F9oYqF/uA/pa59x6wfpMkRzIrqDx+
jV8TGBue3WpqKMu58NTZlFuhfRevcYAhTLkCvhK6wNaj2/7ldlVtirrhuNXEbJoI
hvNJRDSq87EVPUqOKgFD/IV4MN8X42RvAzsjkIZZ0HRbR7kGQ2GwfwZeY7EfsJ8q
F3qBs6LMmWVshKGz/KtTCCYoeXJscKDbhEXMwIS7vvLoGARGY7tulDYswghxzVuu
qrQLyYOUoIR6ZRhK85/bUANVA8B4Et17Hqg2TbR2sIHI0h/vKG4vlqCTbhQlpA+y
SqCb344qtitUlkLSYUmyUoYQpnJkf2/ru0V64y4kG9BVta+ZFK73BiCDBkJbX27T
HmL95p11GULnB/vb+T2f+ZIc8yJlHw0BHqq8pEML2N8hfMmBYzv2OftlCBhzXRU6
P69ONRUAf+y7482+UBsYPJ2waf25ANj8qLqFtv8QTE89ibAK0AozwdzfsLAvdgrJ
fNnx/TuidMY0I9a2ZcC2y4aqNpEAOKIgf5gEemOHVEDcSHI77ABXMdpIOd5zZLSX
BW24CIEhh7+5IgV9igL4mHHJB+iXbQtKXU2PBtE1xJLASdwammCtum3Wdmpd5Rxo
OqCEPYArbpLQ4FZHV60UE99b/FoPGyEvL5gB33mEdAR7zUJ5qtIrEG80GHs70hCl
Z7QycooQYbJAkK1w/P33vMajqtscPwCMrYq58SDvbRynfuuYCT4E9cojcmH9nB0p
7z9A74twggevBsxy1L8ABtulbc70BSeqfmEdMq6SPhB9ojdh4q1vxXG/ehMt6N+X
KV2zVdsI8slnw7cgMS7HyF+WESV6wAFSKerO9iZPlgVL2TXO4Y9XMObEyCFtTaEV
4n4uUF18hzg6F1JZ7i7txFiy7DfdXYlMXhxlZ99kC6w9GzyctHxaclZZfIrecxD/
3UZYPf33zrVEM85M4ET70I2sfXV2A7mexKjuwlz4ki9BCo9a7VFxI0HbuApKLyWR
T6h5WHUCtTzN+EYwQKl4nI+pqiW6RBotB0qlSR/wYYfNyjN2uPElzz/+Xeh40YPx
vR+iihjwqWEbHfFN4JtsbseqBXPcNpD2r6Fxd7wNJ+6dqW7EisFmG7vrhYJd1qQr
89fIGlp8xiCdUgmGj1EzqLP/Zxpl9h3MDza0gKxTWd2nf0ebNfxsWE1rUEfBve9+
Sk293xDMN/ZGdNhvvYh12d9pr//Pmw4ifbXhRvBH88nahgtr1AjpPfC4X8vVorXe
QTqvoEpxcics5JSA/EbG0kD4C//WvPh0hCS8PqXp64vVM7I1XhQaDDemMSJRD7z0
beyPMdYTDarglMGa3Wknr/TbUlXMIfRZ8fxpcSfiscYhc3Qqx4NggItKMb4PjiEq
wWMaLJSrIefROU+W+pRbX6lIEi6bJfeLjjA2K3wWQsEkZzUxSAtYgi/Fv+/kC4xG
VPBrYeiitdxNkGh+MZtMkvnQnVoDy1Ge0R+OUFeD80NI3F3hhR3HFI/v1ta4VdOI
nkfljYkMqIsbc4YYSiXJ5PKrZGSMH/dXqncwY4YvAqd3CSYJa6Mu82YmMhFAaCvs
GT4uafvX9bEGNrIEw94+eBhirDD4nIKp6B0gctrTbKhqdfT6LAEz2H7r9olMJawx
HfaqKhZDOdNEdg3kGHSLK7UZi+RFqIdMwvJh/kkjmckDrLhI6S3UL7MUQ8BHoZrM
/a2lDxEo3xMOHNkv3qO021znHl3/uvc+44D8gGqOIXPOJkpDWfVNDPA0ZuY9iSVx
fVz9KQWU1BeIfC7IuY0zWS4izdc0KvJ3bd27K061mp/b3uCe9VPB3utRqzQY847G
WQOOf1YLA4HX1lmfHOPwGXQQGZXIahfPYmjezrlmgnvQkKUQNvFzbmwZJBB52Qct
6l0r99GsNGOlthAe8PL8Qb69zW94f4L9BV9gdaNJQa1oh+wUmQ+NAXdrXiaR/UUe
4k40chZs8zIZbL6jdzv0shtafazBZsGcKKnhX6EqI1NGW7Oagpg/FI6B5qiclxKU
DxeXNlE4ia8MhGl6DSINdJ3GhBEmZtehq86Jrg6wf42HiPKPF1Ocjf/wnov0FnLZ
5TMkpTKbfBUErqvyRa2Y5seumK0yxG3TCCjnNHkqdaOklEw6CiJNj56VYqqpIC7n
6fq/0Seog8XsfIqJ66bxox69to6D9kqNiDt2svlP2bKQKIFdIJh6ObBJKf+QJUah
TSW8oZWFiupQODTI2cxf1pC6aHEpN8rzML5KVHr6MbHhMDtjsqMCrfOMWOMAhJSB
xj9T3YjT6hRyTMOA5UUzoxGYJmDh8HSsQOsRQ6Z1zXsXhNX2R4mzlS9Zi95jpylB
MXVeDdR3FGnFXTIm4w8YNmfK4Uq30FijLKeLsHs5zY+m9+zLIDp08t/I/BMJASQ2
QEIrJkw3P7tTQigG6OfiJKnsguY+9wV83OrDbj2L4RLtbtxgDbn5yPxn7mvHhs9m
ySBlTjuz/pk8PbJ0zZJz/wS8yzvhwPsqs8cfQjEDBU8KUg0kH5dOPygkuPAWo6CS
/X2W/986tfjP03HpU45rwolfyrjo3xTxwoLNXwhjaAk1soCzr1jBWFzlNs5PLO6y
dnpE7g5Oa8jUNVZ5W5kGR4ObjH1px8xQ9cBmtK+qDf7t63Q602On8M/dMQJkmXzB
jmKJ5HlUbj4L5R80UGGVAMkKdZvIFYI/vUe1ZsCdGqtIGdmKiJvtLS6pFiOknzyl
gfJdVsMm2PI4zNRa9Url/JbOh1yS1bSABHMzpxsiVsWJPxIyuPrFzdMEakeNPWOE
s6fQzTG+x9xlzqKmay5xcICTeTTSy4PQCnUstlzuGCmpJVfbqZgCZgeD+Wb/E1LX
lg3RpPSu7X9+mQzk/eL5lnACgDMfsJHVmg0mOmqgUJpW0ymz4qGsao6aKIJ6i1ze
PoPdFecHPY6mfM0C7UJbuH+OSov0Hdw35KyOCajfChLW5hK3yA2Hd7+NIeXuwfk6
rmI+xPj1VvbQRWBppA9GOPB2TlB3U8FB/tHsKhF7Zuv8HyamoDmvYHbD2gMzJ0KK
ENaiKML1h4LCBHtaJSLbX2SM8VlXbbOZ5PY4b+Bx6ELaByBAKzNUatb+aAFDEdEz
OSuyBtpSvPIodhe2nPA5X6Ly7yUGEuglYiR2V+xdTp984Wdc84Puk2Le7c9UqOgi
91Gx7BoPYMhJQY9/F8PEgMAFeifhHyUEg0Fpc9JAHlhHVxRc5dd/gTbekDAA3ger
kjqfMxo1C8H+ZduYVfiujt+KtjseoGvgjkM21B56sdFDkIkAU1ZCTsZIBEgPmf2h
SitDodFWrg+Js4NXhrEdB6h01fgyoKKh+tiWkaZYRUmnkRF81SnXl5DQFRko9All
LRhwvzDbLBPn1bm620OmGkH20FU2YR/RaBHsZZVk+QlL88tkC0XzQDLY4xggVH6J
d66rWvlA7L5if+9e7o0CnhvVSFzu1L5hiAJqXB7z5Pa/JjNs2cFHc7aWJUre3LgI
PLS4qxoOBiJiNMvXcH5rY6uHlOF0h3hyXoQC7oTaPFmQkT/uSLugl9+aJViKY7Fb
qXeb+zKKdvAXuaf1ASpjPZRU1p0qzUBv1rus/98Px1X4CpZeSGRa+MHsav55gBzg
RWb9eG34IFmx3u6bLn7w2UXRjr2rp3dModynJ5sL5bidlu7g3i8pF2rxnt8OUaGr
RUTzpmuc6wuRnv0wLsHPxXj2v9nWx35/85b065vQEzT+/4JaOFLK7jDidKPs4loE
o8C7wT0IONr9Z2tBOs6aydrWgCZQdVcJ77DyUy7hJIwPP3n46UAWjuNn+s9gXnrY
Pqko9UNYVsbNEFH+GHYv4eEkpsPFrCEbOLFc1mcZag7QQT+McPeleqbYDwN5kgxQ
Nw6dHAPSFYl0jEmJtVr6euOItarnVJhEYgp1J2N4W/qJI3WulPJNO7xqX0PkL08y
LOHqXEtqY0V1Cl74js26lPBq8sIQZdwBgsAdkfHNsUOY0drpVoC0jhGix24j01bc
7ZbEbcV1KVS2FKIL8E/93M8rSGEeftRc6pXbINTzmwuZuZrT2abGfgBnaIP/XJeV
i84+i3wdEADeKcDY+73ccI6dIFPxyetRxWdnpcn6WzziR5NjB7deHEEisL6qyT7V
UHbhMBpi27ftKq2WXCdPxLQxqlY/QTaXAfmG6d2dBNwyBNYFHgVvKccZGB3lzB+H
f7DofXf72WC8CtLIdUodeQstxgIgtic7qjcmyJ+Bq2uzFaJjAodH5hZqERDahlfV
zOtN7YNRZnqW8e/3j08QCWl4cxGZeT3XjoYk9oNu+P1l+MMTXLAmAc/S5ftdtQtu
OiAshFmX82YvcldpiamFQL78OssN3yjBiOJpvdCRs+57+ReM+CHrFkUKw+SohrKB
sCZvkSsBBO1b1gMTVyClpOI2VPFpkStHPuOC7BAYHYtcNX+lXDf8kUmJn7DEfbEj
hKSm+0yvNZc9zY700jnsqP3CjocdL/eigXXoVmdHLMzmbfi4/5CuRY0nA4gFywLc
5aTu8XSTTXH7ztq28fnxU8bg/UP8zl3UNbhggPqOatdxIy+kxTJEVwJqV1JZaNzr
QtzV0TtD7s3Q5/wzjwW8iqionCX2ut42RHBSRODFr03BVIq5qeNiu7hjT2ymDjY7
HRd5EkfjcjJhtEelah3TcwzpCfNaGz+HSHBt9Voo8dOW3HYG2zwnNOuGGUKVAPaC
MioQSeSqx1p6Rjg7xiJbE4EeezSaWie1vDf4AspcbxjzaAaOW/pzMRGiCn6STd19
r/IE66ShRyQr3/iuu8anOcK5aBDG1qRY1YbrABW0BAMxQ9o8PxbJxr39MphuMGN9
4CjxW4Bpe6Yep2ciyJyd071PyKJlJHybjbZyqKvQfT5JbJIQKiF24cc8cBkkVV+c
v7/5OnxnyV9l8g1lK0exZd+QzK2+q21GKUOewocSzTOGj1p8cf2a6ZwcOJdrl2no
itBEl6p8f/FFEcukx3hqc1XC+7GK+kIwB/huL2ch7mX5oZSXvJbWmIHFSzECV8lg
8C3KEa4hxU4guhd7vk36RHehUXcagsc6TRmVxm71mMZURgYJpWn0TTJyx9/Rmsab
T7N+4t9b03YYP1h24Vjay8gogNpvfNcF3Lq/rhimcb388MtfU5uZBQ5kO5MF7oE/
7dBHcskg5/8S2pSzf2HE302zp3mCJEdgG1OjmyrU9AWSkkZfA1HIdIjOaViYrwdY
wM56Jy2izJHH01JEq7yq5erYerz6xeLUuXrcra4ALs0K/ol3rXks3Ac2bsj2OGaJ
hMPbuznC9pWReL5e4IYjGWLMOeAWXkEZtrUMWA6tNeRg18fVQG/cVb7A2DNe4hxY
eBbcH6kUIoSlipSx6RIMbssrgZkd3iV4MH4ezWzmlx8IVdc4gELjnzoSa40/6nfD
rJ0HaOWyEEWszGS+QajUNh5DPEJpg7AMalKaXFYiOQ5zwR8pwaz+/cfkENvshSqk
I0xj/Q0HU4iNLvn1z0eDfHJwtHTfiiMFOeX1DLPj5qUmpQfOyE+KPrQicE3zBPkM
hGbSACW/W+lPOZwswKyg8eTTK8w1Xa5NBGQEjaEWM3QU/h/QfZFgcg7PwY1fr+PL
HEoXhFLRGIk3T50YhNv2D5O7qOW0l9hyt9l7y9F6Uj+7nMI0hQvpN8KBgXUGxGLw
N/DpqiW5pZqxxovWGk24ozjE1aBPe+Osw575bIjdtlWKK2Zn3n6hJZ3x5+CNGqwp
k+vyMUXEmbObSYde01mPoteg818gFSgpGBo0baRnI/1OZ/e/qtiPUU8S/ispPBgl
95Kgj6lA/qiFDfMrEWImWoeMTekDQS//9O86rt/PbCSBi3TzBI1Kfq3Gm1KnGdaZ
yNt8gtOVBKghWPXI+Cv0zsanN99ZnOpuDuhA9FVD/bmHQU/8Ap53LO+kxt5dcAd7
H3Q0paVm6hNc6/ROAzul8Qot+kmAd+Je/3/k0GCTHfe6JtLJFOs/wnZEhxFxlxcM
CHBDNLZKFgf69745PoEnguXuA0Si1vi2oZ5k+O0+6ZRt8ZYf/Ko/jhreZaQyN9j8
Crz8ovQ6uNsdhhooOPdiU/klXdee1Totw8JB8RRzw1LMdAjuhiD+HsfwT1lMy0jq
4g8ieTovxbXnGyRLdcuW7/BS1CozGCYihxyjKzJIDUoH14I3O22okdcdQTD5apxf
UrTgtUwjqyXsfnjCJbCOUbQ3JNv96morw1GOiacHaHO5NXpOgtFRL5YXA+J5Nj8i
ZgZyzahSHFOvczdZpESLAAQ6Ec5ke9In9llRnQGpJlmT4tfvAWa5TphHg4c+BaE6
u+mXw3jvq9DtzXhfxMCS+0f+okIBMTDu9zWHldD3S+jTX/uCUM5bTeB/+hPVxGx7
vmsuqkZVFJhwXRj5xBYkvN2jXwZ/bOC7J9NevIIiOUKlIU9PgGEMDQ1Nz3eioit0
XQCHuFXIMkhTj3UszTHqagHJXZU91Xn3/CpnPUWN+LVcYFtmq9BYHBeSMj72fSQ4
1AFpLq0o0sh/XDsU+ts7R8x/evP1bJVdHhag4GPZKwjQx3JTC5wREUAp1yPeYIQ2
Gix4UpmK/qRgSI4BsnALxbKbX6zLbNeUUc236hErRufTZHQXEqKk4O0cJw63M3EI
3VTVueMYw5Pvqc8wY8HBve/wk7huBa4buVl7Bynku3f2oTTYRC3aZo9YcvlGBWeK
E0f8XbGKBgbr9zA+JGk6QN1hEUlkAKYFO+kadtupm7ut7bcdP7Ik+IK4JbmaolVB
gBLUKrMavYSJeahYNl2Kvc1/m1i/pnXPFRbAOwzpqdIaw0k+FS4PeX3DbCEWYRzr
p5HGVcIzS6xuJQFyaOapk+Qhmz9I7IUW11mG1dYIcHzaG82bsX3bhG+yRFWu1fKx
cWA8/Wt13+I0ZZutGxUuX7FbXVhmxftJBfDQSLc4oJjhhphWUjMAoj6ByHp7+vnA
X7XA2ykGxV12MdOgWZKsZnpKKDwZgXswarWyr6bUF49F4gQQFTjMd/5WvyLmA2+8
tl3mEvam8va0akIFdSTkN1aOgJDMQgRbNsKRiC4MdemMWNgfFzfiqJ+OyWaApRM+
CZd6YvzDc2YBSSGhWOsL3ZkqL7/kdQLc8nDsr0T8TTWTrudlLIARw4zwYAhIgG5V
ar0KvvNRg7PM+Kmav0jet/djzpZjSnMCaMdtNIEMwcxytxrNC64BLb9CObfmfchA
TG7gBtJJPLbmisurSGYQlL7zOI6eRhRyR4F4Re1sXZ3sIt5VSIpPIUKqUoHSGPel
gtyV5w7FPk6X2eFwjVbi3Il5UUao/gMBlnYGgrEpnUbeiq0dnxMxtLuLvfiM6TAo
rKz2z21yOfsN1otYavaTur0IeCtQbToRNBkty6O9ISjOPXX4oUOJbrINPu/iDGIi
+dTRTP/w4hDqDW5JL9cv6aSpNqVojwn9VKyk9l/FimTHhsChwUKM7DOnH4w962yj
SQj0nkya1eDqZR5VMWewqxCTwH4MJ8WSE6zukvtHFw4hn8w0L49+UBUE3rLO53Sj
zHDDbcamFDRjKd4LmdL/Fy1J94/x8Z6/sB/lN71YJgkAGz6ExQTPb1AaAl7ZqBzo
iIrGYpL1Zmmima4fhkl8OgztAAu6EjVoAY1EmIQtaz3eIbB5K5o0+r4E07Rdpdfk
aF0WT7ciSUJZn27UPFRO4eJ5iwK9wU4Ak56aJhS7sn8I2pXO368qpqYccwVC3Ln3
YIKsPYMpHOTIZUAHaHfRLrIKlZsCmQZfvvMdJH+7ceJsWrmyCQDwX76fgsG36mgU
/p4oymW0OO3f0+PkYvGLeiLGfUVgkh+5+/IKXEJtXrT+nbyNgJdogQpCs785Kn85
3Vy4lx208msMLDxEu1PX7iAH61XcQX2hIk2A8+KWvTklRG+3n4nnb8A5PnVIZagK
N6VWu46z330z8iiNZ1AFwftJi6UctYNfJBy1uH20b8GPGUtEFdhafiF9e9pKbkta
eFnecrM5S1q/5AHOkamTT2QIbYcB1k3BQoNcdhx2rlZ4zBCT++/VyCXZNzTd5MLZ
4zMnqee0GjjxVran8yfU/EzOQy3TX4Yzt3MJpmhyj/sy4sTk5obp9EfEzlr0B3mv
ulo6/3D4jz1VGJvjmZMaljdX6gAFMXA1aQrlo9vYjh5uuaCj7/vUwQycxpbCned9
GXHkxZA6KfCq3AZ9DGdvTd17REnRHle6sDfNB4yN5MUaCVWlHoBgeOurYId4PwEy
PZ2KSx6y2RG/XRcOV4yMm8JQ1hmXRGaJkrDzVDK2g4HFbdhYJkM1hVlQZUDOrEEj
eSpkT2NsDElEAZ2IsDqb687y9oQ4Hcn51y4vtHEOPEt46w4/pxsWYSrRJWqMYMew
pDCHfeqeB61Gp/EU3jNR1FFJ/YYRK/JsZXiA9bWzC/BbJxGvalx8CYOzlqTWJ2Qs
bAFoOX6F0Jzw1VMQazpPbytUIgrIm9MYRe8oOAVuRC/5IO0iMOS/wxKW2dvKO50D
PY90dlHD6GdyVorx4heaMfw1YVXSC6QR4XqSzM63nzMWxmajXgtgWl3dTIbDzQv5
uIzXZSfe/J1AeNXk39TBxL1xyd8E1OwhGkEtY9VUhP7tMeW3+UuRO7mPlZx2/zyA
+yuC9ElcFspYkxK6QsQpYZA9s0TWLivMfXDjx7v8PqWxPqEc6Ou1LZY/jxSM4mKt
ToCUe90f9TpzvWNlwplKQ0hRuzVeh3b839MDAfIrZy2BX4AL/KHUU3p7CLOwrCQA
yvITsJwKuY/b6HdVUOoC5uXj/h5BAhT5eBQuJOfL02RonmsSQVTdfesxKeMz29RP
g4xCVq8igZH37fkeUhw4uCqEcDMOArRlsZd4o107a1qAivMQpMMTTxSIxIysPLGV
Jbwq6NZEylzeWKauACZ/ArHqN9+8zN00XG06xUDDFB1YdYKgpPcfbpcowDo7zlI9
l6vRLuFSjwrljj+BNGEh+izc2E7yq5WJ+LoVhQQWT+INlO0XWZNkECgK0Ghad6kN
ayQmeCUGNMWXWYiuoOW8gVGbwVPf0oPeY+b5O7OlHtI3Zx8jzWmlW61Hlf2gwKJq
CegmHQtUKdptHLTX4Bs2A89dq3uoCpLdC/ShRZaUsaS0qdVIDLTM5ic/l/IfthU4
ZGMhaqrx9KGHH251kgp2KMl8dcKcgUmoPKbYd7150MMW2BQJ+b50/7NzGTxK+p1j
VK5QSz04wKARTcfzPMNW1xjimwQu965i42WH+x+sbgrXbMLXVyoTRqRPzUscTj3n
rlqZClzXDYq2vwBrdoxyBdP61gIcCkoU05DaUNHgT5LCFKQan3BdZtlBDL/nC5LE
G3hMe5t0PHYiiPBl3ZzD2fIkiVCukZOI788ycVQWyqmEBaaDy4MK7/exPPEwADDr
McHhel90J/CYbQBTFTfQFMUnWKx18p61ywJSXL7lCmUbGswX10UC2bAkbofZaDI7
ZqxVBk6Sor9cRC1NW409ron9COwcMST1r6rVj+H+CuFrD6wkyXdiHA3oA8RXHxmU
i+RFbQ6W7ZPPfa1pCn0lX5juRlq9S4segyTl1TRQWCmAYlHBC9jBxnflyIpC6yty
Zbh2WUbIEry7QhZqzcmujfSSOpEBKMO0bZfqFqTBnT3fw8RALI2Z6iBHC0tYLCnt
qJj3IzBDX/ZZ8Xt62Epm1KschawiRaMntNPB2xAedfqARVsGPBWcVL9QGyTBUJZE
nePPZLfI+e01bbhbN9hRxpJE8mCdz4CRDfIYp2nqBwkCdimPh8RVaz8yC4B2Coda
MdVaH0qxzVP+LJ1471myOy8gm8iK2mFm9C+Nt7nKenE8uIBID6NqF98e+o8vis8C
U7iCiNyG1gYZpo3IKj14fpOz7F4cqjeP6YxqMT92A2rCPd+0CKeQsrPNkllgjmIE
2+ygWM3AbG85SNq39v/E+sC/4LmzFdGqLC6US22EPm08SGUlNP2C2gBRXNP5A4Ws
HLzdwDkKadFVVYZUgc7Ea1QsKeF86BFGAtJlv6nQ0EsxYsqhlVmLu3nzRwYJAjaI
twLfCGwXJEZzkgev3cQyDp/oVg+Vuvf9f5+5ZydldTeVR//tJ76SSYzNLmyqcmYx
roLKLOCOvp2KBKReZo74KswBn2viiRn+q028UipBvPqlURaSggtPhs17jWXIdGZ/
3LiaBS1hlAIrcpWbjWK+XgfzX0Lde4atyh4KiMxEcgpTxwyOsMgkS9Q1ZPHfrAFF
AXP8fELfWP9IAd3k5XuQyHHvyCR1qn1/UJVPxOLho+CZQRQEFYu8dPmeh7Ni4tk5
0MrFl7thAazXyvRzwj9mX/Xzvi6fcPSVaHO6RzsU8qNv/LOmmACMVb3v07XhpYDp
JjXQvu+HvDHw64Bo3qOvi2XrZz7g137IdRYnVAogXip6iFVAkJby/Oe8eQvoPAxQ
m53gOKZo4npeP5CIt+RkJa4Uor7chR9VXewOsnK+Rk+hdWbIKVz8chp5UAN34VPF
ZxasWp15G+xeqL9rM7hbkx62dbT1IcVMLh1XW/wyACVOpPVxvn4oC8iZIHqGM5fR
mzYgD8SDHp01icyuSj9fJXhmamBeCcJ/Re0FEHWBxhr5x8pWVRxTtFUuxlYYu6O1
7WnWHzO825TsstF96bFP0duyubsRJtmRYCv+qU8bmTR5+wKwOOPs5+6fT2KRp7or
2aP1aEytg+lW1YidiBSCWO4Pswv0Juf8CZn0OAM7AEgJfrq6YhcyLzVy338S+RqB
UU33JNboHUflHzoRhZag7M3XByCJj1eMX9RXZlzoB7coECUWfktfJoq7UWVecJaq
o5gU2YjHAZy92A2ioPkh1OZHrQk4vKYTLipCwyLMXfV72agGGcdbeIJqGgOET21z
bOmBfxc6GhXB3NDf5TpqFAG4C+D41uhMKtNZhqanQ3EHYiImxqquy9tgqcjTrTC7
vdF5WHpsevpYA42gQWS+u8eHUEFDSTBl/9tdV9jw3GoqAFq5NfnbDeTJtxV9Vw53
sYo933Dp0a8GG/MtginR8j6IQZZ5hoT9+h7lgKHiCQYBN+6qY8gnVeGqyLXMNkMc
2F3OL5++i+Xop2XiM5E0Qx7T26r1wFu8c+iY1HkJyGNzf0sXtuZLuHgpirtT11HK
mlnmxsYue7jVX0SqtSpaG5q4CgfbWFB09GxfIfnGhraHztoJkfoOv2QFV4LFRHBk
PxWysA7li6Ulbq2xCYjG122FUBxRuxQsreDs8X7UPoUSmBuERNYVxiPyvdgTdLSA
UWmsEwmIX7Pm5QsEm8MHIVI8LO6Uyir5vOLWh2cKcszTNqX3O/EeSX0zgA0nHTOb
if3UVVwNFCJu2MjiEUb3KFVnLAl3R9xB6BWP1yGV9KC3GzUGjS/W5woZnk1ArVNE
CvLloVnb9ooMVgvCvMKgngzRf2rG99tq3cgvDmus9+45Eo3vPXF6Gq0WREfNWX/b
fji25j5Op/0mtRHoEsVHx4ZXU+FqG0a1pjYV002tHbxkzWclkFnwUKobc7YrFINX
bswBlDMJysuVrxFg0AcF9DTlEjNVOD2rfJ+lIci4chaVAC9rSjve8fgyExmSPZ6p
MqEY9Nm8A149j66kxIFphoh32+EL0t/k1DvAQy5zOim2ZdlSbBo6VVJpy1ArWDId
ABcoms3R8u3qXgyPR1wC1meC7WkuxRs8+N/q+2XA2iKcWq9kLsqNB4YknRqEN3WV
RUStnyTUgmPg1g8d0ifLOBjYcWMGLbiPuctElnXDt3VLW94KYcqKU/lk6J+8Puy6
8PwVS7jeQCOAOjjfECgYlOq4+a3V06sgFNlQ6NRyqwghuYXkwudJYRoxyU3HatxL
bRoqNsgi9r/wBox5pfbPxGn380ZQU4HHQZN0b7dCDKup2eL+YfZx4BASZ9JMlYD8
1F8nOyyUd0v90D+C5Xel89gzahx/PzQDMht5ccaw4+eylALq/eSv7/O0JnGsv2bT
wQG5qydotL1AwLQrOdeqVRZdP/xfe7ew0xpW0uVLaZO4cy5CyttI1h4Rmv8FsKIY
Krui3EyGaLelpV50VB9bABVySQ0JzNabEqb801oFo+c875KJvsOI2PwbqkpCi1xl
8XRJo/BgPDJrrGTQ/LD6Q6dZ2SXfqq0oNQ7iFfYy5SN17mrDjj1ElrKwfQQp+BBY
uPH3JUimcokS6Dlb9hMYkg33u+2MWYVyzElkgVmSWBD26HP9Fb1WZVgGpaiopTBY
2ksuO/xfJpFqF/rJj5ZrZnP+uhBOV6ksWb63+327+Iqx4+REaJh2hvyn4VSN+VUj
gaEhVebPq2NDtL00RIXsmGu8wkxFSAsKFHW/qOBoDlMX9UukRG4dE9sBjKh/V50Y
S4wtVWdJfJ8WZWLPb3F6W/tHyRNF9vxqC1sbKmGS7/L7SyBZUNb4Ws1r3khR2n6q
msJRsdaCYyF7aL2J7lqrNUAZgepFqyJLz2Ci6xwsN2tcT/UR7vzNi+3hpxdTYnaH
qk0I4FxSjocDBbLrF3hoX2LpZzCmC3O9Tj/t1sbNeOudWEWdEgADgKV3a7dlAPl+
nTa46mMm0PukTh5fNacnlp33gzedA1pLKsufmOuqaLI03HwQuoMbizofO9Jh0C1w
upv+rFtJyiei7uL5c0aoYr3y46KIn+BrAxeiDeYwPMjICfPKyQWN2OYq9B+eexP4
mYBZ4NsFy0sl06iJUGIpvhYSEKKnTWwhJriJS6x8tENFKA6h5u7y+qwHkzJl+VgV
rRQeJyr8o6naNZJdJGvJGbtoU3MEhYyfrVYaMCvzxMDRREaibk5Zd8cUVJL8ER6f
qSu/VWZ5mhi8PN2FnMwZi6J4QxedumV6uca2UZOdXT83Rp8IBWhNHe1m0hfr0OBX
JdmSK/vIgybeY4hc0S5XEtIFuitc2aB4jp2PVmO/YFE4epY4HswCxH7ZBVtUGfeW
wpbZq/qcgq7eaYXf9ouHf8cHnLmfuhpwQa6ssOXDiGaapETZqHOmNHA/XfsqbaVb
TEcpeuO8h3SIHsEJg6GawT7TyFV0zAACj4P84KJ5lQ56qSZllM6n2LQ3CRccJ2UJ
GGvxqq+R/EQ0R7t3od8aKgp1S46yyl14KTHiAwKGKDWgG3bovCdZhMx1DoeaVmMJ
sV/nkfM5XmHhbVJDAxm7SG7xX2ioHSvX97538tjSUDqGMLf25uYbyUk+OL/bHjuS
qcveic2yGNMcyIgGTVaXSZUKQnjVjIGe+Wo2pOf343/SsvtnmLKZoGhZqzs5z6cZ
UAu8J05fdOd8cVQ0zwqtmiq8qB4X/PcLSJY3ZZbGCC5P49Nj7Tz0iw8tKJ3Qvz/G
zd3oRqBuG/GCtjqxtDjyKMljzbQct3L3XyXf2+zibqk1DSYyhEBj/YDyut6aVnvR
JRRfobEk+2CsanpiFXcj95sAiFt9Sy6bCA7PPJqvTbxmNwBohqWw47SrW6OhsjWn
IykVj8MeK7A6KcGTiMJDPSL25/GTFH9G1kKrP1idEKBMpFCWNt0O+loyUCt9OFEo
+vzE/C4mCfFo1rbSAluTUIdFFsKTDXWBBdkAQid+LjEJ3Wz7ka8dF+VIZ9j5uZeY
XM03JxeVpnh9o0W1K6G/qcE1lZsEfb/QsQpnMPON48+GRxVcpc+lPt6sfDwjZkF8
5grv8s80iDSTAEBSFJ/zuT6t2q3Tk6jGLx9+p7TITLWE1BZT6B7gSWE5jpyE3Hxr
jyx+6b2K6foHf/UHpFmAMnJwKkEXA2dM7QXh+sD2/NVdFk5YmshZLgs4T4NwMbKY
9vTJgcmxLbYk0RVCY7CB5mktLmooBdW20X+0Q+zDa+7uFvbe6najnDh4JYppwgyV
WHoOmRDu2avPsWfU6bzpwBy8+XV2Q3UgIJAiwB4qUVb00DkUXe/tU9CqdiD6LOx2
k6idD+ZrGslTHnxkoI0kovJglXwy3CXd/Cr3GVhMgpF/kMErxGd22KkDDI04vDF7
mBvX/uJclEuOp8tJ24BONFoYrZ4RIahUgndeIcTGHyy5X4zyGVLhjtpsjT3U/zT9
yNPZFWLnVK0K7plEvmAYyzslOVvk+eu1Y92PsRx1zg7wzsJ0KTnWoT46zjhD+COI
Giil4rd32vIfaJSA89ySeraSpcABVS/4PnuvWo0RAFDbyubQfnOQcegAMrOXXgXH
/G3w3zO3zrtV0v+g+9+frs6w/eLIM6A+s6wdTtF2NFAlLRHYwOUBldViI6RF8afO
618tWwHl4i4gING67/pbgu06ZNjZ1CZBKK4bW/c6FMvX64NrybMNFJh6kCkBQWMO
KlqY+k1VvfthUhuIlFcOTXziaRsioLgwlkE3Un1Axx+8OecYveQavYmOzTX/zFIs
0Lv9xgZxtJlOWbkc6NUAMGyH00ea8MXHp+84WlEkF/oHO1zcrOFXHV0goQjyNSHb
eXAkfyhVczj9yRNETmmfK9hk5V+dzhmvjY3cs39vQU1wCUJdWuufMitUtF7o0MKt
03+u4uIUgzXVDfKcmyGbatXpzwVjCuzKMHC1jyt1mn6PgYL7dzgxyUW/aPI6ODLL
d0NN7MJ2pJeXrUf2CgNU3yOGyNQatJ8G1jj7aR0+IEsF4/YkJMK1rm88FP/drvjS
Ez0yx9FDvVsryyPnHQIs5/7tr8ZH8FOKLA/TAB51/FkRztwGX3lMG/3emAiBkjHb
T3s6QNgbKCjzfkZj2xTzlFx2rfdHWqbdTmMIi/+opavi2zv+ef3k6vbOcM9OGRBB
z+ztHis38SqrmQ3PgDXFyOz2gr4iDf9P57uRH5G9gwjiBTyECMI/NerWPgyhmctP
vaFviaZqE/oFAYDTOCsiEO6H1yR0iQddqjIv3OTbP9pj4BCDY02mxLIcCK0IaNzr
nNc3nT3ezD2ObXCHWmu3nAAb5KkBJI0XhIGtylemGX6BNsDyvwd+yCYvYytE7P4L
3BpkhMppwhI66vWaOP8A0+3gmPoVPN3fLkUENPWxQTYuWZVBxC6HgcEfQnNHa3tb
gOgsXeYbwIBJkJPMeysXTudoMbmVm5F0fvtqYBkWAltxOt/yzwDS0s3mEfCikWkn
+QwyJ7JjX2EvXyt2+B4w1mn7Cje8mw5TJDYms30PL4mVEWELI2EfOkft5MpGwvkp
sr88PTG7QffMsgJzqlEFWB6OP5VxioVwjPh9RR/2Ryp+GHkyqCDKh8seThiN8pgn
tuhSVss1QtuUYpg3psuKJ4e/DUqGdGhI+PIgOVmOUBgIUwp82+vgDFOLgSPyB2Tl
IldCOTOZ2mfZybpeAa+zJqMG4Sh+iciWNUEdxLNbwwZ9e49mkkH8RpQXxkffZESW
7XfXLpJvaS+fy/NuXCDPySEqzDnu/N99ewnJMrQ8j1a1XETNKZW5IL5F8v8L2oDg
/5QKiUjsPvotE4jRSOArgeIHpmuG1dgPGSm817jSciNCWybW77O06h8kvHXlHDns
aZ4FuWgApAuNp4u6SnI2maEeWx2/0pVaTRvHx4LgSG8Ue6ytrf+9e+VqtD6ACico
yoojUXax+vVI4WCvozlr47jNwuKz2yRwgGy0nxFPoWL3Y7ZyC42lXklwxmqvkAKq
RKmXAldOzE337flj9BAA6J+FlfDEmIkv47BBlufgi5Cu/8gh6kBkULrUwpF0Gm69
Gw2TP3oTOKDlvyqR/EpIWXnZKVnHwUIgKD2/RYHwKWMln106l7F0+0upPlMMoYxa
NaA+ZtbELifUyYsO4gPrAqi/WvmM6M06gnl7sFDQ/6JieBld1aa4V2astPQsJG0E
f7R1jPm29dc1fyggF6DxJMZKzwYXBtIbJZ9PzCNPPzR8l+GChpxlKu+5qQP4dq9j
6tP5MEGPp0P5yxrjj1tBs+e7YbzfkrAJmaGmEzmDqj1PRkLaWG5K1DB3I6lESFIm
P7dlSMINWwNyVJH9idfzyjFJm3vJNyHVa8gvnFKx5jvqV6qI/Bu/kr6MSsk7UDls
A3Xuyz5TglJF9KcT6in6C3i6lGWHSiqWvihRUYWK1dMnktuDBXUuVsr9Sq8kx8wX
odHB+e7vOIYc9BNZ3SathtyUhMbqXtU4vCHFErnxpjnZr3twN7Eh6WniJo53AZKH
LA716IP3s5sevrSAt+U1H+OzOn8AIaCJnjN2+DAcArXIcfz8dw+dEIFzzO4xwcOw
OspsZqZ4VWUrtWzuqHJGBYcfqjvMH4pBmUAHn4y4Me4XLPSKA75EJsIRHHGpIr0a
wAM2pmCXbUesVOoHNh7l3pzzlf7bU4AIQR1N8L+rid7rtoG/FRSESagUtEYflIIT
/SY/ie3pPxM1IcrjFMEQwSUQ+AIa+gHBcV4g+UM2tsqfdUqZXTO9kmhc4x7p7aBD
HMS8PMuF68jpNhTThYry35peWfWXKra8qSzv0Zzwb+fTYnAaZXnheyFxxcuLoSMb
dcmtjb7afu32Hx706hUhNmNmLIjzQx8mFahN12fkCd7pQ2rmqAUcZKyEiLBuZq9D
JVodZiYJFF+VRtSp9CQOOCgBNZ3/6LAdwXrnlJsr5RXR7k7CBDeiNxQwqff9s2vA
t+KHLxe/uhAPNu94LZ/ZPUvfaghGuBSejMIh0xsd3damneuh4ORzogfp7G3q0HVh
jzIRC94D+Flx//m/0lEQTu+jr3YrkivtPEvByMS+PsSO0jw2cCWQMAz/sHh7K+3A
wihlemmnrqRexMLbUhjO2hJK3sbm/GgkOqcQWe8w/tN0Kd4csL8diP34vQiFPm5e
yx9MNMIwPTJQcA0wWMFd0o5Xh1Nd4uzJgbQBAYxi3f6zaAvTD/vFGfBn2mwtU7F+
vEBE3rCtnJaRPk2vrHBx8o06vnqqNPPANpWqVzaWIce5VBJ7hbiy8hWmu/WwoG+c
N2YpGtzxG1W96Q7G5PLesRenjWJA0PmbqDKqW3e7FB0Ds9nD5qFOKlK6/uM7B64A
90tyF/fLd9PO71odsFGbzijHo92fM9RaD350ZcPPoZHWAh//7R8eI0LOc5GwiNJN
Yuks8SwB9+4ds0UYDGXBMAsbXSZr2pLpxFeDkbJDhIwDg7m1Yufh59Jm/zIrcPzy
YMoaTiE/H6KZ1LamXFyNwijrRSvhLHfF41H4MOHzdrdYDt+5gfNAx9NIJ7yE+Luz
keqaYuxhI2JBr0yJDOM+6nu+QAzjVq7kXFKTV1oH/MwhmWbYSvY4uXLCDLWytWHz
Gy0kOCw0JYc/ERBQrpqOigXs/Q4dEaQl3UeoPWGMnYm5CRoLXgyoisDGRXWy9LvO
tqMraUDrV19K+C6Qv2WSGJ+kj4eelOGE7ukaHdaIoCB7Txk7SNDUt2xb0Clv4WtC
zK2uH3PViAOkjAOHuPplriEIw8FBfbgaB7VV/TJML8u8GmZSaMlcEHGz4y7nI6Ko
KglhoQjBDCEzy49rQdZWJKAfaMT+v5AuNWAsCyDiaCLJBUlm4aA6q3ssaMsCJ/sV
Rlkid1/DslIQTf3c0bwECIgO9wqY8H82LRPwJmAyiMfWpIQVpGtzZHCtvnCu0l+d
/02ASBYdIfBcpbXAG0zr92+HFL7t2LEpA3UkNQs9AsddG39caqakzNgehP1qWApc
q7UajaLMb4mgCc+QBBX8bQXS+cjffqnb+ikpCa/Zu2BzjHYlin3KVRsxNEzj3IlG
CSzoLnx2VPUmvwGC9yAXIBRkN0zkEyfHHWNOqUKhluGsMEt0ObaB/ButOwVFg9PK
igIU478+DmOUCsb8muahkb2D6Jvtw+1iDybfzk0GOt3nvKfKgjVIhuFzNFFToLy9
nX4C2FKECwHzeVph6zrffpbtFADftYvTwpzAJvzIovng9e/yu2QBANdoNgHzVQPf
Vz/qF7Fv51PnrZdNALQAAWHwP5nrYViZZ/NRoNQFkB4vwmE4sR8aul7gvQL2Ou+h
rXeNS1D44WkAw2ccdKNaIuBigWNgiH5pfCfZtu6k4ybpnNZRa6C2R+W6ISb/g0rI
eWMgHMimJPz0Nfhw0K/bAN4SfjY9gvloZwHfjxL3sNGH7JSPo4X8LCUp4COSUThQ
5cEEXmERj8PnE2HPEJrgSr+/36QxWYpYK3QWRTtDMpKnnnK4prBjWZ0fksd9nBmE
ItSgB5EVdiUBRZLbaXUTjKLqLTf/89x7t7Jvh/SA+7XI+eRGfqWwSzY5W+W1BJ2J
Z4Xl8T2Kc9ud0ipyL5EiTi/m9X4shfEpTpepfzSYpKCkJyfg85l/0trs0rLhErvr
pXpvD46py6PDIYqk+8YqijK4CJmoo7EIleMS3kltL/Yc6OX6bJHwwAue2FFe1ucp
Jfhs3UVLUjmruF0N7qUCjGaCB69CUhNHkcMTsKed7y6xSKHq21eA7gaFjvQXXSUx
msyDOnz1zwIh7LZ6zoKVRcB5tROHBcyuSS3zZ/Tv1UjTPs3qL5E+J7ue5MW819Jd
j/xfijWG2+ZE+25Y+M7QBCkcbBBQr+oAyzehEG2LTC0HIn97BmkJRbdtyE8C9Sd7
7gr3tn3hyMNlKGKMr69lw2ywIvmqzkpqvLrVu9laQMdoDWpIX8vkK9jCKwYgGJdA
Qex7UODA6SJ0mWUUzGW9oWTrlHqkEnDGZ31q/7FPk0MlCyHNe947izw7t23Esdog
PW4IOMXLANMV4UZgrV0gVzLEJDjNAVqkrML/JH7S1OpZaqoDCnjX6oe9EQxOz7bv
ZqvsLmCD4aXl2v6ODJ3T69IaTzjL/hwBN5FVGwp6SVPjOmjhnGp/Q917JgVtsaQf
UU2R24jeJBKdK2a9xR81OFp9L3hLOAjo2F6+BgjJSHmYY2dyB1IFRvPXLMmEDv6M
TPdLGz7xayPLzb5C9+z9o0xWGR9H4chw4+ZkqjpAuVEricsoLZJ0x7OceCD7vPkn
JkSaeUvfTySpLdxMjU3xVNaO4aAbv8Wqx2koPY/FSYcjMBjR7j8ij8cZyEIqz6E8
SQR9MwCFg5Wb+1RBkEDtkViqNkzNuFVhKTOgakx4H8t7D8jBa8VM8aOYKwLezV03
3Ip/5WKPs/Uk/mU1PFsfX50icrkvi0zxWRISxiBNzfrvftBzzxSdrbVysEcROYfu
NPhL73bocV/WTpX2jwECk/PCQS2je8gDB3Pe6pyJPYvjTRil8GSIXkrVaNHF04G6
KovkpOo8hjMi22ByiXKZiwjkbAHjnA/skHTGTUjv2N62soAjMS4kqoulbPrYhvLL
+E0sMMfhGqAag8Ek2xNB8S0YBbGcoRt4mCyM1C7ULrDSV0AsBKQMyiNfAA+HYXX5
K4AEAA1FPc+3KZZfIudU8B1GGVtaZ64e34ce5AA/4dImX/e5DKe0PKapr54zGfB1
BwZ34/B2DMlvlSc2E+aNdCSOqYqg24+E2q3/vKuRGwGkQiqAYZNslJa9r2bhbNnq
X9JSSXE9ThlUh79GJ4t3N94aGtAEWAJK75H7D9Zsoz2i/4znyw5mkJVcvlW9JBLO
BNeqXiw4i8a43igT/AqOWgeme1/iKTcREQKHXbzzCpzk18D0PMB4/qRcaXt7Iuyn
ScAYXBgaFa0bqgNjI87RYYfFhZg2Sp9J1HXAmOLiQ7miTRJBRoL0700NGVQHT4C8
tMokhkaS6MyIOI2qpcktFTtrKjz7lubbueTvkH7nUM8kWLPsv3mHg8GJr0RRbDfn
3mfvwYNoPdyvKs6Am2i1groQeOJhkhBW0Ri/GWbGVbUZYW4NsbNJwOtPgYO87Npc
JMyp+xA4MVVMrEPcSAKN9mjtZBfz4onc5j2k/JL5NKpPeqyetVaJ37Wug9m62JWi
Ei0ckydxiFhbHgAfYl7P/dsy6Lw8iRyAJ5m3RzRsBawKD2Cewj08EXPYsX8CE0a5
Vkbpb74q6s94D7Gn4T29fjLODycefD8tfn0QFc4EQUVyNgpIriReq5cAHdLHSAuv
VQamdixaKCbV0j6fOr2Dnm1YnjS+zy8J2GSaNfGdFqNXeOJA+25ZpQYhte/J0N95
XNnuJgjDMk4eu+5ZTZmvcj9fqKT/P/dijifnF3M1tDJr9OUHG9YagXR91YdEjN4U
36qAIvx+a3Prh2vUvL2mBu+roZQ1lvac5YV1tke3qA+KIM/WIUkAi+TTxhimLirn
pjl28J6q1RNkBp0UcjgWstaUj8vmCzna4h7KXaLXY+SdoaPOPjzMnvT3PjQ10cWw
Ia37cVCXWBjgVOpjCnGK9CQn4jtEE0hlzKIFCgQ0EBOMrXVYeu3CPSX9xH/pTnH7
A6Rx4aHlZE0MBEHAky6s8YwgDjMjtb+uDShBWUKlzcMdSjAwyCjo710vY9MXkIBm
6COAJSXAd3i9LrpCGUaYda8HDEOeEn9ZG+DXVvpWVQz2Kup1R64wHl8OrqEKGk84
ZBAqeeYNZ+q9+h83eDwa0h3fd8YoYgh+dMzz/QGG6o0BdCfijfjTkBFLAYnjq+vy
DGVEbWFMZmZzsP+WHp3BNbQ9sJw837XkkphKDof2kow8hJgweIjwjDocFvvDRZM+
7/AnuNClmBKtD6OmIqAXva9/3DK/dCpk2zQaToQqzgoRGFbF4mWVHEv3hLaWC52k
N40GCnff5Go57EHNaUoPfj17NLB55HwLprihv2o9cwZLXBfoofXN0qzyGbth/Pi8
qFr2+A+dADoOZscII1qxXnao0qo1MC8/QpucBiT1cq7DP5fwAVxLiut0gtmO6KOU
20krCKAJPvU9iRvhUat1Q0VGWD4fy2dXIngnmL5Mhx8jzCUfPz7cQn3Fpxgkf2kl
HMViPpWmLAmPideWpvUYICrW/uixBPFSxTFBHYzouNGg1++WBj+h0DGoHw0+F101
kI/9M7Hqa+tc+8ltHY/OV2NtIhC1/PHwW7jALhiJ/XSDEzcDgwBlxjW/hrguYYQK
dxAcN0R6R8BZxTSKPrqWk9fNpFOLr+ebC0W9JNEMlKhBcPvJiDqSVV83AXMyjiUR
d3asj0FUPRGd7EuAbWz+sp2zRhYuHMGdgxOt24fqmBIEPLnAKPmpbfEJR+IaVYUN
jQKZ9SL1GwHySyJV2tLmA8f43cmrH1wHEopB4ADWtun/0ve+FKOrynrpWshdg2Fh
IubzOJ5f/seycMMOPeVrXXc6DygF2RwNzofaXNEH7O2xSdHUryjYxgcRQ1hfsoyb
OY1aNSzX/GQ6M5nQglMg4yqHWCVl0NGQjr930y0qVmFzgsl0PpowSECXFava6KyL
ZRoBxLNSvhRNJ0JbJ45yR/JIsq2E+20rl/PmG6S7i3nOVvZIUU+DF1vNgeuqRGzB
6BTs1chz60ZdMCSUDkpI0rJv/2tw7UNAhJiX8PyFIp40Aatcy31GVWSY3SDo1S2D
nOZ4GQ+QRGTvFVlFA41BBmwMuc6yNkJP3052JoDVwtt6izeYqYyKMDvt8bqmissj
Utw0N4vsA3t3IPDtnS8RIA+5U4qxULYqtIfepyM7/6LnE9ZBYDGhdXzZHmb/tvgV
MJmoWM4SKh6DQP7CnpAS7oKEZxLpHTdDLrgouAdEV7ccHZY+V/drz8EqGR4pLNhP
/n7Sz/QtQ8Ssfco9KuhNdenM7YkyhUW+vV109C9XBcNnovxpxr+i4fTNYWahWP0Z
MQFrYQUiWin1MstD5sFbLDuoEggv5UudRILpRvP2v5ttQVBIZmE8tBJljBtnOMUl
jvf3hnFgTWNLpEfd0qEkRwAwVR8HqZS2OtHwBeqgJq3RiYPq1BB5cWMKlKT3zUDo
CFHCKFrcoJfrIbtJkUDUhamQNiT8Evh39CGz07oDTCmGGwvNIHk+aTSqk6SCihiT
PsmYEQVNzDtSPTBEl4kowtrYy4N8gReUXlhYrmq8LyHPpkk9r7PIjirr6nQLiH2v
ZkntrK8WzZSxnsscjyM7kik94FrdBXIpK1QvMMuYrLDWw7NOGjfSamn6TDHvun7b
RRou7nqdQX9tWcvBjyWubkCJN0w7Gquk6Ceul6dLswnfYcH0upx8bgeSkev8pKRe
5PdSJZpSIqLByXngvXps9gW6DXIoV8mGEgs1C2I3C7N5S2Rt0bKdQun8fLikPWum
YD/gbK5VX/eDVzZOGiOc+NxGaHSIvCXV/DMvz3n8rZeubV/S3pGOV7xZrKrvOaCH
F2RAduSSlDZ8GCxgy5Bzd3um81EQsYm4TxX1Kl1yq5ac6vBhhTFKnibYcy2QpztT
eT/6fYWYfcqeuLtCoXHxexqD0PiVq++VUJ/amaf8PQ/iB8xCFydGHXJDcy5san9z
tuA87g77gohkaVuX7do5kW+FNHkoKAJyJDoIKbZa/oUUvBLfdKWCEd+6qMk2ZMwA
O+iaV60JWMVwh8cmNZJNWEHQkJSrpXPIAcD9J8x94swg3Qfa+fK5KHgbtITCYJM0
+/WQr9/ijkiXa0URn9eVtAFcPmYxVlAZ6KQfzLEapTkrgvrPmZ23V1IPg7HvDP7T
JcV1TqQNE9gWilhA7YCHiYfehtT0CClvzNBpZ+JgU+cc8bVcBjp8f4BjAs8/uIso
Sgcy10nFaJ705qNaimhsLKPrKL7+zALqljjA7jLxDgiju0dT5SLJ7fojhA9K/mIJ
mMPvmsI4ZL54ecb2eSAb/25zQg+4UyyBu7l9lgxen76rH3xqCv8QMb5V/Zn0wBkx
va9xUBocM9ZSzbfN6aIWETNZn81ysNPob7WyLjJZiA8Tfv1CVeYqCo2lZ4U2A1O/
DwDxygDHn/vMjL01NtFFNYHsaqfdDP15tZAp7eV1+dohSoXa2vU4bHZBJ6Tk5DUR
VyV1a63jeWWcTCf8b9PhYN1rvYb1rMmXLe+E8+IKGjLsQ/veEPeLOnlcqjjdzns2
lDLIntSBvA8WA8LPy25M6Hp5M9vhhSMKsAOZVCknVP1Rkw+3e6M+Kl1zb784JcYo
1E1k6nDgFxjIJujkRmtVUGiSwik1ifVBeLaeZ/mT4aq8+ifMA6bpcW4DB465lb4P
K4qWPFJbmZZNKVVgQdJw6KDMtCxq/A4ZwViOEFika7w4Czz0b78HOkwdAAt3mWGb
XDzGS3VvY2VUzLXcAqsPfXnm0vlNQNeVZYN4WoNTB3Tu+Vv0JZB0Az79YTtdGuKy
PyHsodzPCNBftr1XwMHzElEHitC36oebveFbvLbcWgXYaaQYWQj8Y2OrkoB2sOri
qxX/iht/6mfac+QJnmi5kqMkysOfBFnd7plaq7jfIm1w+cnzLx4+1krpLd7A1DsZ
p6LmOUb28Y3gcVFPIEgoSOiaGhHZAXCSP5zaPpc8+lRR6w61NgQ5eFbm0Sxygt9B
4e2cjTXik2HRvMOEVP4ArU8SwQb3e/uWhzBl2UKH1QIAAJgr/koAv0YOtjdS19OC
m3VCAdT7rUPs+Vko/YZaCJIyH4/cEilPn4BEOezhsIciZ6Km306LAuB6GeXoFwwM
wMqfwURfoH+dyDEhrbbBV6Myge75f6Ri+0cPiIZ2vuC0Q92tsxuHpMnReYDNqxtS
359J7fAwj3uueChoK3JXHisN1djNTEhU6U9lUbqGYR1QRiqtwC8MpJG+OhI3K9Vh
j/7csGJIOat0JbKc4acUmVTOFXnTl05qbsosLWrE5qgp/71sR5JZOY+YHqQguhqF
uqyYod2XZujRwyvyWxk3LHCyf1Ye0CbrKMUy1lMYkUkJk5c4a7vtPFiemydgPASN
sR1s811+I0j2lJmcRHPZ1HQREs8rcdOeG75CtYjv2TTkdesdFEsgddVm6MPIzwlH
FTuQlD5LePcq5RtGRLW8kEXlpJxFV+ItyJc/YE3gvlrNIIUmgpaDMOJYYnzbnzMd
gGnPyiMAGLTO7I11sEmjlGRbrNkjNB+MvCKRppMDsdAJh0fq43b55bnvsNyspT/M
mNaXqDWxuwUlJeynI5DwanC5rbqtwhMrIksfs/jx3pe8psyQL6P+0x/fMUIZqHnI
CFwsH5Zb2fgt3LCT6FVyX1b1JaIcpbnOL6Ly909sidni1PreaG8gzLCLV16FcbKz
y0x2q8bf9DZp8u7a9Tu7jHSsQ4chuhQ6i6XdqxgaWG0dY7YDzFx4B6DjWcQ5gCaB
liqdkj8F8nQ7tak3YtUb1efGiXP3HONK3m3LwfHvReGvtkE6JcQEsQlRF0KSYTiY
Erjz0RPRUo8XLsGHczMo63/5maV8WcfYZ8+WVpuOwEjOpB7lj/dH/keNGW23gyRK
Zz02LwrS/42o5c/wEGu+wtMX45AbzfB6RXn39+KQBefAXozwKyHB1vjF2tAltT7c
83xU0wGEJS7Dcccn8DO9L4lRl0+e0jfNBNIG9elyj5YX0Brt/9ltnISwAaySW4EH
vhE09nZbktIhKst8jmrlZb5pLIkU3N8yhDJWxxNiqMpFj5DWFDjiMDOe/8G9s+xf
gQPqlHxfuskEw0Lp4DUgazmVXEb9ksGXIuhPThu5p1Qh7MVxYaXWLPFCatfSX+eP
K8qKiixpPrfnjMFQndpkNeg8vqY9TIcK97OxfV7v+KEgbreja9aMhWNii42TZ8hC
V8jPOPOuxCMiNUeaxQBPN3b/CFyfh+yctN2chzGBAGoz+2bCWcn5Pfs8hFQHRK/7
fuBHBqYXErWfYJYkV5vc1Rmv6gLr56aOiA05RuaA0orUvr8gHGptdeCDVX2+HoA4
QzMyDRXatrvz5D4S/8vnmf9l29s7Ec2NouPzoZgwAS4sVkTLLgBA122owis5ALNM
hGcv4aVM99qztPsJX0adeykmruTmGSWsIA/VxfzVXdBbPGmDLtoopPgXZmydGWTO
oJ6uf3QvTKPsbwvmcF4KRqkE0oNAUvlcVIi+rWNgP/J9Fyd83ivMu+eVcSK1+fCe
5TKbKfdtVWHmoQhz0nwc4otI2zaKhabady/kQlcoUJbWHCmo2AhzBRQOPrXd1y5u
nMafKrt4HkqDcv35umNR3xV6qWBP3g2+pd7ohGt+PHz8EDSL2cJgyEGRmlOqXQkf
RuqmPlJPDcm/9PpPh9sUq0HldVjV2eb6fq7vxzBqCNYSiV8XFBVmB2gQgqfszpGm
ANZc+sHfINSiDHGIGf22pTZLn/UwC5bahctOUPTGHC5BLCYOn3WJolCWpZP8DrJF
5B36Blj2TFmq12URLb8o7shW7BsztD44kuNoFfCoiF06I3gTzw/rBr6j8lJCA3oY
5w+UWptizpd/ApUhDk3klQoXTVRtNXrRR9yzsCAtMcomE04CJ5fHpweXKaxZcjc7
MWHmnbynufn9JjDGD0HTDWTjY5R/eTzqQRPnNH/ZOET6OLZzORYYaRwJtJ75TFli
bkXjETUKyohrP0hhBYHgfQy7PYPvduajdE8bUEoM9oHwzztgh0NjGAklFTNyVCtc
TLdMqp4/lQhIlBdqwaQTL8yDgk/CA9KrFtFcGLO2FjBbQEpzmxetAUep+t5Tm/aj
ES2HjBSxA+G7q9fbbOBr1bTLC2P2oLUB9ehh31/JMccfBLB9Ol8IIJTasaYVa6HQ
R65j1Y1VAgOX1618c8MLUf6eOTSlHPdSOhSp10yjecqMM73zucwKDv9HEeDnVaGG
K8214yBFTLH0aAVNw006uaojN9fehrHirCgMIsxav6UN0U6u8TLZR1T42lIlc4D2
qQDomdEPXtADfE3a43P3vHjcsRy0KPwZ3LHil7awPuR1B47glhfFCR9Fe6Yssf2M
I05HHHi+oRDWtbXUu3Y4W8W8KFzHMxweZ+P8aGQf0/VO2/CIZLSP7jwnLoEXdqPu
jD6VKn7Z/Dxke93DMpUeCml5LAwFm5PNYurBplTC4yuU1VtgVnBnkQrxg7lNjarf
N6QJGk1nxecNfxcWOxrxUnakCSTJcSxYlc1QK3UJgi6STBH5HrU9PL5gZKV0zYex
5eJIRwLjtphiTv7OUp1kHuXq5KxjyA43Bw1NLJgY7iuQcPXpgTazIiWSIqMDKnjI
0wX/ljIGYwXbVfAljL9egh/2nj12Poynzsc0VSH6Nzb5IJpqtNWirJ7d+eE/lvg/
nRTKFg5xtCmvU9qWPVzHskPfbkWKqcRxuy0/gIlAhBG9Ad1QKvC0rQbeBifRjbdv
mUR1Ji0AeiFfJqtmnvJi+DI4ulYpMdM1waVBG7aof6in9U427mbUUHAgrd1SmO8L
6WtzY10Z3HnYrXD/EqCPizcd7Fej4r8q42EONyvV3iXLLE2abGwkAzPjKSwe0aGF
fkP3eh79hDFcnnj3k2gniPYOlxWo5m+KeK/bLwHy3eVInnQExVbThNRE1lMFqcQU
XEstg6asqRXYYS5EpmRyn9QAPTiaB9BDmXsVI+sdpxlb0D6ajeGk1M4Vm8UaM0HD
ariqzw2+HE159fox6POoHKmED6y/Nt5+Re9KQo3NCJx+Y0rADU2H2egqa6T16LLL
tcobxWJScxTzpQpQVoaCKfkPG/1jB8+DxPWGlLqEh9tDT84/jT08G3R5zvrkODxG
7v0ubRd+MtnGCO1cTu3ckj9FPFx24qDam7Fa56jewALxFnENG6ZVqD/oyin+V5ca
xAv4SAr5oRQgqGoKcnIddmgkbHBViZgHYeotEB/ug9d2WPleT9yToiheXxk3PPyP
l2TAieID00DJtmUTw4nFGpFVpQKQ3dceaRQmje6mcHxI1EiE+XbKO+N1czhrjoD1
7Kz0tZ9p3oDqAUrsWhCLVwbz2aG6IT3ClO2N85Ej24u17ZA3YBD0abcXK8GNuZ+I
xBBida3elGj/hheNnFp1AUTk7dbFRhUW9CMGRbqXCA7dzWlCcIx2fmkBV9D+yZFC
A8HdywnHoFbIrKDswBZOKI1nCi4utXezG11QfoTEXFG97vgjbjvaP65RiHmITS3l
LrSnE3EbXuODWtVtCc1zVUUFqPfARVC5xrwCbH1G7L8+qr8drsSe7MEVxNn4XLzT
JMFxYf467R0zJ6wzVvQbtYbLHO7D/Ppa5hHmf6GbqogWmXB92yXnnkd0XIfrk+3X
tyHqc7+4tic3gLm3dClEWKWixoLeWzcMWAEMiGOJIw2kaSv7nq+8sEspFbQxieQ8
wrhQ7C7qd+id3Ib7fCUklwInMQW1uK4wah5vMbmNZbOUlk3WK48YwAMFKVYLySe6
R9akGdrPTciV0somuvoCO6fbhOCXbKnIE1g6OTXUjaKIXi0xuvP+H6+Nh/wKThTl
1+RPawVAPMGUDeLGA1kR2RAo7mh17nj4L9Gb1TxDCn2uzjPODQxcpyLWt0/QmwsK
X9DGtLEYQG4xs7rIi4kvJ0LxRfQXGhcLDZlLcwYsAnDKJuXSQZ8cVRC1epQmu9WZ
ZEvmVTo1uLW5QeRjPfIuLKeom3oEFHioI0t0DBtOxhu3s+7GfYxre4eAS1rNUJBB
x3soSgT/M5od+fRMXaSIyMVDlzXuhmGHMwnRahp7XX8zeh4f3et2nZePHhoDT047
a3AhEi/5Gote4oEzPDXzP5m0JZ0/QslQMXBeluf/9n+HkmTsQYocMSVDnpD9LF+w
kXmBJKrE4RLQRu65aMU/kerFJfjF6mZcB8NmW0Hy87mOUI5Li8Bmcoclus/RKAlY
pniY/rcVHGKGnhc630SvGXBiQtossPWXD7s3ki1jOtrVUdB20U0Nz/6vcbRmf1L0
MkcBkawIr88r4WIBgXmHHtHOTpJmcW6upKWJBToN6R7/GoU9d03hc40xQgzfK4q7
oNMlkls8MiS0sbnO1g8URg8Qi35E0TPUAQi3civVUpwF7UkDcAZRZ4q8+oLLtWEi
blhvbUS404lreeH/Qd08I+LGHzLC8vG2AvRhUZHCUlNtvZgcoeqzQbWPb7Lg2kPX
yezkDjBInaO7LcByKjNAhtFb+Khl+6IgiYHoBG8zTxy5npZW8OQ/NXmIzpxosvlN
uCi5LHT5HA6Y1v+e8gGN7Tqc+RHCiJ9tyiTlOhXNgCXVFXoe+GkzYdwUyXJfJesL
l24AOg2v9jQuGvDA9XA8MXP8heoc56qj3BThKPszStNt5kGLfnYQLnZ8YTIOu1PM
ZPhs4hnodYKUvjpHHKpNBHoxlVnt6a2w5Ytb1fO3XRYM8+MeIU5QEGqkCo3m3qAk
FlLywTZ1e+SjMssumfWAe6oaWM5rqT9tPUaPcX/vfCYknU5qpwLi/foUHYpxjI9u
vfL0d4ylkLxEL5zJkNT2ZTiqsIdMUYZ2HuKfgs8NF4lIwMApDrXu61ZXpDH06yO2
Vce0oGClzMjNH3Civ8KLjvQT/6uTwV1/mJipvM/1MAi4MBw+c5UZASX3HiHmR9K2
wSANvTSU6MUSDhMs2g6/5IxUufJsKRvZlMbOAH+VM7TkT9wxgsKO7XFomCJzxSso
r8zkJ/aAzTpn9pIiWAKdOkvXBbA5E+hMivDkjW5NG0P4y9GQHQ1O84CyAt/zAWk5
/sVZfQ+vbm4qhl7oEpw4JpkCqESA6CfOQ3+QtI1Sa/mSoMLYo+OgJkbpM0Bs9zCb
781mkasf1rkvoZHE+0ssnWu+Cj2HTbTjJERK4qwCBKS2RNK1sVKl0ddtVnPsOiNT
9o3ahkO9/Z4dqmWRkTE2753eds23/iEqF44OaB4Mbwl9aSP93zj1vX9vsxI6/Ljm
AZAXt3L2zp2PvKPilwESqaPHP1thQGXayisDk66wWllRTUsZ7gA2E5WwynbI6fgu
Z2XSKqlwk68hGNKc2LXEKxrxtn8WSsQUIZcb/rXiLHSY5OF90YNoSdOKOw8XJ0NM
zMUzhowIqUrQPLuvaoEgymYyN6imyeHt2aaNKRMDDXTEtUINVIy/aF0RQ5DfR95M
41pM9i/kmgZ2jvzVaMFT98VhonIo3yibEGKIzOAsvtn4elpVY4s6G6qhfdmqIzSi
nlUNyVKvKDMagns5cHHNjJE0I0ZV+Q+1Dm3nYQynKPdD7Ue0q7ah6EJt5QEgw6kb
yE9V9hdz1YRL+3kvmPkgoOFDW9KTwXBRyWQ6++i8NZZVuZ16m8Z0VcY2u7rTb1Y9
cs6Ln7FP/h1+Kqo1ZY//g1npcGLAMPTjEVbP0ANVm9GRnw0T+nnwj1QSboboXC5c
RU2YdcDdfIbolyO+eLpJ+TaEZuEZb/M1vNejTzMtFCIMWBvKvSLoNDmk1D5soGr3
aGzDJjMjtMbo4r3DCq86ytRKNDBLp795/0cKFG8L1p2VpV7t9Cg7aXSiF/coRbBP
TJoApsHjv1dZBBNfxZ3JY7ZEHL5D2dPw+4jykNmHnoTgvsk0PrdghQ6ITcYCB5/b
RbRoxOi9r2L5rOq5hRLC2QB/nCGp4IpDAJhgaT7uXgqd9Gwbv/UkDWhEoGQqkE6a
baEEdAT1MdYCRrRIgQGpdBOZKCUzDjZY1E50Vkbs85rGsDu4YbhQgEPFrQR0+ZIt
QTii/mvOZo47TsgayGvt9DT0YPO7JlMrXD4GLyjlS6VDtj+wFJFlzJEQFwzD2NZ4
dG8Jz3DId9DvK2eBzrlhE1IZW6xzUsudCUVaXVPUvm2Zq+tSJQzhqdxRg53cIkwa
hqM7Bd29WFiwHpq7p4n+XFlYFlZcwiDRBDjbZP+N6iHR387P7ouHKlmRislt7Oyb
4+iPWDlAxWXhUtfLdjq8+usSoFXRWE/a6oowd2siX0VmF7RibNXHNWrj3ky4sKjZ
uUzjHVvGLYZoQ9VT6CvKV2g26w3PcGEjbEd/qBMtWMFwkpRypXrxZ4dTBTvPQOY4
y31DlmiTVjIxq1XRiekWVYr+vjbtSspwlIsI73DCiTeBgTWWshwTvsvq0GcfhNjc
6KZegvgvnYUbHVrwmBDDrf1RkImmY611QyhzB+FwGKPt9wQrxOYZGuC6sCfoDMlw
mSbwpiujBUmBgNVvhElW11uum52bB6U0c2aLqbp76G0gkHxrKqmsvgIx719aSXjD
0QPEYBI6ePlvcZEJa6JRhjATEe1CldphFWLy++EclUXBNmbQHa9Xgcqc5f3kA9Bm
4xr0joXgCU+ZXh7TF3TpFwxILaT/w9MD0zCh0jBKZIwjXvhSMyaXOorRtgIkqq+8
XB7ThQaosrl5xmOmCvg8/jRW3OMkbVXSsCt28wzOHpJ2b+8xI7XrVleYD5qSotg7
1Zr7b+0uv1qZw8eqg8FXGOeN0XsizFLEpuGyCXmuvUxBgiSNE3RrjE8kVUJ6+2uu
9MnSU0vvctbLNtQyOzR04Gtatn4zUVkjyRXgbpXpWtkWHd6XBBI1FWczXF/1TgBC
+j9mlUF1OHt4OKT/ArsoI3sdnQVNXmnvuR9S5l//uSItl3KPXgrdFXMomH59+a2r
E9hVdR9/NKW0FC/Y/1cgXQMDwFe+XwNeZxshBjtGlMPvNVrFaplWeFBb7O6Fh2wG
ZDWKZ21edRrlhTwYa8bz45JM1SUCSuwrx7PQtbAGYutSIlVc0q32PV4sXzA5KjUX
qAa7FV/wqgKnxLKDwiH0nKjaky77aWPi5FRCFHgz/bPlLLhB4ABg9sEeJiWJ7ALq
95orcGsiB3eOLANMapRIGnQHyiMYQ6x3wfVCcIhTS8C0g2pqs0RaoS/fDYC7pXQ9
DCQr8MNMrbVpdd2Lpa9wo4WVzBDMloNxBZQAeVC0fug/a5WLHWBsycp8+WqBwRm6
TmU2J6VZnRVs+3S/UidnvCucB7/QuVOsr6K11jh2pLozgxlz6H2urdKWXHE9AVgZ
L293hAhEaojQZyBmnUks+0cT3itgQGsb3Is0eGqtuA4S6XrLXDN9lusgeqRK6Dy2
0nCodchY5N/JdZ0WT4Q3lCkH0Ty4ng+thVRZUK+kij6Po/EzbaCYRd+TVvRt9lr9
22nC6ebOfwuXW9FC4dV5bw8K1CDnKjbhOQoKHyN7Wje+d0ESTXWoxti5vkzDlqJ7
KauUTHbXv5M9hGcC8vO/hQqjEykXYxF6Au0jX+oWMu2NW8lM19KXvAlyxwGkCV2u
a2VsLwgiPziqHuxHLCYE1y7WUHoqWWOeqFVzC0iYhWl0zvFTxISflnwi3fSYLO9D
Y0FhkryjQZKmsPL2uSQIEWv4AE4Ti+hhVEjAzI4E4fX8ka9Mb3oowH65wjMPrrzg
4hITvX6bV8a1d+FEpn/l5CLqYX/SxFgscfRA6Ys6AGtqBW+FyULtiJGcgDyI6NlX
X0rqvpONHj9wD1zyoIJBUq1Uc4vyoQ79sclKW5hdSt98D5THq+5++NQGUNgPcC9D
j0sdz/BI9jy2Cwt+ZRia1oQS1a7qV/Zex5+WGdT80bB9FZVxZgZMFgggglWbOWq/
qp5imJSxxCrRAWdMJCnbYUU9Qzq/KxbFgnATIKzRfX9r2zNozeBU3lZy5yqnMPtz
1Zbkw9o2qq50jVhRrCRNc9IKZPdnKWU2F3cMQSghVHvd8OuJwqgT4pEKBm4RZgxK
qypYjyiIDXPjQJ4TD9moKeESIjNVQ71rQHR13kbGR0YStbE6j1J0vMCjQo1jPsfu
dc92pvxtMsL7/9M9dLDu+iovKdLz48SWEVHzLODJ8PUEo32yXkhPBvzuvyqWr2V+
sBr1fDQRtbgE654lqjE8rlq8j07Cm40TpGX8+S9Wz3IUxlUWY74VBgMwdwRPxGH/
imMYu29Jqx5Tz9GKSyZP2xdDd6INyfMCuVvMdmxPHq5QbFTkfFxhZaxgPuS+eqQp
ZbkiC0RF6DcYluGFx/laDYMB5Ts7ma+paBtdsTeN8TW7SfMWJBxdxb4vUxWIfDSy
R3LL5b6REFKy8ETh6/HKXoomMBwlxBvctHZcgYHt/wzvbVfwDo6jdxvZ6sukDFIF
fWOmXdvhXjK+qMluMTMCXb9kfc3iJw+hChG56Guol778XFwqCGlk9XnE1yA7LMHw
SExugHXlmlX9k5TBqofdscmjPcDjxw/u0nVGq6ssllw3jGqwUzYsbLLB36eT97t+
b6NF6CNCCRUoIy6OyFnQTU/KmIfnsHAV62dJ+jPSSL0xpm4YkeFVaZHH2gOYGV7B
LxGvNqc+/j7yqKLfsB0SM+ulTH4a1MjdV7JMVqHZ7ne3ReEnLii0iUEoAvd3BNyq
l0ngVWelfqZ/hsYyMycgqSu+gVRV6h93q1YBXIlCWQ2RHFsecKTh8yck31kL/5J+
NBYvhK1zmeTDEJp9gL8tkCTGDjIM3zBvHnrwy0xmijydNZsukG9mdB6a41BV2lc1
Q8nEP4qqJi1bTLc+cdJyc6PgV0vlEcLpLb8pLrUPrpQ8tQPKbvE2V4FUyGFgb1AH
dnrdUG/dVOh5pD5iQgqs381nIcuEeeBICqZa9fML8G6HqoIaNJGZE6RBrTTIU9yS
Ymd8AsUgrDGck04QqTVM6wve3ShzqxU6ipLBhccZYsc29gwHLIVM/m8HHGoYBw+y
QDJFg7I+1y73be0D2gyJu5NbbTYh6SZsCcUZR/S50dghpL9ZGF7tIo8BDXa60M7f
pLMllldK1QI5cDdLz2OCv1ONkO8Io/NS0hVPIsFDeERQ+SzBH3KiDPcPt84iDLHK
mMrm3w904etuK/YxWmExaNcbhDUUVgY2i8UVEB2sqRTAXwRlX9TDjUTWVTGjvPR2
Yfs36eKx3QkNpNknRDXp++D5EUM/Jctu+7avdpxDSlLj6C/ukoDqEdDckLIdbChO
Qbu+yvQzC5nuS+98ey40UF4J/opCwPEqF63wP6PgAZjUM5Sj98XQ2VwdcVly0IAY
uKosIOuo1Nlspstmu+YJttUV1z3XY6RAh6gKfpGNgtWU92s5k89b9nxDx3zUkF9F
NeH3Wzn6zXRO+IH/SrmjPVwCFzRbijmTPTsBfOe8vcZ74tluWsDh8Tirx5Y63AZS
zjBvjMux+mLKApK1gAL11FDSj1W4Ze9uYVLMV030Ocm6f3CxZe8n1xdf+1U0vp9L
cEEnJ+D/c2Au6ytYTmwmR7lH/liRXqAC3rGXvkTR+0rj5NksFYJBYH9oTkULGE/x
bDXZdZ4z15eNGWL/zKtVmbL20Vj0LL7yrvL5+PckOyTclEWSnQ/O8KI2LPnB4AZq
A/++uv6rQuOumntUhpwvPWVI/VJH0uue+CC8c1wJ3+skcpYZVNWzWkmBh4ecNbT9
W5nverDemLrgVdqWKwVJQK/illF/qCaUyX1QFWqros45y/DWyjgq2VsxOTWRzJMv
FQJ5qWrTNv+EXG2aFqE2oTb3IQtm0RKPzA2osEh3A+QfGPaHUrGxVrz7IVJ0wLMj
UnyRh/A+ounMQaY5jA5JYkAr/s9JiW3DWMrTn94kX8fXV5zwalJ0FxgNiYMEqEzw
6USG3nEv/wejiv6Q+wPfjysxaLS9p50d7CCnr+3ldvfI+xrkQTx78cSPjG69QJAK
YdmMu/ieIi2ANvxskm1t8wnmGsQmgoctLU6o1jTwc8ngI06oSRSilefUT5D1abCp
lrRWbwDGkuj8jppoMfW/BoSa1zAuBPIqH3RCIvGn4/mARxjAynmYkiKW8m2Vf02a
/gVbFpVHTdmIGgfoyLztn8RKqeGhVJc6dPcN68oKqRwc5RyqVfYxAJV+rmMKnFW3
hR4oZPLAADkCyBAF/XLI3LIwvHaZfnd1XfWJ3tgcHLciJDTUEcMZEEL/SDrWxFFX
QMsqA3NhcpGrYsDrM9RvyiIG6cholThDPJzl10UWUjfrPZ0PuWgfMkxa0iG7jSFj
BhrnIwQm3B9yZg4rkw08KihVTW+UiuyCwvzFaOvYy5IB92bKvtqiH+QbNdmDKZfx
XXu3KQtRliCZkBFEaKFS0tIsV2+8MeBE7BeYHX/In9UiGSSa5cy6ZA4WhB+fq5+e
zEl7OIDqV5fpJhhHZRX1Vh/oCiQI28pAq4udDJI/xLOFcBNauHE7FCCBPLYmE+7L
+C31bT5PY0E5Il4qsTXijK/8eOGXKaHGDyACF1WWGnPHZkgroC3vy3ph8scv9irg
me3RDv/L977RIKw/P7I47jFLZU9ayINErHTHaVp/zksZy0HMSBYWQ7t5Pwv9U4B3
RmcgufQtJsih4WUymyW5zHEfwytOojgdL4fenRo9MVwtyeg/vsZ0veU4L5TpJwpm
IIrUbhs0FOfdXRQzyMsJnEu7aoH2gu571GvIDP+xwfiTb32d2N58UIIBLtc+SUkq
STrhDWPa8Bs4LYNfIcWffC3vIpsXks+prLMgQohZK042q9RVxedhNtjJKgN4MwqW
9JqSMxyivsmpYjS7v5MnWkWke1QfLXJtG9CZQw8Lzt5cdiXReDPFkgKlDlPUVH1l
6jC6Gjgv+Bn9/v0cuNhEZE1Nvzt7BFAVGMhzSI/Oh38FizbeBNLDYbXRrfO/hnJg
dbIi7D/HbiVwnWZxDdDyJ45bQ2hXvhizVWaZmh0CKrFGJk8GsFESaHTltt6kTqAl
UZjFotVdRPS4iobeJu/3aurga0VTCJWFhMTVzio1QZFaYocV57Htg9ov39ZwWi8U
ixlC9F28qyCe3T6eeGFckKOVgFLtWr9TmdFoUjTE8RoufXeslA0nLhyAPO09da6e
D3XbL10i31JigoQdzbZGw8DewqheaIoVwJCY2h+MNnsDVJNBeYhyLd2sP5IhxZq4
vYaU3HqwlBW6XTSb0eKwVAVWcj59vr95ZjDuVyvhcE524hFW8n2h/MlLaixH3QY5
FWsDX71LVMYaoRnAe439mSIdSmoA+So5ngpiVtzL6YRTcU+c1N7gL/O8n9Zjj+0B
kYY5zIv06T23pJyeLsDX6gOp8uldniV6wK9H3Ee+HD90YbjCYjgEi4YdAtuhyMBH
wRp5bVYvNX6rigwHsUfoEekwHe9h6+OdCaHO6EfBjjRb1eLxeZtQx6ih+4k7GCSk
oDaAzaPkIJSQP7GKs8GGgBkKJouMtSFRIlBf4709Bq4deOkbmKFRrpufaQGEhDDl
VoMkbq9sWU5Hz8v6eMGTOjDQnk+YRJ8R12uI1XDuh+UB3csSLYVl2AGYfAKjBuK7
Xty2K4cbGncrOTUC2xMSzdC+ryosfymBHcSINLjMonJT09WIcIsvL8PQyZzs6yhZ
WMILQuknb1+6oPvn9cGZ4pkjVXiDHGDWJbcFrAwWCN8qdblgm3iZo4OC0bS9u0bN
l74YiUIryG3REaVz0oNcqnKkuU31/8LM4TMSmZyItYxKNNNMepTSy5uVpbPgEU/v
7eyzLplVbseSTFUcdRokPzBU8xFEoKzY4yjPgfzFgJ+nXWQoAeyJ2UoTkpbdebaV
/mdoK2YhnrYkAlLDba3EDShmd5WBnbEvS+AEgzu9EyrZ/SHxW3VJ+933l1XhxEJr
evY8r7Kx6gdzPRzhV9CsyrtCIB6iNWJmqmV9xIfdNlo9R9smSsFsO0gK8mUuqCld
VqlHAKs+WUAjM4uR/dDchX0YKxk84bv/dyO7ewCUy8uzq6aS+tu3LujtfKjhLvXl
FLHPYE/8oS5a89AVKCEPwyFubG3704G8Tm5f0WXUGUT7nu0uRh5lxy0Gsi7d+DWI
nVeFlRS6AVXDsztorjavkJd0mTRuQdFvRjVGdXCs0LRvG3sodvkWoR1TpD8S31Cl
qG5DmDPQB24cy3w5oGWERlGPnHRtg1KTqoCzI6ErZVwFsSnlai5DykW1Fx4DURVB
cJ1rPbXGkmQP3zRimFiejVJjJ6v4D+juaNSLbvUZ2Y7HH9lVwAxqs+aVB0HWzZDM
JhGd4tuNWj950Cr63zj8lmrHV4s2RB0pSJw3nVXDmkwjaLRUsiM85jaUzEmTV2jg
fItrSN7wii1A57Tmb3KoPz1zpaCOVdMWx+v+RGMXqyhLIR2BX5GpPaG5QUh8MACa
lN35YMW3off4+Nn5KBHf6USJTuBN7tGxJaK7tOfkiaW12nm66IghF5xyDKzo4yQJ
E0on9xfBDP9Hux5rQiLgG0Sqcob8C/awyXc8B2gwOyXhamZNm9b6QlWN+u878DEX
16UWelAMabmN72XEtu0geeEzVLVR7WtSDGJtsSMpb1lYUBpo4s/vFdCeRp1Z4/AH
eNB2DS1LJg+PPtqDxVoTBMjUiVRTh/DwazTY/ck7f3OlgdgO7fv4iCeA8KWWKMPb
fZqTDj56kEtonGfnFrhRUGaHFtEP9HVaPvZ1jxIQ7/J99uIgCafBSVxCKG3KyL/e
8sABg0A68F2tMdkiam+EgH664Xj9rZnNrbVwncz7YrGzeHv8Eg5xCjXOFHjrgstT
hZDNdmdy83PnX9k2dpTcMOCtQsyk2XiMmAquTcqp4T/wjfNuD+3nM3m5N1ifBt3u
yb+ZIzg0qwiyVU5FLiX6dlidKll3Ad5YVJpqjUt65XeAalT+Toeyhgpt7ns8sfOx
7sa/D8qSmyLcjAHWUDd2aUZMnxLBKtd6HLaTyYoffJnBaf/Pnl8LgX7y9UOkkZqA
htjH8tg5UeKJk5IEBdk41Ukvjb4ceg8wpty5rcWnvb57Svf9smhqB0tS3GXBmknN
ZqiA3IOUxX2SwVrUAvpgO5luWsAJioNr+LiT6VCyCixXNNAvWfArg+KA0lKi1ZMH
0DCmlqc4RtiyAImCGouWAblGHc1RsCNDzlLV0rfLAVFvuEe7F2fXf4Schi9W5d3Y
x7yA+z9l7I5buv2JAIy7TON0Vb7XPGnfLUMd4meJm6YEv8vVoe0Byw63KpPGH3C8
YpW7uOOeS6cZGa6R+ofQqRfuWgje7M+1zIqBcSth3EcXZ8wH1Nz9GvPH/3JznFr3
wpeym45lrHdv/8TbP71KH/lxXmXh6Czr4N+gFwZMyJ374AqWyHKx2VZJvZeJFXXs
H1P8cq4ZVjZ5sIECrh0pDqfBhse/KZ8sF4ApbgjF3j1mX6N2IVLTstoB9qvdqpQc
naeOYLzDh6nnSzfEpmpOtAN9iEyWez4FXxj1RsB4M0fLtqVqhb4GG/jKlazhU0xr
cEMrBqG8PYFOGYmgBrqpJfn51avjgfBnqFKwg2z4W1yN5fuXuOIstnp7Gdsrwh2t
vMyfnzCmQpxmnfLbNl4eNj8RRVhuJqYwxTQpbRRrOovcSWw1do0fW1MFusvf/dMj
ATGU19768cZQcovswdCEsSzUMMaop+i+F2FUFqyz27lPXLAoIV0m35NYbl6Zx2x9
1m9O4W/iiM4/H8M50suyHJ3kMtyeOjz5b6Wm/FRrySWSUQt/K8jBzY8d1/uelAH7
q8COPTQ38TjiEVszzTQRMsra9lIGtBQzUjtM7AiEwofSGW4ChzKallChDgpOj6Ew
r9Td3tAzoOx1R4RIvcxgjmPAgA1qMbXFG/myiYwTmmAcnlJWetmrQ9ST6rfTcZOh
iIwIgXCJl6KkleiR1s90l0hmp/KBiauXlXiXLTLwfuzQQ0kCO1VHOVOsHKwxK+cc
8GnNVecWNVMEffeszL55dFI3ILELHLN7W8pJGyC4Z9rugWy0S70GL2xdleVc/mIq
NcpvlwONi6pG9yYBLjIjIOY47xWCvTYfWVBhJOeMIhM0lmsSlIcj7RwdiGuyl8bk
Bd5uQM9szsxawQUPh42ZoPktK8qs6gpSa19cz4LygvQQCkALh1Ay8wfAqXlljW/e
VA7tXbn2IIlFD3GqoCoCUMpP3dJhIHxOtiTqBWQ1899bp7vQaGRPkYCKiA//XgvW
tMRUypfkbgIk3/2v4CW4Ns6BTTvIlZhW8ZwTeMpFm85ZSb9RN6WLhlzioXZevjY2
DLyggBErczfFT0piCBJOTAaEd3klVzwL8QI03GIy/uddz5DNktikGG0M50c7hqJf
JrYg4DsPgSEU2oBeFM1qi/RORSHqD35KfCafDSQiZZ1WhqZlgvblEWOgKPX4D3RA
mQq7ehKNrUb/5mLls7PN70n+gO+wfzsAjRzjiT1ihZuAe9C2M2zOgJWNCeaW/EFD
aay9ZEe9Gx8+qO/hdsiLAU+Z1ipt49AloxdKIj1V8LXN/kiWJ+mJjUO88BIcqa2e
lRN42kM4iBeRIxvnB7cnwzeOuIG8d/mqXYXDTeF+P1+Xzqxcgo0XHd9hDAagLU3S
rSrLIG1eBuNMQbZo/YUb4UzqCWXQQ9rDbntm/dTkaOH90u/VsLjkT3Yd8nU7tCQx
HYAHro+0B4mB1Tk506HKNEdg/5W2PfewqgziqFQjp+POCiiUdmg3kJ4aNRSBAWs+
Oq8L/zPl4VYgmGUo9Nv73x7t7Nj7178UEkeBczFIW6EFd45BEXpzOD0fEWezrE18
QFa5WkTGV3+Ym5Qc7mhyYcAvHO9yspExq322tfzaY3/BRq3WZqB0J08usq/ppWLj
AumvOnRFifwms3frB+b73RPNaihfpII9wGfQv0pmqnRLNmylCxA43yp8WfeBxNEm
YNovCAisiuQhJ4ZO8SAl/DsLCY7w5u/Rn/lj8K+4wVOhWq7VV7W+lwICkAP+aRko
sG8O0XZbkSEYDkEeV3stH8KCRGVzskHJ2ee9nJAS+UrDX5Pd69Oewd2lOTB4F/E6
9Udb5nUb0z6esnLnQak644IMUQxYRss9MrKESmtEtrJWwTvoUXFyws6QjxK3+U8/
3L75kmcCk7XCMsKGhRBCLyuu9hmhkWwsq8ue6+tjAq3BF/nvSF/nl5Nd7I4O+EK4
UzqSoZCe2ITaWs0Cfeob8bQk+x6z89kvstgm7gFwHuqd6+m8dB4lNxkXAN7cYRQs
+W0Rlfn2teMxp/7GOcWNpQQfxCOH7nL0w/FQhrbUsy29GTjM7AZBPFcU/a3qiD+Z
hqPZfeqJG8ArabBtCJANa8melOyeGYCj/rJ1BH/2TXKcjSlvON+7z5DPGK/GatjH
iW7UTpHGtters7njhaU22qF+DQQ1ymvJnipw0CpTNX8VaGetxAIUrLTUP5FhHVO2
RODb8AG25ZzLP02TfuEsfrwoaxcn9zT/n0/n5N4ejA07Jj0iQb/OQ/C6ibwZfrRW
TZXYIg1j0PG+Qjd7q0wHVUc5UDOCZSoPgJTWKxo4XRnw8DAyaUuScRDoiiaXrChS
VK9hfTPPP/sYjztt7UizR/WI5bcfPEi4lr/x5wJnIFsiiPmdSskAPHfgpwNFF7Pt
jqrMDQmUEnPtSZcUjBzh0m37O8LQbrs2x3s0deJwi1PXG/WwSohbNNASYsyR5aSk
NkrxQ6ywNhiX8do7H+Ol5EFUZnRkId4Mc168uvIT/HV1WxetL6tNTDbyZi+1a+hc
JPIpluHW0eCDl6Fv6XhOo5XbW/AW3EHPAYTfsQnOTrd4I+Rwq+1cqrjx+4WAru7x
LWn0j7GtZjQH57POm0+emrb6uBYb7z8bSjn+901sUrc+Q45iNV87Va3cs7dPZWR7
u2V5nJqj2rTwVSqa+7dc6DZXjS8OX7DAErTJYtkgW9k7yAsMtJNjnFUnRMtUAQNS
ulXr5x5aQKCT84FKQnm0kp5BU151zrbsoYNmg7SvZeVUwfwx+9NUyk62oDloKQLz
UEP2kR00/fov/45ztidHxC14eRvMeuE8t3itR4vZRBAPvqiILYB++I0FC5r3OAEY
s+DgkyX/sHRwqBgL9ryNwBFGYmU8jEfpJ7M5TP47ADBIXv0oUHwUlP49AWl0Ontp
LBtm6qAd3tp0y0+HQyPKw8/wuUye3Hzzw4g7RQguP6ppDMFfk9VjIp0yS1q4YsBY
CNi+lcerGihv+2+8pXnowYKwpOOF6H7e296Ubd/tykG6TkpxnZxKPoVxLEsrxLYo
Ujhc3/hNtrzEOKU4BIDbnXX2zpoaZYDs9KIiJlX+PGkYdcZN63BASfdKPfNuR2L8
Es1G2p12MNSEcizYg6vMoXWZcowmosBSzkewOm5yM8lKJjMvj78r+8u8zB2R/fMm
RP8g7GME/2fv9PT2ZAGSL3HASEZi2158fgFRJehjJtrCVtICZ2A0I9tFu3VErfPW
V6eBFJuP8n0n5HKwtVuIlJS5G75mbqtaJYS4CoqDXXiqz5n8pCPIi/mxF4Sd35WV
+RrZpyzJOyLXAv491sIR32zFi/Orl3grZ6XqeZIb9NdSk7J5+raaqhdsx9Sq+0xj
M7vBDGD4Zre+qBRXCka+WyxtG0h2LGUxl5oHOnvpUBXhen+OiaM2aemfZHwYuURY
j/+YDK7pd2ZP+VAinpKFJGJZdPE5GCa3cshXMwYulkY8/hpY2kFwpQukp+jE+SR3
cDKdDhI/XPo7Ph7JEnLtCLqXGEufv0SbexAN1gJfvW3odGOLodqXAAcNSV+IsJNA
IYb1b9YKYH/uKOMhnikmrlI/yXAnM8nmqQ+OogL7UVf7+QLwnAvzTvnU4xj7Cuwz
XpHqpQwamAHjY2NFg/ftFsAaZfyuhdETsoWPkHElgxSeDECJhz1vvehiozjLCrgP
ig/oPikAqh77r1TWLgpp3Fhv1c9LgX9Up7u3lbkg4AUZLXT8bF64BurPuvTpa8AE
SYS4PTUdUxgYien8vxiYpTIvsie9YfbECd6e6IclmW44wSF34MkYlgDoXKUldCZb
hAEzKAYo2/n5rIINYA3QRDwV+tN47J6kPvegoT6VjNA4qcC+vYu/T9HdZ78wKMb3
CwCcDoL4ANDEyjjxDYYxNWcNiuF423lFP4nVueT7B8pyOE7YFch1ykM+geMDKYMe
PU/yTvus87CUdH9gt2ClvovKain7XVz19Prm55++pEYqFl8MBa4hTCJgAwBTkZYB
SAIUK4/KsZnUqslIp9QVy3PcjbBnjXWYmmQigWf2J1QIEhmkZ5wX0D7f2/rsWRoQ
`protect END_PROTECTED
