`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UtGoWkjdhre/cP8KOlUNPBc9TwOoDyB4Ggd8MDdU6eG2Tah91eIuRslDKNnMAejF
nXw/E2GjhV/8GhOsxYFDAZtBldxYtjS+0/tPPJyEXrUJkICxGQshfNa07w+Wdulj
uazJIkqFogUORnfVk38BVNqSgX0PuC2oIOg1zATNFOWwrDTUBDdC0V7Mch/f0biW
S0CMOD8PJluwd3krbDkwyIqvMdmPgYA7ZMuIPfz2typl5/zegkmvePEF+EDrcu6Z
0ZFHmhZJW6vi50fmyivpc0g9+f5ZlcVHZsppfhC0TtMxSSMvL+5Wm6c776VivngK
bV6bkoBKlo9ORQGfsBQ27rpCTkSWCRAW+pHH0AI96oOokkNkZMWopj4wRHS//vyP
u+9FN6z2cvVG29vyVdcBXtsLpnACfvu7WcqrKGZETc1wODmfeuwhX/5ckrmonlyX
1GpqPJVn92S+PVlcGy5rKBwm59W7rybQWmTCauOlhi8MiEsKGKny1+APs6+laMur
bVzZgw9eTeG6lBRN9OdOrv0trSZ8mhhGHlVqdB/0t4CHGIbFRmV9xUw1UXgFxVDq
FfkZRgF6VkoPAGPj1+axviQIHEnxhGH3+Fvf3a3bYMbQsN/R7SJ6bOgiliHSaUgl
s90VYT7PLte4Cg1neWcKbZz/CfnDD3fy/s/E4Prk1ZpneAMxmvnHi0FN0cIp4+j8
Q7bbOzZCIM74A/Q7bOSsWEBEMJmw5BHEb7z3sVkB+Iq2QknuKHEN+Hdkz0w1dKxf
qqvrin+xph/9BlRvpMsGU+1nYhB1XPLiIrzs5omVcJoqSiCTIUPpkAQ8IXnoi0AV
bE22lJJRiYyqenGf/3imD8CP9sNAwp11XpX2PyjoVpY=
`protect END_PROTECTED
