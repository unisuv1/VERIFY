`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pWxXXm8kmZIe+1rfCK5bBxy0CF2Uu4bPLN0EyijhYqwhUnHWbNwSXHJoi7yM25wM
WGGGaB+XX1N+utLtb7rHC6pyDp9uA29bCONenrLaEly4g3E+xm59HKkQraQmTih5
dgocJNqMEq2lbQZF1U4KXofdK/4MPXE1Kmuj2hVru+o7wAPGs10611AU08VaHsmu
EvDH4BQSt1Vh+0mrURH7xbDYqebBMG0jVIMScF246tUtkM33cMoj7bIu3vYPYuPi
1mrLG/x0XDiRqYnAOg4jnVD9+I2mmkiARv5eUiysZfucMu44KOO4AhBCifd0qiVr
4CCkNXm4jhk0h7Xgk366A/UWvhsb2TFh3srkiBtlgaF+OZtURdmUUKaDjNpYVPEc
vKuU2qmTJfc3W6YMpCSksze4myUjdZdgE2qpWxIrYk8ftWaK1fCv/0mAb5y5JHor
`protect END_PROTECTED
