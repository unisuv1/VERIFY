`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IyRD2Sl6RxRmK/PGeeuQrusXseOt4S7cW3VuhDcxTNXLvdO/D/zcF26lPq3D6v0O
tCMY03rgrw9sU3Uf7S0VkTUJph16Pf5bkIbPgHB7m30I2+BCWlx9EaohcEYJOtsV
OazzvK9Ox8DSVF0Zysmw2qP0jXfeEOJ4uFQ/lly4Yw6h0Y4mh9ILL+nD7+R6LwL7
`protect END_PROTECTED
