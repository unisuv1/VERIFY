`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4fuz+LfACswIgPgDLDpzX1urJ6HUOxKDkcsBqnCby3z8NVPfVuXEmHQc46WCaMXI
R48dIEYPfH/wxlAbz+PZ8mT0PCp0Cb9PPh/1MT6JIPhi09oL4GI+0VHLyRLrZ9/B
Q8E4yOG5ECf1fFCcs0fa2bMgz9z04ysdk7vezgVQGvyz3DgMCz3RuqAHjzCywsgl
j3Cj2O/28zQFKGbN82WRQiIZ3FPFNKJ/flLJdjtLWkIZMn67ar0tCn6ESWAZYVny
0+xus3bE/TsnS3UtKrFmdA97cNm/taKve44o7NW3B0S6a2NGaeBBfNbsdWA+uEtd
Mlcs4YceZyYTA2A+9d1B7JawH50DFZ9ds0w+/1ROxPrTS8H73jhmCGqEApf12HJZ
q9HPIJbOVGdf+GDp7Oh6KvaQMtbuW6xhK1zR54tOIwOPclRQenrjgA3lG2rdn0Zy
353o6Qb4+36EoAjRyu5WkgwU6cXRO4i2tyFnoKpiUXDCq1PsEH0ACTjQRWkLc/Q1
f+yh7iB2TDOeOREfmsDKimzFKA7k5F9kb6tIXX3qsFPC3W1xnNFNfCW7NQC52h46
P/6OiJpcvFWA6og+SLFTBScrLS2z/TSIdJryvPKeEbwL5oOpxtRzbQ7NyOuxpYVm
1tqPYRArW/VC6LfRqSALRNBXIQKh/AIsuayhwLOH9A/kgLYUm/GWcsN1TX0UWKoT
Z4KCGE7JVTdLfbdHhIq854rAaIu8NtdfhpnOasUKtN7buMRBO9G5BaoZXcX2hEPW
2qNg3AjsSsYsSVBLeZ7mSLcFX5WgUc4qywSTJ5nzGSc44/Ayx0Duxq6EEYO1m52K
9WZnt4LCW15/CKmsKzf5k0+2UMhTeS3C0gHDm7oHbLdudh9IMCJL1ZS4ItBDuc7p
lX28UztXrdnI4uC32RorScmmoIx61DIpOt80F0u/4QQ/97p26tOk/AwS568QJC/C
wgvDNSNbctPsX6vbXW+oXaUsnlnG7EEoZxj9x0NayUAOHCyfSSUHK+D6MN5qJAWj
nmvseSPbw7xy4hJwEwF8A0+DTCc3cQ2fWbKhdHMkrEmZI6txjmm+eFaJpHhubREu
ki2JZe2kI2dG+hSJpp2RV5wvKEA4/q+RAAUK6FFnMZAnW+OzjuUmwC/NRZOwynsV
wxEkoHRr61EerFLuvyrvhgNuhN9IY7AXZtB+h6ei+Brtsgx801fxJFcVn/5EKaFw
XlKUuXRGVxJFHvWWdXUg0zOHyGI9pDHYgynk2mls7mxCzzH94aYwXbKwE7IqBh+q
+SbwGLZW2CKZ4whk8Bj6HIk7z/NClQywZmiCLRkbMS3E3tHSQBwCzEmkSi/twdbs
u8VDhEEbaQ3OAHC+YtE1BRpdVaXHgg6aCpxIxOP2dCZR2dKDvN0CCoqh+3bbgR7R
E9VqJrfFNtuW08jcVGmxRIwS4bs+96UWUQod2Ftmq9Slgy8XQQ/R2NDZBGxNXYqC
V6CpRujHkXV484mqhaSXTv8h+kjQilI1kdtjwtk5KS3PPIs24ITKzjj3lGHk+q4K
QI41t2c5I3k3y8lAwD3waorPFN0R6oKd4mAwi8Mut+gsv5qrZRqxPfiNuBOiI5jB
/c4X8vn5KsB9aE4mV1fUfFzJbRQoHH4lPeEATpPOgvhOzTUfKbC3BbaQu6+KNOdw
Z1KcFWCN3Vx9XYssfV5D7HEL1mn+dofdJMmQG2uePxjSUHjw5XtHssQyUrAtNuRz
ugoGxQHz4EEMJUKSsvpvunDY9bEgY/V+h1xpD066G+wTfC6OtGzqWZYB7JG3zhVk
AKEH87Um8WvTKFAWcWCMMBfaO+YRqaoeHNF6OHqlGzNXTQ1ixr+0rzLDFWEP/XaO
5PYOuDHMfrOPosWg5EJG5pZ1SHhdVyOkHIptStXhmRvMcAhDMHaKGOiOHXxvZa4w
DntEbZUM+gueVRDakRGOEEgrM5lIwmlJgnlPiSpp0RkqJBaDs6I3VzEvAfhHtMk+
sP4lBh6CW4ER2HHjEPIjY1oWL0hakSYFVJ6m/A8bLGWvd7x8XGhZd4xitONz5MLB
hMnlac2t+4gOGORSCTSTxu82gCj9yTS/876c7PLp3js48EnTMOuenxJppWYnHtKB
2Gw/P0cK3caS6zNWgQQGRpVLfwwssGmwE07OX2y8dKG5BKOHd0IcLBwBbVNvKMDX
YZJCOmLOPD9h/4RWE4er6pVwYo3mT4TcP499K6ZTqkBS2l55Gg5X1SbSCJWu9gyL
KGBPKCydrOmRCXtCndGkbt2YIvEyFoaLJqyNVaBCEbKyhDwWTj58hrXZWlVyHhkQ
XppEOs7PBjyqkWufrB5cRKpzsavvaU1+T1NZHT+koLG6pnqb5XU7j737JO0hSxmu
1Gpjj4pnU2HVIuRwcgSH6UtI2nRydPsWmzHqbq/AbIuipwWuaB8fTZxHOSjmP+13
sZ5jwxg/tKb98fTgILTXfxwBhHltggotABsrXgz1ucHOPmUFcajlrTcPJraQ5FD4
ccj97lamrmnOI5upZT2YfPqAnOQQg+kr1IT2UH4p2dEeEZ2sK891m4edzEtw1SI3
sSrvGm/jqssnnJwzD3bPEnPl+7eQfsNw3PFn/SeJCfDU4Y7aKs3Qmy25l4D7FTvi
2JwXHL+vWNHA5jLlfQQ4hx4ZY5C1Qtse2L23WstwGMFOA1FJ7BA3HSW/mEOZuO2a
6XARA4gVsTD3giLPZ0LtyjSeU0DEoQ/Tp1QjnckrEhnDb84FiViMp4wry/7Z8gVV
/anYPnrb4ZFC0QUXloMTBsWhLqOZiZhsrTa9NkSVw+V2AwG6y1NOyuESHYYH8oS0
20ytd3sGcRIR/roaSefiFACfvs/7j4GNYz9lrwqOVd+xnaEBVd78wpXqn4sNTFDf
f+P1obxqP7tWn0UPmLMoNpLstUFx0XxW1qlqOCzYCpK+gJlY82qk9z7tSKGo6BML
FdXbRx9vsPU648P7YbvIx/bz2dP0IGhp9Tc1Bn/3ZH2BsLhXL4krkt/XDkG4tx3s
7IuSG31kU4nWc51VdkeCY1G7DYUz/wF4MKSy3JjcCzX3AfSC4BngE7nSMs98QLBW
ZaNnK101Jk3GvXn0Xk6tTmRhB0Fnp6btw67/Aezg+Rsaz6FSlMIDrTDzdasjXg3v
cQmVWcXHIKCWqdLePs6QUOSGT9CQMbYrmDA2KJ3ZPJJaXK7c/1a9NVZk4Q4eh0+J
PRVKN6T3YwmBKKg/0JSvIcFEVAHYcRtuLo6+A5M2vR+YmZtjeOelPJouz0j8tuV3
4ClgnWOCTJn9O86KpVRSn7uGauoHONiupSAEOV/TNks6WxpfQl7MRcGP+/QyY5fF
GBMPCEmYbZyAdkEWGKbZ4pzDSlObWQMsb7S/HIBpmeUomwZYe9Dp0dDp9e1nJQeZ
2mZ1hk3RDBVQ08O6UyWlOZvBSYT9tAxUSaVkCFtW4uOte6ppoaub3jhuL4NELoaL
eq9xXbKJ7YFs3UkFdM+a5xyiHE1qVsQqZhTu9qdmz9cw7Kjwn7k6CTMH6Bav6N2S
KDuc7WiBRVGkq7v8bEWRK8CB+G5OabcMlX3LfficecRFc+kYxBkBSFtWeqEBvNtG
kl4358LEyMtwDYHFgAY9P+k+tsSQHFEoQQhvnF8oXlf7H7KGyLqVsJE7TeK4Z8W1
NHGK8K+2UAK4bdAxAggYB4rmW5uugdHDvU1SjzwFMbXAF17MgWYMAEylT5EP1BSO
0s1YEtkI3EpQWJyHSk/hRt2ccwW0OuyI2Gc4rs8SulmTW3qR3gHClWQAwLWidlgB
PM/GSElR6CdziJLb+a5zN2QDK85DFGC7yLw5+enh63r37CGmOQ/cJtjyFYs0oR2t
y6UvOgH1WKkqF/qCRPMKhZqMjmzMhiDMDcUVxV7Bl3eldJbs891GN8xY9W0z0D0t
7gSP2bJZ4JLhiyf6gEdyxxpRp6m2+gYx+iLRYrwDMydYWgJReqlCbl1ZWWxFLOZX
vfB4eXfx4fYh7+hcWJ/qFMGfprVCA6/t+xLtfdvk9ggrIz8n/+Uissr8pDb7makP
/pwkEvDOSguNvPL47Tw7BTrVbRzv9iDNA51QiaTU+BSCB1YroYgp7TvjJ0n4QhIQ
6B4ycZmOEnNwVUBxvkasQtjjuG989HscQvCezTsnJ1O+IeJZpdMaHV8g3vzKSVKD
qu7kB6T7tA7wN2/9ksCKyh37jHlXWOrH4lzs2peAELKG8CIscrCMlJGmOAR1TPpA
zpBXfnZKfxjcr2bwGFkLYXw/Vw/rMhUw+G/Pj627iIseOsJ6JVzglSlQ3X0aO5YA
5A5vzWTrRkod+KS3nCQ53talwrCyw2DkHqBBkb46atmJKOCtu8ulCjwKgrPIKuGm
thjhrTaODHm/mf5rGPBPaDkCYFe3N/f6dJqQU7qlCGv5gOQeHn1K44AmdoyYP184
O1sDh2I5aEgKtb/pRJyL9740x52yziHN9tMYJ/+yU+guS0Zu78zkV3ogjro91/fL
vKXdPKmskpuXvfOBPdC3YuZIfAMBjxn8W+zXm1tlCvq5dLOwkhlykqYGMByqOqVp
1wJoszeSoztjZVPDl1vV7Tg3I/uLU8pEUzwuBXgCoUjB3vFkNoav51gFvplJTNuA
nJl7hJmhYjexPHWm/nCGucxdN+nkKMAfFkcxQ2KfwhuQSep4vZLz523h/6MQliNX
rS8/Kx+KDFLm2mclQ/HWAkYNJYWHGxYY6oqANELPscpQGAH8re+19WsiX6ubsqSx
zfQZHP10Kl3ZJy+7SzJVYjMSBoKr/zRNyrpjjQHh0csArHsl7KSiJOvyUaeoBmLM
wGMbUGkj1+hjK01pQsSOZaNcGbZ4lSNKBsk9WluQtIscAg1d3Mi9i9XOou6PTp5x
b5yAz9EveWhJNAg5uwgQdp4Bb9WFUxC+yjvcPerfC4mfP8MXPxT5jjfQtI/dqZfm
77iVuZATkEny5b0dKASdDtUmxti+Gl1mys0oR/hqf3zZbaO3bWWCSb/PpQ25rZGs
46TVXVf8DVp2EnhitimZVPxKjL5ZUrXjZT1hy8kRuTr3ECliKpHSVbrsRS4p3vik
zHWNhNRyVfyjYGF2aTWZj6g8mFXUklNo5j4UOsGcupWTN/brV/rllxKqU8gNYmSs
68euVCXtGRerEHc9WCiC6oGVlHa9MHQhGajLJzajVJyaHSs4LHVHXG/PtXaUsXOR
iCct/pZYr+8+VL5TotxTZXFLZVHGQ50Vxd1MtGcWN8lu/CadH7EX2r2B6CIoNgLH
ZLC2TMm3h8103p4PqZG0UM3JNypD2u/2prWEHaGnNlPaza42hIJIvT8mvrreAJNU
9DEZyIp5qQRmkTEvIwhictkpy2HyxvLC2k4Gcbm+4oNwxNmkO7MRGTOlwlyPvwvn
JSdZU0QXpDYntQNtkpS7tEfgefsiQ6SoG7sPIJ132LgcDOOhw4q0PCVb2ieFr44q
tDowCW3xSKElL+1plneifAt0yXclzo8OLeHWHtYSZq5IMseUQuGe9k0BtgN0Nq+1
Sgbu+E+4IjmmZm02gYY1S/evVmKlSi4/2Dkwn4inpqZZsSrnMmPvDuKnLvDzeeim
8IfratANyFN4SyXzuICMl4nCn529cj3Uqgf6QzQJ94HRL2qmwiETSp2ZqJGqcjR0
lJzrcffI3EpBwAA1ngU6yXOkmUh7HABKVbJGTwmHtkjGifrHzo7lV4dV5vd3G2Qz
rZBgG1B6kkuAcRhbeprggoJn7GARJcRuZB8zKSZBoYZeo9mQJk21vtEUorgdcEPn
jl7Wb7X9qlf8cVMEAGNOjzVFcZ7RYtZjHNmLK3o7tto+CvvkiKu/eEucCLNMkTRQ
zFVzuZVrdomB4Rg0Dv4QIZwUsdJQ2iiDpcRD0ViV2C4geBRPL87jTRjYsrAY2Cnc
XVC9ZiYYkqHeT1ADytar91jYmqg2bGLEuc1fTQ8Y1QP3Cg2zGf/EahhLl7HHa5Hn
03J6a7avRAmU4bHI/ZSj0glrjPfR85AgfQfpUo4sx0wFFt+oTAXNdZRRlXZW3Nf4
CRktiw9AWEc14VtPLFmpkb1w/cc1KDtZgQ35iiatDRMYkmbFeCJzRqQjAziFBHxI
Pecm04XjZmB+DPrczj0QV5QpdqokQeDJy6D+YSJkl9quFkxOHxylU3r52FDOJ9/h
WwXoofNb1zHFJte/jNbDLA1ef8759zwo4ThgFkOX2TggoLPvba9I/ykfAJmL/dW6
HEn1w7BMRg8t+oo/UHe6U/lx4GaftgPNgHcXwd70av4BuhMl62eXvqEWh4jlipPr
UGrE8YS7gY/G3fgfLeIwagaRDe2yH3dFmlfZCA+0yS2B+TtsbcwO+c62gcI8M1w7
BHBW+8Q1XF2FsTePKd/2fBzK9yCyaxcW2t6Qqkl9twHholfWpTnVmgh9vnltMXrY
txF+uU/R1Pm/61X9yxO692BKcbF12gzJYfwXK+vVV0a0Kwmy2BK2DV8LtEOzTYI7
umtuLH12FQqxjO6hlfpp9VR3eC1PgTv81UP4mxEKOV1+m4YqrfXEvBEsxxh4BPbE
KoKqMDXrTAFHw8UF6jZODYaaBr/zecGTDqa5N6IdWSaR10B7CCLo3qH6IfFKHRjt
IJ9N6whDNzqOPeVnpfyUcBVkZwRgE831QXg+sLIIJd8Nu/zQoHI7JshSolRbXS2l
72GM9tqz55ztiMcZUbka8JAef1trS8UVzi08CHMt3k8Pp9xBCJvUrk6TNpitZZ0t
EsnLv4cB3ef5xYpueHRMjoDhwp0m8bYLyTovo+4aDzU5DgjwZME3t/oDeoJjwo9K
IPCULtowFBxNjo2FwHQZkPzE8RgCp6jcQ+WPSJRHRTuT3zi2gwFPa6JqguNvL4K5
WIzPXuyZ28K+2l1jXK7T0W2WrC/xtfsUCGUZNIpW5TVzPNLonejNdYoTHcQwSTfQ
dXPp6jthfEqC6/mv/MN91L8ANpcquRDCKdcg5gY21ykZss0GNv76dbrh04wMsw4r
rZcPqfG7Dg757q8NWU2AkAeKx0rINORBcBK3FoBANKhOxie3Qjl27w/L5fIXtvgc
w9iWcwi89BC+lJoqBLIqLBrZyzC+v0/U4D1agNWnQ92c61xRQsD3m0JxehuFz610
MHN93+cBUixBLEM1iS4CwWsDAxLHiGvQZtqFSSDNtpOqXmIluIFw5G8DCeSc+pUS
M51U8ZsPtyJYO9s8n+qJ5bV6UgTkQK3MzCilH0L4wDFxFZN7Hhj9plcRI/D5jzOi
5P+Mj85Yv9DNJX7Mj8QDH4nA//JJTMCuZYuFX5Oor0U0WSlrLamY/rmg3FxR/cSL
BvrhA729+S+zUl0qYIwXuc60yE6DmyGImom5U7NDonhUiz/Eam3i2PDR5UR9VFZT
eQwcvGG38B1RCHBx0ODMvinesCrtu9/I4nhBFKTvTp6tzlWp3bhmh3Y02ocK28pj
W7wAIUC44YquDwjuj8g6ji82RD1WtWJS5xNSEICgBKqk01JVhhRKIjstJsmN1BkQ
6YZrDBCivB+fgM3/k7ttOhNAkMH0ZsABDWur8R4s1BmeQ3HLQJVo+3XNsOJfuusr
wBVU+Rf9NhzECIYPU5Xb15sBH3FKVfXcKfTpBENBlHy7Pnmseou+J9RInbdqTIiG
MZlIChdJ2bF3Fua6hGlInNqO3Lhdm6uhGfT95tcJ8O+bmUeG+QIQfpXi0Bn0o27Z
Irb5v/cquqYEWzI6/vlMeQFsK89RVhjC7YdFPFmqE3/lwUXh2ucQUp03ogW49XNf
55e+ZloqHK7GtUhfsCog0XJ6wY8JOS+80lEFw2HkkFt2P3NMaD1RcMRj2QaMQ5pG
B9wLqz55rFRGc2305ryIyILcZTxzzM70QBvWxKvzMbPn3VI7OJWJInTZWe/z/GXp
SdVLUEHRYFXITQngfFRDDwvtL4vZ0a1GXeXDtubpYtoVI25hFF6OqheaOhTzzhAA
1Bn3lhB/tfUcbhy0zK7Ks8+yM86jX0swSgBvvX3wWy8jYPv/r8TeU0GYZ4JUQKz9
EniRWu+je18uR8zJ6uJKuk6QMDuzRbhehS+7BZ6xqk9KCVK5Ac/cwMyABQdvHSPE
Jz+M3/JChFOM8rhMgRfPs4Zhdk8GxUpD4INoyAydIOcrE5MwuBtd0OMvcIxTmp62
JtTPBSlCCcDf0JtrNOtzCkQd3RE+ilErQrtIqUEqlGuZsNceRGTgPtZvhDEthd0O
bvBIJ1IVGQrPQ5gZgRWeyd+QeEC8p4ElN4x7lUdNwmI3ndtztRI4OqjY6bIBlGgQ
2xAkUCtS80SUC4V/416JsXx6whB8+ydH3Z6Yw/Q9DmvmHhJFeyHIPNxrMwtDat6Z
/+P+YTRIp+TSITdgZtRge+ILT+xQZGUpbGVGPdyzYnghiT28+cqWdrGdT6UmWIho
YH2aPXv+qSVCbZdwqaEkWe4Ewq5U4u3Is7ODYRT5o0EPOEf3kFQ/k/3+JW/w5T3C
aXhg08sS758mLltjiW3EpdIJin0glT0A0ZnLrlzLcOz3Z1IKR9pSTOuBbsDy6J63
l2ZPjfQ6aQXqjTkg50000/BE9mllAZBfyEz0tg7435wWyKF77OmyparAhylo1+J9
QdooOsa8kS2fAAMMoczkUwwNw6dV172Aqghj4X/KSTgeg4ysR6YbaFGeImoxmqci
HizNqdU+X4clOgv8ukpqqIUsa0n0E2UsxXY+WbrxzfEYB84vQ0ikh/t1Dg5ndY9X
o1fY2xWoYix6Umv2/k2w9/xAbjDEhnbiA5stKVKuZysiOXPLtZYRX/18jn/Wg1Ks
dStlZkZpMILrEfJDvMwY2Kh/AGatMM64JinDteY0kIcm0mceG4ONhjaw8nEXFiC8
wQA2kbD11Ik+ZZh6IMzuUTt9rg8PaAat0O10aGC2l9hr19gf6Fyqh3+MiaxOwRQQ
1y7vOG9hvhB4OaWIcERN0HHgqc7JVbsR1gLyN3XpxAHrN+dWT+WeceOVG/trlU/f
Oc5xWT6ZNnBHLMQRHK6qWNiemi5bb7lz2fDPvRpuk3im50NCHfD+Q9L5xPYnZj3m
xGInCnUNOZ2WdVVeSVnckFePY3Xt2oqknxEa4fNMA+4VDXExony8fx7S1mKRuqbK
6afaC53haYdzau0hwf0Kn5NcD3R8V8uhklm4CQnw1FC/Nn/LZHaBv2dPsl6WV2Ly
glq6LOC8aOzkS9/lEW0YQXvOcGmBnP7jT2eOL/cC9E5zpO2PblrmT4yLzPtzzzV3
1mswPhCEDqMGfEjt3TYGpguTnI+xF6hBUx6BWNh2w7r4wc4QI74OXCZvA1R1JnWg
Ho4qHfsM9J3WlytZdAbHEQ6wVSeEut43oOC3/4AcEdRukJL/g0Xe45PIJ2QclZHC
W3+fU2yuKNRHR5M1QacPVE06jBq2HHRhLpyVjmcGE9umhvPwN7JFI1x5cNFkkdH1
G6xFai7Jwso5lrUOnZVjNWPoggGVQNXQi/Ukq6IiI3KODbxvpo6SAJaZDUIxLMRC
WUtkp5w5UidFXIEeIIYnSHemwl9VfipjGG5iz0TPgMI=
`protect END_PROTECTED
