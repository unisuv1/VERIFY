`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jFoed7/hta+v52kWuZwpOAwpg0uo7z581Su8pMdNfuv5exgGEo7UHBe0T1wXyVUG
Eswl9TXrV0Uia5t0SMsYrC3IbPokAKnSCsiZz/O697f+wFUMyBOGF/QbSB0EMr0z
C1ppJar46mzPWlyJ7mpF/kaqe9+ozvoE4bF+HBq2Ycd5F1C7Xjw5uVsUGdzHBjOQ
6Nuz0/hzI4Oc4+YuzGyDmjXcYXia//NM+I4UJ4q6+ZtiXSsPjKwOtwsiiiU4EWm2
oyAMySarecKWW105iKwjz9GPdeXht1I51e5mI/ka64px8SQhcuD7xVXLW7n6y5r3
WmiHGkHLndUPtOMduvui+7Ql0FvhQ5RVegDdEXdaaWxkdpWtyUvkTJinATW6awdA
v5t54SCk/7PtzeTZ5F+8Wn8Y7ys5Ueioj0WciDEDNwvPEZJp1hZno9fEy/LH2IuW
Fg9mcjZbtvVACKfdnXRK0JuuIjH33xDJ9qqcLPnv3kp5ndaQODtfmKoLnLiz+N5w
DQA9NP8I+H5wnCPAr+LloVujFCKI/sFgcGkKJ69rqJCJLHw6WbV4pg5/GLdL/m3O
C6B4icZCY6jEgQ5ICyxj32FhKtAW2DhYz1StYQ6VOIcgu84nXo717KWTh+Kvmscp
fTycJ2D3oCP2WYQzJ+nac/YkYearmX5pDUl4SX5oJPpE30+MEooxkEP+uNWzdMh3
ji+9LgDtyAgipptJg10HT5SW3Mlk3+DhXQlxGm07kgxpOGv7LfT7cJHrwv7my3+n
WkMgOzrEr70mNs/iyQXMTzw8joAjSvSfw2A63bUwKQbTlTPQqL8K5nVM11vEcbFs
YgW6Yu936KQPQiufHb13AflPbVCuG+O7NJkUv7HHZ1sF/ZULVAPtG8UsDByFH+nE
HA9uAUujeyEs3em0KNR+MiijcdEW33YZmZqbDxRu20U8GcEasUo76sV1ab+DD1M6
aylezwaXpJnupexVfb8mSsv4kio/y+TM/m/YF67/Tn689KPXdaZs1UH4GRoa0sAx
0lJXtIM+b4UadMQsMq0mebn0BevLNScb04qLGYKNyzMeLxIs2oN+BLfwSPBOFFJm
3QJRpqumUnmX4i4i+nW9h6TpRhiLE3fGmzaN/8Uvc2g5Gda3+vjJnw0tTpL/1I57
YZ7X95Uddydmq0Esr4mxiqh/T0nmFoDUad/1wQblqIBBOHFKdfWJX9c5tWIsp1RD
5m9siOnWd9Z8iQn8Pf22RFcLQj9Xfgmved4IKT9br1W+IngvK+A1jxV+kk3MLAgL
E20wvAW4HjvpaNAEVG2EnAdgXf4xczXAD2415CeS3xXdrrePnGD2mdMdb/Qy9Auv
IFNx1+JbzewzRadcQRzGpvpCbjecZmP2uqzwL83lGMhjWa7pmznUPxn9zkcIOgtd
iu73NGr5T9BSAw0xYbLnrM/HUq858Hrx/1enrc7820FpQ2kazQBQJeR0OuJcRKTS
MddK18yXc4v/q/7q5FDWWoz5onT7rQcfU6QHJhmuZTmgyDhwcnIm3c5lttAneHjr
8Xjoe42dj1cqcauud3yTJEhcCMrAbaNlSr+gxdMbeISYYjhphVSDGQAP29Es+Ls2
KBRQ8Xh7lJ9RYFB+RKvNoXFgxm7R1G1dKg0YfoaiCVxScXaIyFGLlocG08u20OkY
DH6UuShdo83cGZgEwSyDkYyOeQ8nU9DThFYQiqmyYY0GnDbyPpPixgD8ioMt+X35
8FHb6GZNbPwGeHNsgeW5hWXWmsX00A5W01HEXMRhU2TIC9/jOmRhNIcqHsmuiPxo
cblVANq+/puj5QyBJQ9hP6I7AFtRClrdQkQNplNtu0rb2T2IOhx9WKsGdPPoScx4
Prfqcsi6XV3ozwck5HULQRThXAI4lZGr8t4ikZeuSi0twzE6cyEGPBBzXaipqyGB
aGUIrsp7gZ4gFILuUETgk3lpQlyX52przPXxHm++PVBoh04ICkGwzAf8jNyV8emB
RWbUqHog0wMfzc1pF0HUITz6JnAintxyqpK7LyBQvPpY4Z1aczuHS6Q0ma7ZtCP9
41yVW8hgJTZKf1YBrlA31cII6pHbocePjcHPfAZM+KBhZmhA5oUg6H7kt/I1hgNF
KBOEiOF+EH7au/Z52nbgocWA1L4nAFuE8ogCsvnbdPME6l2QGcXGSCvnVqmRbrh1
+W4/de+3zY2N7yoR4faTRrWw6XvrCSk48fVkUBsZTyLzn4OCnt8imtglMqNBA/nQ
/WahEd1usmQosrEyvu2IfSdg4rO+Jx3XKy36V5/bO79TI3a8qojNYgjsxUmtfjI7
nt2skSdUjFtDoyPqNBX0/1bLDClRLXCs/Vaub1jCs6uNNlHLUciL6NnnKx8yigKP
spb7/qEVn2csO7r9bw80P3ZR/AYrsxGNfmzvsEn0exV7//98U/poUT9SDxZg0LTf
uk36F7mmF/nAeLFuiw39ptOE1iQwQBmKrTX1bKCxVKaAfda4LleRlnbIqT7uM52X
yU+cfhFMMii3rjenhTI1M9TX7Je6voIspOXjtFX2OIW7YuHyhCTO1PtrY8eWHs/u
iRbaB5xAaK8OPd7xsJU8PkhIYrNzNst2WLzQ3coa9RSMXD333l8IBqFDCVlYKrso
4VuSar7/NXTqHEYLUbdf8zCagEIr4fgHNoxUOeGg6J2bTT4ivYnlziRICquOrVk8
4siSNe84YstjzWDS1bv4LmcHC07iBaWbD7Wl4/Tx0Mr5/UJhof6OmErZXieRfyqQ
mY5xTuLf4188dpOBdaXClrrzeQ1k7Xa46IEa8nOlbF/blHy0IVSl4lRgcdifr5i+
V2bm1LhSDtbiUNG71QPVOqwRrrWeyVwyAZnmlRIy5Sm5WD1m8fu0S8SakrhChjMn
Pv1tPJkzYioz2AewUX0HSlEPASpJMEPXUbr1mT3Dn/AqeUMqKVE5cefIiKkkXw2o
2DSNNNnrJjMXSN16S555k08aQWEz0RME+5kuoXzAsnb2jLCu5wo1sBVF3E8YIjYy
LYfTZWeghIEZnmKvXoSR8az3I8KIckQhwDnG0Ya7y6IrBOn1uhP2eK/SgTVHfJVN
TSaybZ+0aesFwDnYx0Zqgk+ADKzNlTOr86mRLzM4w31kODOFjOBrVPAF2WTa6Kt5
BrxNbyOwwT+8T5/ETKona2LUK1K7tLgHWGODDCIZA22RnvDnB6PPBSdhmuIpRE7+
GesWhaea/SBGQNcP4iDqQEtbmbO3RWvMb+HIOoKK4ZdIkP/4NfkyC+Mmj4jOZ2fx
z0WXHR+XhIdePUGMdKtDbLDwBOYeJcZMihU0bX1gaUCn+z5hmLjAz4DZ8lP+bkPX
DVGh33ujjBwvIbisB/HeLsOWyBMv3dO1qIPEde1IX6fcSWonhFWOPBdx9yIiBXJ+
8IcoT3spXOCWe4oPbhzEZN4lF3LcdPhjatYXznOOX8BAt22HaYz30jKT63Uwn1MW
zcKVJnifLZK+MvO2KgGBn7KlxQsvqZE5WahdRZm+NGkUxXIoKl8Z90hTIRKrn7kO
8sMXnWGVKw4EhGoywGae6x64ZxEXXmQ1uNz667bxHfAaJ04Xp0NihFsE1UTZlYFX
Xgp1NHXx56AGb8oZiurH+wz1vRxEeX0TyGztkSD6pgrztlM2PejjoYpzp9XvI1w7
BWQV5mZrdoPjpGIcmDzNH1Wey9XNmu6mDxyiHWqQgrHg4OHeafqGrWPegsSBwlTd
nYyqk9wtwMLVfZ0dowpL2Xgn/Q3OYmHJI8BF97ikZ1lm1LSyQs728VeaYllpTv5c
64wPrR8a6fZ3tV1uvJHzqrUtlnpJRdtvIUfsbD42P04seis2lMO8X/yJuMZXvL9J
nBj+at65vqdhq+iB/2AMk3idNsHgLzvs/7PAoIs8pjeJQ9ZxOflKO2MDty/3QyAq
Gn2YlzPu6nxHvYI8UJ1uC41sQoz3EyFcmtOyRA3gNbchZm6wF04W4SPMR4ArsEFx
+ZENsSxj76FiAoS1E3/vLGw5injTuCvnMa4zLsZLwu67KCkWNWX2DC2i0M9Du13Y
6R9dD20t+IhSgBFCpjqcludhcXRpXxLlBwZ8xfZXy55Tou5D0Bdl5DVsVc+7HZKi
/JTb7BTRL+i0HWIUFG68/VedpZJhfUCrwuhKqJAVPPlSVAjuL6aQ/3DcPxY3YSbO
67DuHMpPM8u5imr5/Pccemq48Dl4WYL750fdWhS/IGNLIYOcZ3L0yC49yuS0vWtI
W5+0CcdjXidD6N5t1pVHDPUTEABBUHtAQnNdptwU9K0KZBkA94ZslrRqE+Tqgwi3
6HjVgeM7lyawffWwjPZV89TePx1mN+JJTpksuypHEAdD6d+2bZkIL+RDazQOa/uS
AgpI6Pxu8d8Dn7cCk9H434peNsE5JkJOcMmYGzaOMpDWz/bK5MzSYUCsw1jgSH9a
qOrM4ucyUey8+Oe6FMaPChBy6uNyZoK2mMKN8NDTyfkyyOPj2rNa7WYCu1DVYhEu
vDK5MpHuAoK70kjAjStBeqvgkbiYNPyA3bS9hr1Df/8T3ugqe5R8IVeyAu88TPL2
Xz0eG9GoaQSWmI+f5VLZ5BTVSmL/b/pHUyjBXMMbadqKzGaHvcFEJ3M6TF2JpFJB
SYcsOCdGmzuJkQwuRp/SPJeIWKGOBxHSgeGhWd0m3JQDRNiTYmoT/o2iIqHbYe3q
KLu2w3wIgCNiIOJj6OMDOIRO4db+0ruNcoMnEOh3BYfcGzZYVTd12g8aKD77cP2i
9No3kyt/k1dv8frMTNiHg4DkOnft3st0UUkav4igsqkEXvAWVGdWpxatrhjIv9Sj
Khf/PkHbPm7mWE23sP1D22du7JhzZ6CZd4plJDlpVRVP4PFslEeoNwIZRpNkaFb6
w90U5C523GMge5+K7qlWNJ0Ux1FJBZQXrA902x2qiLI7jIPnNbvCj8Ut1em8NQoy
gwADeGwJpb+LOWKbNfI2DNXAXPL3lzlLTLX5SjRx1WLwsgN8zrrPAKXkwWehNDZo
o3s4vcombW4Mubj7jiiXab384GuK4AFvVbgmisFuI5LhwFXr/bu/ATn8+ujZdvBT
CvmDJy8TEmBuNV+HdwuhD3E53Fh/bzfP2bOdte6WLV9XxXSTw1bEalD4eHvPfHYU
8YnaP+UicWp8s1owQ0kTT2GOYRGBV7gstbnGxLCuWbJBuRlZJ/jrvdFH1s5fm35B
M9nvPhmlgAa3ryU0uoXLdgRQ1nyrXv+O6RVx/1j4b1hvH2AFQhN/IAxn0E4XcfnQ
6kv210JDujn3a+iujTs8piagXlpjZtI8WyKmwj9JaLK8ATrTXtVhUz54Zp5lkLo8
eMgxZgGbiStE/g1yMrbe2wd/CHGdkRdyuyvX+D2skabMOM3zTvJvAYesCIZp7ypP
kxURSZ6I6V+vCimZnwy+dsAj5jswn/POVHB/5KsIk0tcqEE7oCkvuve8xG0lqocR
UN6EfkZipsmEHhDPp8L8HwN/cZZklaCnD8nvsePDt2Uh09KI+dlreDnXgW/YnWkR
hsoMGOftYBUXkgSZgZ0UA5EgCVgPULr3TaCH+tz4fbHoNhVc2yLrbDYhPM3kNAeK
PU5Imo0OllBC2I3lmmJ1drogirIvyFdVzLu+BZbMXrlHza8JyVOafKb4ZDq45Q5R
sFZKWZloyFZIRO+DFPcQhJCrQcW3FyyHN1eP/RbYiNFA8QM0x6UMB69E/70Z3JlC
dtA2zN+zo+izyacFwGT4qpFHnvqQCNv6iiCszXveDbTBQfdB/D9GWrpShJbugRPY
hDH9aPCsdlHTW0DvM+C+rglD418Dt36KPkVIy4bC8G3I8H8NSvt3+lsLwiCDOcOe
vO1t7cOMlfmYWlnuq4Of1wWKQTYAcNeWP2MK3JQZ8iiu1onDw2tPPR865oSCY5H/
MYRVwb2hKpK4k+eozo4+UCEA/RGOkxnSkjCttfr8ckRg7eMxztxEfBs8sbWMy0OH
lAIdQr1jiXaoEYGoK5V5TPZIZVcNppxSn7ZGmtJG0kwc/mTYqFvFckC8BEEim+sQ
ou15P7hNsDgwBVwWKaCRLON7WJRHPSGrBddE1nCrDva6GQF4btQG+iMoUCRFVM6h
r9f6+YiynhdhAZ39a0DriMXqyHSdWSdfcdNPdRf4LtHsx8TlqFYvxdLWQSvAFj4V
f21A5I34sErF6M1coF6V2TuesY6k+RmLrY/t90VwkRbBACmo1BwGl7UaqrUNSWCQ
FZr5LF2af7+4SEnvH0tfmdFPPGffnc854jg6PRegOzOKgpL4M/7Xs3AzBjrVzDNj
5WLILLVK0gvYPsB0+VmtRvrcxLiB3/u3sZ1B5lL3uBDBcMttuWc0/69CC4i03sNI
KNvz7GJ+C1OHPFt1XFWgM9E4hJEj9tl4Z5bKYv21g2e+p0bCjo8F46cvbJDyYeBM
/x56cMv2aQGOkQZ6F61fVu+vXOMk9q7XHeTm7YogO1uo4bgO+3PCQJQ9KKBgsxmx
KR5/7ILD9u8hdNH7YWOt8Tq9EjyTEWLzpIQMeBHAhjz2avrh5K9YCDURMeML98iM
m0uEGuBgKCWq0dUlrAQP9Sb1oXkSUJ8QHABn4SLUAy0KC0stNsO3DqrLKE2K82FI
n+24HNSjXiC29lhIUxg5K6u+cKZd9cU05YwT9Qp46ZqR/6pLEBLz5c5nNXVXYkgV
XCa4RVZEua2aYGiLBgeHfGxVF8HALbrlDPGd584Cqm37thHIE1Rk9wIMzEgtOaHl
RjiMn5GY2QIn9m+MQw4bxhsQc+j89XbMX5z/B0yuhW55pLeVPULjg8NHl+GL6LCK
Tm+kG7DFXBFJ2UmUQl6qLbMbdPIuayDOHGy1e68X9HyvedSHuNAJ0gAwXuCGacsq
tVLtmm//RJhY3kTKBAdZkkFz1u1w2vMzT3RvxnSLT2fmSFdbFsiTOu11qR4nKm6N
+9a36mZ3J+iWPkkVtp8S/lez2IRIKB4a7zB872j9wHYPMT8VbsACOBYRyRQHRa28
0spY6tvsmOv3dqHNP/oNYtc2GnvzJwJ5z3pD5G0mGkCHGzeLIEKRghya9/Vb3RIs
5axvbTCL29Fo7c38H9mlylarPvRk2oLOG0EELXUD/CvyCZU+BT3LNk4Rk1WqGT5d
AuDpyGl37cAy7X5t0IrXarXrAzcwA3rt8uSx5TraIn5Qy5C8rKpAIeLJAZYdwBOI
1whR/E4z2C7nVB47bEwDAR2ZQagCnWhfnPEMOeZ2I0CQbDF98CxGpkcTg/lKJqn2
ZOtEB4Jx8c7twT64Ta4t5uU/I4HNFGKbjFeaMpc9mgjWWxH8kWyURMvqrIIOutKn
82bkhCunLf5j6/eChL5gWGnKjXaHn5/0nfiLlQagdZrKXG38eqJsln2WjQvkYEPd
tgkPHn8RYb5rPYaGRSaDaEPJ7HwFm4jOqTsUjwLehKgFmuccfAxm4Kh3qBscLDb+
n89VP3yG+8xfL20iDrBWxlbWE7YZ4oov0+Cco06GshTDpFjshOvvj8WnZF4bgtvV
LnXWGcTMiBmjcPrO4N6CrfzP66CoVXsCHV4XXMFuzZi9jbXXCV6IfJP9Rfhfxtcg
jNIwcgbhL5W9t1s8deM0WZso0pFLJzUe8/3FAgwVl4ZPHhBj2rlA9M9GT+9Qq4vR
fKLQPQRulrvS6hrPXXzClKCbneSbA+1PzJwkTcZqNU3iLQ247xBX74k9F5leAKCU
7bq2LH4YHoQFXtUZ+2iHuh1XviS4ZChniaPpEvVpP0IQ0iWIKnHba11S2uGiJOpQ
w1q4Cj5HSIyvC31Cgrxw1PGvznd7+J8WuThmDiGIDmYrSqASwWVeocwhgHALF7BZ
ubJ4R7gNYwaKDSGhiPtCiIg1vaOBplSl74UHIfOvptI9ngj/IcWnEdgcpo9CP7BI
zDEJYDoeetJ7TJLSDJNN1CXzR1V3S6n4UprYv4X60F4AeBGetN5k1/6xaC0SWMEa
+ZbQltqz0hfLURkjIEWKfuqMDXBEOUJeCFiWL/33au0H0yh1FspFlUddxQVNO2S9
8gp0LZjmdSlPYUe5+/Fm8s+8X5JazVbwm6vF5+YOU7JcTKkiQyD9CJQ1M1xL56p+
HIguAz2J6N1rGuvBIEQqk4wGHaoCy2xBv+GU5ouhRL2PtgrxawjJelp8ldhzXILf
8pgnVvZRUu+Tei5+n/6uegRI12ypH1rlRk/WyBXxpOf3/SQl4/Pnu8vAkA0Wqa6X
AOWrmG12iAbSvHQKpo8qdQkxJUut9TgGaNljF3jxMb/fTBD5GV/I3j3wm6uWI9pc
TmU0FN4rv5rVJIsNNAmIJzeigYcoQY5kLcKFdzJ03izSKvOzJjKycPIuQ6SJnvif
7GXYmtcH0NINbP3aUbHKQVjEaj8ClzSg7NT66pW5W06nLl7gy6PZkJxBTVDYerhF
xFbyoUDXR7tclq7JRy1Juz4uuMh9ZQxB316S9/OKia3kEPpVaaHJlHCj0H5kxk7v
PUYxq1ttAfzWP4qJyW+F5xi7R8cvTEN3+m7Nvf0gzogfY7xMWkZp3KjkG08XqbN+
6DZPuoZx7FLMwh5uFBt33jUy5sJf1bYYlt9lWfR9p/sbw6Gdw2xuvB5gWmKRTlb6
GWR20K6H4HzVpxN1JvunkyzgXRFXPgFcPysW6zxK5FvOjEvtdl4JvNEeunmeE5f2
RWqjksZEb03C+y1YYQWTYdLYhEYQUuTG/9ouQ4vSi9Gw1S+6E+TiebSxboiQxKaQ
fQOMg63MYsJPaqCskysT9qDhfdtTxvxvcCaNtpyI7KMJtKgXiMEOPV27F4tQVohc
FmHyCj52HRZhNzrrjqxJPUbWG2NU0nVKwFFbvG4PD13Y/XQGZZWGqTI5D6VC+BJa
Qm3+Nn05Jodes26QZSttZbz7KYj9bm6YvVnUXOYg0NzK2x53dY5fNCHlTnnM9YFz
aJ3U2Sb8NadJF4iFPHOt8Hja/vSGQ/4+p8ntbrWQU9WLg3iS6bS0ZQbaFX1aGEDI
IIrLC3awdsI4monmnptgMW6cglUmwoFgy/qnhMMaNyoSlU2dDvuFrNjbKbFtMw8Z
c/BCFH2mAqL3npxl2sdikcp2IIz+N2dxjOSae8aqVzdtfsUclOXfmB/Uvsbrga1i
4c8Mstxk7G188M/j1g1L5ViqA0LGfblr+IkyxrPbm2eueFu/0FpKxyUavRrZ61qh
5btFR87m0P3VVWCaA35z4vOwsL5YxRVS4AuA88hYFAPBXhnqyVRi62pkFyBTWN09
WDCu9S5U/R8xvmorQzoZM+roSiM4QlrEnyIEVHt78sFvojeOlNxEPIU+SUEXYHvu
RAmMZNiW+HVfi0BYMDWPtXSCezk6tcU9pAy3QQip2sU6+lpiQLxu+EIYWIm3BSpR
QbhoxOJ8GhtKeF1NwXLN4aG2fvEAbjkLWIxWf/jh3V1EcNexZzf3Q9CeZMtCbkkD
jMGHY1Uj+YyRwuMRvtVLjZNoYqA+zy7ikLYuyx5qSBryfQV2wvhUmqD4znJUjasw
ZsdFaHlAku9KcXRu7jorVB6SWF2FLHAv6e/C44QV7DargAh9rxCJX9pdWKUaaEbv
8b8O6xB94H6gJVc9+omczRABJc1Nenpu0YWr7Enz3u7PCFO9RV5JW1R6lYe0bpZQ
iJ+lWj9dqPmyvndpyzkNI3D1nZJiE0NNopAgv7TUxdcPI2VI67NDiO9wqaSKvmQ1
OrHO2qK7Sjcp0FskGRRLiirLJIJJSnUte/xEWbrzhss7qBeY3dsrEm72KW5FtfsQ
/tIfkSYfDcEkPVus9iIqpqZb3QV4/gIJqgsDPAZeZXvOaxs0xKKhnMOz4fbfGOvV
zuj2JC+A43pas0rk01+6OlNW8LFq0Jvo9FuzxHJbm43acAh8huQw0PYJIvAo+ueC
bdLgKM7UKF59P89ZDAjRKMkBdBwDSR1dUA3GXiAIC0ulbWbqXnkwqxt3Z8kU7C2z
ITN9fB73Cfr8X0UYUPFL302qg1LU/wRuA+VKuHQ/VHf4R5GwkgQzhjn+MxunaT9H
Cai0VJaqkwMG0G4BgVz1QJUyMuPBCUvSajZaCgIKzIEKhbKNNPWcrhYLZWAFVS/p
7wtjzRgY57MLPJikFZxksD2oXKvM4uj8TpzamfnNh9eUjGXAQhLO2nQjbwmb2h/Y
soGebmwgC+W2NxgH5IjuZVPKDhevRM9LQ7DnO6aJVkaIU6lB1RjAImnV+xwm8ju3
DwQ2mVtwAUV0fM3BDiuuaMAF3HrlsITXusXk4hiNEEgXmNl/HB5srtUjsfs8r1et
znD7onggguQgnxQ91A3mMVv3IWq2iWO4HwzRyUK7O4jsuhnI0oazalVMcCY27xiK
oB5LRXCZCXwnhBp8xYWjeXQ5ObGp44qVg7H8U8ORr48L6GO2YafgDQJaWCw44Ss8
L8iCiWk/Mk97k2YNmi6lHl+WUbnsiVTJNNUO1z4y7iy/2zoZv6Tgie30w6RcZse7
KppXl6aAO2TEkF70IyGI4xTRV5n6up5Hb+17v4x2G+Ul6qyC3MXODwKgNL0z4p8m
oF+ciNsWB3bsWgCSCqKe0yvfoNLFKiQmeSJYq0A/roS4VdgpN3KdTxF8fn089WSN
L7ECfsPvlTfsNPcyJzp3r50Yrd3Zf9Bh3D0eV9J0wQ4eAOLItVDTXFfxh78EBfig
QBJ0VpI7ElSK8BdMxxRxufma1AuiO/6KJMoT073TmnrOGOoBddv82xwZZkGCpwSC
RUtHaWHk24eCO/ejtC84f/cUYP/0YMEjn5YZD0sY8zHV9ZjkckaaFTkUIgD5Mvhc
4Y7zC+FOdv3wv6srucDP/DNn4KEVHWiOzdmZPzF8xFbx9KdS3HEUplb0ITJeU8Uv
FHXDTXOHI0XAy2G9cNsKdy+eXaKszjGCA+Oudh1pjTn08crGiFbAN3s6X06F6yHU
KfPCSM//XGgr0I3ZbolKEHKmTUhvWRZWnlcnk9BA3sN4hytKojdOeMd0LztONaiA
88rpTGYlcszcf8nslhVIRbFa78WM7BFnoQGBvp8O0RIiTPS+JSAe8G5iOGvw3oU5
wWU2G5hllSV0aY/Ewg/2EvsnpK12Cebk1XJdxZj/n091QBVEbHkb67d4Wky1Vs3y
OuwdIoy7eq76JjVwcyK8CI4tgui30nCGt05DoKUhunJuEupCExtA/XFadXHpAUf8
qDN7kTVEq91c6voKJh6kwQLXQBtUcXMpDq88JVxOM12XXH1VPG0zqjZfLiO0l9SR
l86CNSNm0K1dJplhgxfYvrCL2rFhxEHHbqwsXHe4JB76w9huVI6GPCfBHjmf3IJx
yfZ+OAtk4wwbh3/iB39SdtTQoNi0Fj0gqOgkDFAJlFmkiBRy7ntqxP6ySxY2uSiU
XXNXU+jDD+xMHhBpVSSYQEekv3O2fBLXiDBtkj1f2LoG3tbTGI04s+LIia2WLxsZ
NJrOPmqUDQrZ8L8fvAcqK2Sis6GSxRVvhrcUUMUYB7IPbP1//0i8nlbT3eQeGjef
hOuLIwVDDFSc8zs2qDRsIWWpurBMr1YbSM0nyOd3V0dlTOgXNtnBlPWZxMaR6dTW
u/bdr6kecoVsA4jpqhsXL8Bl5nlfOm3vTFA7Q5EeuGykEN5uKCze/bmIzwabzo6w
xSIccMvfkgElH1GaMSb4rRLML2FF0t2y4JMU7nEs/0gEgTsUhiOMS6j2LOiQsw5a
rI7xxNWIvMhNZThCE+iwn2Iv4VqOKQA5kTasEHFGfkY9H4mQT0lgp5ckTzSHa0fb
sL7++S2yX/uxsNv8mHEap86x5FM93R4B8gwAmjka+o5MfcfAJiISmAtc+iAnpaWi
SUmtBAOMQE74BikBp70OkbfQbQLi5jnNinDpl8aUT5r7T9HeKgpITyPl1oO9k42z
61q35P7rvMUwWm8hJ3DvfGd0iyiv8JtoJwPiZzsCZS4hcKs1PzZ/MBa7H4GKUVHL
QEhZRlbWilF43EDITLfVS6sRMtL3YA+Tpx1pGqOGE16scUq4GFeM8tSDhDKbMIDj
xnvpVoK9Yrw13VfBGZdsGcJShLfkKY+tK3iUwga/kyE+iXVkviLqvGpOodTd7uDe
rF7+WqglP2SqpcWnTgKex6m7OUpeVu9t+upbKa9M1nc4dQyQBrV18MpBc/ZPH3Me
2JFpXIkKT/gnz4XclXLekbCZjQKnfB1H0qYGZS04J9FxshrQN7YehHmZWBh5Ilne
fxhB2B8wNXfyIbSJ2eeQ9RUu81SnA1a3gt2mQT+MLvDdg9H1OhTJ/a0YJPtmIKC8
oAfHbibfJ3lY4iTTao0gmGECKFlamvTMHp1JBI+cAq4hKv4KoeJiXU9dFi1vNOBD
NGSb+J4wN8wu+LUFTGjJKswNz5rLcQSWxPRpsklHLXrbzw57GME6N9T3VI6c7bwW
hr1ngqM9VZvpdUDYMWuP8eB2jHWfC5jL1+w6CNOOv6+UuEMwi/SDPBIz/Kg/zzv5
KI4bJlrwjdIa62ug0Z+xCl0U2imy8L2NHMeBP1BCycx252KS7HtGNWsZchiZXOUx
yr3SlEPaf3QQ7+nVoYsbyufWFcN9+hj4X4B1W+ruHgefnOsENnM+yh4owNTZFQ+g
ygQE6NREbqUnvW1kgxB7RuFdQw5dk68c4rxDxnkh4/EdMGF7nKOr2GdplM/lQFY5
fqSk6rDId25iTDoTC5MTmGoxSUJuMaMcm+3ZMnam3ZudbBYQHkIB110mAzc/3twS
nb9AwE2x+4mXiT0Yz9WiCYXgJyjokkHFnynHS0fBMh6XQIYRPzLr6lhBxFfoHkAj
ZIQ7vtjRzrS2BKdYIr/XP5maOLM5q+Xl6SYoy8k4Ijft9OmpocKD+0CNOygQWN+b
2A3vwwxLO/jxowaUNP4Svlbgzau/z6qAO3h7yQoea67zm2Dh93bgw1o4V3VHF/z8
yNk6DFKGLkMee68v6IjdFv1IRs2K0HVYV+EU44KorOgbioBH6pSPqPbJpYlT0TEr
oQQuhXUZekY1ol7/1to9IIA1gfZnG+2HEGevEDMcg5W8xW6VcuE1AxYM/WGIeQYQ
FRJSTkbRoKRZPRRGT1eHn4GlbtYQf5ykBDTFGeb/50zCpz4FuHHJ2TIB/kij4ugr
BNRJCW6AcB65h/Bay5AZcGohc/pRJd0RISJbjXJ1Hek7BM1o73XQloydVqJSGqcu
KZR9g3tgGkWqkTC5sh6sAY5iNzzOJm/6sy9u5ZHVdE+k178KysNPYSWXtllLjiL/
omWdFnwFOi+YtBnrd/0X8Dhe6/xbpEBZxo/fZXlAX395o9zYSIUaoqS9UQk8jZ9m
kB0gpnGyk/25UtFE1GvJniI2LQCDVcpTdcjlIW6bDV/cACasd8uCkyfGpHxGmj91
RjBqou3X2h941hDqqzKvs9tjogxE6/FRXHEOCvBBG+VA/ellucLxafNdeDZSg+y3
hhlF11117frraGCGj3/HENeeEu0ZavqiFDCWRvQdj62+Ux8uV2w9akGW0ZN/4UVZ
OS8QxUyCAJWs3BM3y1aKE0Q16+hca6/wDjyrehzMVVKKe+M/ItvCNA7+iMHicQcb
QHjlvLy7LQxvyIXSLH3NqRzWlYteEcGw/+zB8Ad9M82UB15oNoGkEFm8tb/6Ix49
L2dMvL0OEWXKUTAjKOa+ol8sCAvmobflhYQ4BOYOICTPLCG9D2DMySvpdsytan9m
AHRLbiunRux2ZNuvSGt/QUmdSpsMjaWAp608/7CdRxT5wsUhJU9XCesTMeu9H4Ui
t7ED2QyWBoyd8OMOc1hWovhoj0ccud0ckYnXFf9fRDU5kl7P7kwyAw2g4CEIzIgr
axauA2XSqXbVnLScuyViTAptja3FOqaEfekJwbocq/NDcBjD323y6YrlEVcOOfFu
SmyWGr4zNlBRhOyzfY3H6j0kj7R9sSD1cIru2FjHfokZbH+3F7JS70pHMCYeIAnK
7co8Hdp/vPMsy5AmVuPdjYBKYru1PVhUi0cpkzVfrFC8Yax2dSN3PVrGv3RGNPTS
wSxmilN7311z+AA9PUrJYEkz6Mgt0u/ED7b7Z+xT4BLIdWXg4svmWGxyWfauBABJ
TYWPmREPuTz7DosIMVfmJDJheqbZywDVL7G1S2+DikPBlqKqL41mA5sRCgCe+vct
zMkWSKxGxqbN3SpVOsyPTqSd01aOHaQeG+X3680X/oTw+0GZEiIsUSaaaE3mb+iG
YeObLiM0v7pALmaFlhKV5dtcJt7vokUPxL81ASEjwPicRyDvrwv/tT+5wcT1Ray6
7CrhH5fCPYzqFGtAnbYmFocv3IwypLFdGUl46gN9LXb1w8aqEd/M2EUc02D0K2B7
iFSArHUR7xJOS7Ys3mq+nCnHwRppP9v5d3WDsLyEiuGdCAGwermQPNHxCliNr13q
DGUmWJFxgY3B1lGjqSz7ZDUXujY/kdtEUTDgKG+azsSHGuAMruiJ97xMPQ8tCduT
+LnKRhfPuytYYQeYk3mjyyk7lcHm1Me/mpv+ldbOtQY0TC+3vkcj+8wg3YJ06Zff
5eR2m79hYDRZzIcWtC+PnX4rYpy7K0FZ1l2SRljwGnqBKiPUoCF6k3K4DWc1OUFj
vAF/C4Skx9Xwnm+skuGS3N8MajBXnqZ3yv1WKdWRHPzsmHMMk4RfkDRrOGJgX7ox
xChydCIKYvPUtl1O3wCtY8NhJXJ+/WS90qzjtVsRAXG2caj6RzOqGMO56vTY86NG
HsTOwGx1SSHgUjPm7YeSEK4zNqgzHmg633AvfVIo/HzPv83M+yP8UOuAmotwL89m
nGoV5oNrmI7hjKGni0G+1BIS1quyC0gh2Cx9CseXoyMm8zreG4V/MGETIzZ03HWO
lg0zAqzDBEP/5bzUIFEoMlMsjws0fwoQJZJxEOAr20T6XipbWVyB/+6fu2FnUSWe
CfvLNc8USABL/D1WLmvL1dD7vRsgVxwa3HATsLzJBc+79LR9Oc7Ilwk5MrhN4X+W
cZlXrTyPR6JK9yvHNhE+U0VjajLzi/wVDee3m4SkfO1dRiY/qLutxAsCTIWdzUB8
CNIpLBXtua1Ay19W6MGs4XfjfG/1PYqQnB735e7fUzV4Y63RsqNRXRBg/DJ2fMk2
D2p7Y/9NQtmIlLaNiEHQJxG15x5itzLRMmUey5n6LMFvtgvW7yQryppzRbUCPeNG
7A7stlBmK5ieCuNqO380qCvqqlbsrHJuLWLmGtUhygpX7MKabSCX1kVC3rfo4RiY
KnJ49NUkcTpgn7XqtkVWlto8wGKayrPZR4V0AqFzYCA7FtFDX6OND64+HqdA01Xn
rEjLm7rVB/brB8tFrNiA/nPhiJPUe2LEMge7baNqdeSX/tA+Pg39wK0p/99T7xbz
q+fJt5ka/Jeigo0yYTcS82Cj6FQRUcUF8MoyjkXSCDoRBoARBEyYjHw3AyLZw8bQ
xq0KLHg9XH7WlxnNQpp7iLXe6coQaQJ3+IH0GUhyZGcnqvK7Q11seucjeonQ/pHW
Lv/Ta73fBBzMgd7F8hD/zA6pvF6O2UaZXRbS0ajowEVkyYP819b3RW436RahntpR
nDc/w6k4qFsTV3G/YGU5llblltou3XgYNdRALIj84xaVJDvxSWQD8yzV1AO0ph2+
BMtHNcGGsSocYQGXu+NfMxHJf3lKPJWrQVprLh5JTf28s5ACFegihs61dQrUkjzE
DhFqwJdo0zZUGfL62Lxn7T8XnVQVbI1Kl48foYoUhMK3h4ZcDkJG3uquuxeKeWvX
R8Ufe3eOSJyaESO8JMjFeB9rNjoXgsraM6Oj3nd6CBFjTbZiAjiyjqDguehtFDRx
VBMro2Pn/ayymHtp47Dr3NHwS+PTJfM6YyYLNfBOfGEuXvsBtHg7G+Xn4TJO2YXp
cXkC5khCSRpc5FL13dVPkYdUIj/XbntEtcCQi+ucwvsbMbjfw9eysES8SzpXKR2C
PpfpY5POQcdlHd6qCNZFAankGeicDd1VIO0POUDue8JeAY8UN/7yP5PrigNv80or
ReCAEzakuzfshS2v3gs/D+L9q3Puhpke1AVGQGrzgeBF15/TDna5ge71VLkrxzst
eyfFK8/JiFAL+ErwpABxyDFW4v6Rw5FOvJT9TzkoeqAVUDEJvp/SRM64kvKWVI74
1lbWELI+Ai4LC+gcW+JsCJb1SM924PoBHUFWLlPcYBq6PrNh+EuuCSAlz5WzLNMT
fIn81J/bldAHzwWSsPhrF0F0Qjtr4Zh16FYd8sCY9JsIQc4EG6o1LFIJ9YGs40lz
9TEpT8sxJ9kBFxLh4ZnfrFmgd8CLvOzcymC4z688+nr6VBvSKQD2vwBbbUm7ZCJ3
bjjgjJO6bsDLhRYqKiiBFcjFjFRmNrN7gxyLaYlQP6ecTBiOqDCCnXj2igGiX8LO
b6ap/b7/n+pYp+zcyHrAVHF8pCJwhLlPyGXbtsreh8aI4qH18prH0SXC58WUyG0y
HRiOUW93kYL+tmiWSptkVTNn4d4v/0AGsvpxB19OoWuAF/gPT5Y++kcpJqpMKLkG
k424vFepAnn12kET0+6zhid+fN5wU7YK1fbLjTdd5Y6y+tYjmdF1OgOQkiKOO8LK
wtCRV1CbIUMQlt4kF88BB51D+2zn7eSaiHuo+1JMqEtcQdPkQlH0ntZmjsD+nNMp
W4uDHKzhOGR1FFAsiUzOLrFHHUX8zeX7mBzwsZ8+wDK4+Am0Piph1bpE33GJe71O
BakcjAODmPYz3B1uBBcHM/So8qQ0TtVNRp9GL1skNuYcWVkHeA4E9LJqrfL8rJ0d
+RWe/wRMmODEZk+Jnye9xhHCE++YJ/CyeUuiNtHLP4033hX6x9gminGFbxXn4Y2X
VaVI6P/7lwjji3ZzwgbtGnz9D7l95iZOmLpikXy2TOCRz0Qt6zmDU0OZpF7nsqRE
LnwH8WZUpRD4xE5fMET3uCoien4QUVSLTYN8/6KGz+6An17oKsUtTEY0uQvUOkXG
iMNVh1+6Ee3S/81XXueuJ1fKpCEGLXf531zSIQXgGMl6L+Q6CyF4V/B1rF3nBk4q
aReYGCDqFKXGnFomGuqlM387y+6CDa4Ta6UfiICUrqKFunGUT+xkLmE30WtNW0fG
NJkkqz+nhUxpFtCXxOO8ATMahypBsfv8RtuhxLejHrnK4921Iu9fYUivjkQe2ZVq
zATE8yJ8dE9hyazVOwUZUSnMlvsP2s79o9EaShGtDTIpzYHzckXR6+cc9TDlpHrz
Py9ZdP4z2ZrTHIlIipcQp06eG27DgAJARrP/dJ3PAII1mJ8VP6jopnyEnYrXU3Dr
u/ut/W9Mxl4Vnn7fjL2yN3VBem1FlhQccFbCWCjooQ4+aEEJPWjdMchogcjlpvYx
eLzrajhk93H0JTbyRnI/4P82v456yMDcZ6KIhYDZeEtfvnx2qHJTwOoShZHSUDxd
D4CIvT+IUBmpDA7i6dK8x0tOrzG3soop1kNpQDixa8APC589ed+WcGNU5A4RkW7h
5Quz/O4UceZiDQfHCRhwMSJZacr/nRvpUD33jgEqol28XYZepzFzOFBAg2eCCW9P
qzeD105kF9F+t4BIZK7wrnnbghFAvgA2wpDL1dMhJENSgQ5oD+WWsp/ZPjdqc15/
QuJOU571qcE3R/cPjeTUKjYcAj4AUfnatVh/dE32pybgQXeR/dBP0igVrrYlgwaI
xAqpkg09PIywIuMB5RGEW6Ea+MpYoyRqPdaqzvPwKge3MpRmmUQN+Ha84d6epKEV
ufI8/q9vkgCWet0CFau/dDvVDvd/NsZfetDj7YBRJApx/Fg1wGyNJI4p1GEsoYPd
UNmKg2X7OP6lsFmjcimS2272mvlUGMa+hhdxLTVBFHJq3NL3uk1iaoKOekg58ef1
ittiFAbJuo6Qbmd3wjGWnqxQrmGDaTdfnRn3TemZeYS08RKftPHQqoUkuZkbaGXN
3YLiyPYoLUIyZqIYCqiiO7LoXuOMumVNRTWnZG75aRhqt/lZ3IH0wnr1m78pge0D
XLsCUG7Jt9pfhL/yGBbQV1U7+FPAoOH4M0r3kruVG28ozkvp5ACgrGH4BuEVuhog
Dc0ppQPgWnO8evL5VUbP9oQPJ/Du7J2kHcJWChwS9mG0TgZ0SaBq8MXqAwLlJo/0
wC7CCX8U3iOqAokPBEF0/WnO7W1pria8i+F1FZHoJ7ebTAc+/6Q8WTPHoRijSJix
g1VcraCas6Z/irMGjO1MAOc7c7OdN88A5vCPr/wU6ONs4yU627/X72wjyaTrETUR
Slhd/7Y7Bum/3nyXwa5YcUURu+WBHkGTQae8LPUPYNSJY2rgpw+5MqkiWB2E/PpY
++wp2CVUWd6NqJ77tfFFpssO7fkiJ4p+C506AOpmv4EL8dKClc6rK1n3zn2Zh1eN
CygTat+rQOocFSKaFLCZn8KLWdDwHZ+/uxt385FYl8w5M8fYzwTUq47ERFurv6ho
xlVx0wvjYdGEd3hfg6GEsFOGSbegobdT0CRJr+oryrwIlT7EfsdlPBjEVqeGtf+T
5hTH/cIIgy6XhvoBHWcL/AS/+N5OfqFMKJXtgL1dj5N/XsdOn7bhxnN2Yi1Dj8RU
SxBeq7XLtd7MtLTNSSjfywvuaBAlnvL5cYyjGS9LbgieAKFAKYt9n2c9I9pZZKkC
bS8NzoG3DZbsho8VwA9rkqMV4b9pssFrKvKlRtnttFVYXyk8YpgZm47kuifBggww
fURpLlXVuMIGgNVHVBvB33cpzShUa+fEpWaZT3cz1YZwGUgd2IWSMBuNUnebNSeI
XwjfneMFd1gEKw2RHRPtb7uKz+i7OA/CHdu0cWz2VcIq7CjwUJMT+lSOV6aE2dG+
kIPkI/sifS1AD2KEWrc1Hp1MK+MDIn4uzYrp8zNx8MGnOuSrmopIq6CnrJERoUss
VI46elmQodE/Se4O2FY9hHaqPD/w0gAYW/QewxZKcHGW0SgeunbgPupzWPX6odYv
6Y1h8vZebUzQCavNdSOU2Ns8o7pvp6rG5OyQLFxOULerLxva2CXWlLxk2obPFVEF
eb3Tl1zyJ5agt8NEG//J3tYDXzLIzWYu2cUnPTiICwuP0OHaoE4GQYDP+HTiOpFK
tyHaAqCmWS9WaWnK4+1D+PG6tvSUpzakDWu8+K1Y+tc3Tj928/uIDGjfBuq0+5de
1j6hLM4SuOhze0Giayo2QkKsoGPObYhZuu68A73C6Hrf8P3b0G4LdQAO2rCPnCi1
Jlq1gbQ2gy4whBlFsxHYam4K+kEt33oe0dA9IRGlcX4lIAJKx9vYg7yb2dfIr+ZH
1JOcxEpT26P/riEuq2Rlu4zov5Yl0N5jsFsG3LlZNnsR3FJEJGxGwQIbvI7KHF5w
W6PfUpG99CE40ba2Ck2ewef7fSPA+WAGoUucmDKjTWC7yjVU/Arvcr/+ws78xEGQ
Tx9UNYeaAjagP8SZdpMMtitUxP+OqcJLwLZRMmN2kJRkbTinMyFKXW/+4XSNGYZV
2vd8drVje3D/mM8l4W4LY6zA8G2n+G3uq8Dv4kimmQZzNLLmndf0t+3Q5fRKo5E+
/n249NHCFXG3ypYo5jlSPwcRKfzD/maqXb/0q+LhVwdY9OttM6oUDnIZXHBv1HHG
ftcZTbd5o7/yqBE+7ibES+vYFcG0Y6rqxp5ppuDBBsZ7N12UUw3PWns3DJUTklQQ
CTU6J67LU0/8/NK074fC0dcehmLBhV1Xvi0bi2J6XVBWbX/UWcFY8F/9gHlLQFP0
/ouN9Ib+EftW7H+BzPNTEKs7jzhX7x8UP7ceyoB13liAf0/AqOxTnPpzV6KpRYNm
J7WhdrRzOyirv4kuWChByyiKNDj939eLcvfLndtJ8j/Zx3LqgGfmP1HdvafWJcP8
FBd5WybSHFLOErwJgThvOBefGhlCKnDcNFnncpX9U9SlTPj8VPwZh5JyHlx/fk4o
LXuJ/r3k/0gThY6fnctjqXFSuuf+9x6wrYvz82ZtJfxNFFpdRaTYZf6HCCq5aR50
BP00kFim7K2MXxri45bm8QDvDfEwYSMe7zczGwP4hD/1gkEMzFXdby+nax56UENy
NigL00+a42fYSNRNSXlZwO8AG7rqj2U5C3cEQUu9DyMfPxNSAK6ItlluIBFc5V70
Gu+bsaodZo3gME387C5ZRNtOgj5PNDyUPm6dNwdfP3GN05O9XZOm/fIQxSSrpcPz
Bxd5jnJ7wEWws4Li4Cq57JwUoKlL92FvFxwJYbA5iZtl2tMX/G9eTEjWioQiVMKq
38mXroJA5Td5q1Q+8PgWNaPoBNxEvlt7Rk8RHIeK65i9QtsGqEmh6DktVZi/GRwO
L6kIPxW3UJhP3kf8JIO+BJT5hKBFNt2mXzdm2qlsFNOij9Ia1+I8h/Bmik0px6YU
+8rTWCocJ5r43l1ZO40CzWi3wPdEqOwS80E6l87B4SF6/pUg158WomOkmeO8xRRo
764Ohec7e6xhZqsISokjXO7MEGGXoC0/nJMwk4+DGWeJr48A5sKl3zLtVxIVd/ew
4OGvSmz9hlFOszIKli/BQEXEe+V+Bf0C6aV3gIZ3noLAGsKtBrsYMQ9Ys2yKRJIA
4ppRMUJCukhClEviT7W4MmRIGq0VdWt6/W5Boz5yR1QMweYtCBgIaqa+TecRNDNV
OZbUK2S3/gmrdWdKdb9QqfEPWakf/TDRWGuzIYcnNDWfu3zoZBRi+rd8iW2DhVVe
g9EKVEm1YuJYvKci9DV2QNLGOgHb1AJAYOWvB4wPg+WMco8JdzjP4F2HrArLtx0N
XutXX8uAF9jDQWtM0AMPBDo98uSOviMAjEBljCaCjtG2GmgD70bgJfDY69KHUifq
sNBJWPcVQB0jEQ4eezlpHunAQkwXUy2NDGMn3G0285wP00EU4gkhw30gJmbNYLtp
6I0DsgQpCxbBivaU+bvB/UdSdDW4Z9lgiGN1Km7TS7tn83MfVbeRRLqcJqIZ+uFn
JvA3UY0UrqHf+cPq5Dr3TJTzPCdqViXaXfDUyGa6ovPBKd0TeMjf0C6HhuQyRfeE
QfZYTt7xMm5uHBYvVgIRV6cDv52N12hB0Yqx+pXm2nydaF/pMtiItVCtpWhjpcU4
ft1OMp7OqQkoyt4cWOnva1Tq8SvEUPnkArIAJ3fTpM/vaSk/SEmUTWD/fkTvMDf+
eEVtzpgtX7/xUF+gxp2rm5amYS/DuZl9rkcXepq7w7ZwnZ1nrXNccTSCySbDcy8R
L+zmDwf1ybY52Is8eJhPpIg4g5sF3xBbNhHZ1RkYmNIsScUM8JrkRiRcGK1E4kpg
I/UUiOKBBOy+V3CpGKC5rs5uvoeoECTAxthxB9/vuLwoCpW1vlyL4KJEwWWOQZop
yK9O6566k9he17DY4nwWQza+PXmEFnZdso3XiKDkPPVJdTupmkvplwyNoj9AKiAr
PNWTvZNkswp3+0X/b4c6oqE5JELaNv2eUM/VRhYmApyAOy21i1EiqZmN8TeU2JVh
lDfE5Qi4h42BK0HOA9KSOSF3LnIQvH53wkm23Xau2q0FgMGldk0+0PHmYq/Y5tfH
wfFyghjcZvFxIj8G43NVO/YGH+RXcJNkpPNxAOQk1yMEvVpMbQ0pt77W85PpGNSp
IFf6pu4ljux1sYoWYkXLKH6lziuPu6aOI74D1Jv4sBZ6VLBdV9D6u8OfkHgiwG6v
8iRpXaSFhrb62OGF9qyko4L4AZrtCijD3aUOu4LtmYCTNcoSKxISUuEtVaf6xQbU
SrJmob7WXuiuX9QKGlVU+ToF6AZdIO7WEEcLGEE4lNq0SSj2glrTiqinK9wxMG+M
9eTcemkJOgP4wO/gRAZZ3oZXVJ9GScGI/DOMqqc9CRusnxMriju2yDx6w8hr3upv
iYlObvbQROdHYvvZozXjKBQeQiBuRZ2s9cQZxbFluVhjZ1z96rcpnPckovzeDAIL
qzlgK4s1qbZwufE63oWLLtlcyx0DFHGmFQxZR202pbv+Cju+37E6B0RhZh17KFp4
I6Gve7xPuDnu2jkImqxgxXlHC/FLA4yV4SImYAvI2fvVo1+PwRVHcHd4WkTER1ss
snF9W03G91Q4WUIhugpZU6/TveSHlOednLZrhGRTPkeJUDJz/QJ2pHuM7tChw3Lf
Z651hcSIHS83XG0q0lQgefJzOosUh76SFlr25pXplOO7rwNv0sVWoOouhFLRUaJ9
QQrPsi3Rxw5EWeTLJhz/FegIWR1+vSXuiRwh7IR3MzAfbiCqUS7iZR9ZDQyI6dbk
xhuUWjgbWNyhzKxAZW7kGbSMYchUdgtsBlsxvrbapK5QiNsHSihjlmsOraIbkg0P
zw2zpj7Lb+MbM50k8bTJre0JFAAaFL9/k+0Q3od10a47ykF7w0O1x3q51ukVTWsk
M/ha8T8yGMdVl8LzLHZtbiuMTr9lzAi63OxmQMxTaMw9jXikesA3C6Z4ljxl6hVj
daZjuIUqI1BChK85v2jr0XQLo1NhdxfRhr+kKyPqZ9+ikhyEHF2Cu4llQW+UGurx
0YgLp4VeCTrwCNNNe1swj+dJKdnVrMlUnX8xHbQ1IWBlWM0h/1Vs3zKz5fKFC5Ed
CGjavDUkMTDIdFbAgPVqoZjVzP0VSci7LaQcvGB41cHAiU8juLmuA8JZfg8VKdMT
44DOiRitxLm5uhpIRHXI+2gZzD0TWrPx2Fe9djjVMTGzm352V+RGDAdzTEXNf2yi
p9RRs3YwP9jBP/bDrK8qVEQs9Jo9PdMmb/YAVtxbRX5Fu2MeiP1WmpJKAAVo3JoL
3yf9sJFysTKpG5AYpQG6QhV/UZ3pbS0fQDLHHUtMm7mSlafHE+yrwwdbjrBLxF45
MhaPKlmnIA8/Gst8OECkAmtFb3lwIBem36JR9nii6miER2UpeBPwtpewMWKF/0WC
cXK2UCJINgQfuTumIz05XL9DK0gk8Wg9H5BbF63m27Pr62KkshgA1h3GKby6bPPu
R4R50RxH/khUaR5R0Y06mkzDSuuQGkBWP7/iWWQCSitiVIwbCumxuvi08/cD/g82
8Qf40/yxM9doMFFx6UDq1Gpl9u8QfhMHUjKR127eAeSsXAC5uS0P+JbITJC9ka9Z
Pod6OKg/qSJ+AKWuOvzYBEIAkfKUmL3hR1/V8PDPESk038UZG/H9REB8htOQYsib
mCQUjGvArRYWx0RAaAcDeorzPDSkYxVryvvQvDiY1NIz0TyshJKDwih+Kpnjo2j0
1XCiuf9kfnwhaIrBIVJffeM/h3aID0aJA3KDFpuWUAZu5KsoW6qMaExFLWrdWv3y
f1rOWWltNxXTjUmOr3BbBBiVBFlpS435UB9sW9nIn7kqWkj7gx5lqBo8PRl4DqwH
lDqipaGPWjJSkxGQmdK2uwHfFd26WX4zcHgtedkcu3SIwf/+jnYyibKYtO9QWqNi
vewNR/H81zUeAv06A11v3RhBKQTScpT1CCHJsqCI4w0Udojf6Etx8QnMgIHWs08X
OD9YzlwFJe9CLYgYMhN8rlO5WZzSivKSj8PkowefJGcbeH3+pLtlg8r/UgToH9Xu
Lo6mL3CwvRVtvtCYFNBF+JHm0+ws73d/me0Ms/+DnRv/nLOlqKZmU2HdCjG4Q3RU
gDaX7HCwkPFtedalJDweGSkPyn7tDHprXFPjtiQQdl5T75AAnRb8fvCXPrc63fry
yGc5tWDrEN8BGQQy6w4n9fp3q9RGkFlPBs6zb6tPJglLh4pvYOJfYBzX13YeiAdz
1+sDM/lmBxezgWa8QeL33ItWrd/6iOFsimjcphCXU6c5NShmMKgntkpBaCFYRTiC
+QxPrnbJXICsddbZlbfQJgRFbREBj5yLHTRrNdWnoT+fv1XTbr73Eh9TeD9DmLJ4
q2xqPL0RHH8+rxXTpOCPQmCn24KzfZnXf5XDIgHL1mX0uArB8jWdvauuzkv8xoVM
XSEdppq9f2BcIRPZRqlSlpFtO3GC31hDOJrDk0j9jwzFNbMtcqcBqUENbFEB/aQa
mCzqW1IX3YRvUww0MNAvRkIB2G4Z5w6YjUJPvJ0Js6jxnPErJ/qGUJj+LmenC15A
nN/59WDG/yHpeh8gwGqxtCjS8/YoeOgut/bJNrGY4bJk3S4qrRzm7IuOzT3XwPwF
FPmqQnx1dfCIxajTUNyol8bFGcHae2KqpcY1hfScRTfL2ZqgYthQxwuqNteimSzS
H3SwUsZO5SWQjh65J5jrGMCbSskxwOiIQ7No00njRSW4jASgSby46CGU2RNDoT1l
RnpAmaChzmynNELyEDdLGnoVrEQpVKGYt+BWhHi7L7+Bm9JPimGVgmvWXf3kYf1n
wOapHR/akpZMHmbx4xfwxUFXgdbBob7eGkY10ncG2LySct/oPTisl45XPH/7IfVU
9fJ3dWWP2cL3Ekowd0b2/saO3bYB9WWvnuqkw57iBtxmYJPsasWsQAzOEn1+mTKL
uqAOEdnheOEkUSNLF0cQ00AnKsQOdMB/OtwVMiurLRzM9bnZL3KrsN3MhJdwsaVV
jyhGg38fokYEKqDXysr/9PjLAWj6Ao74oNeIP3rX0+TOYJE14KmWiL/ADsy9XdDn
cc6GQFDslzpCjUmUJLw65in2LNFPrQ5grrG3CflHCdYgcPvHDB9vS6AXMJ7ceUKz
tRYqFvhzZGj0CIJMx60+B3mmQsuLKyFgQr/ZleWOSmTTsHduFCO/jZHvA3yl3lSu
ngub729Otu+9OcjJJBMTDZmngpO3raBLN2XDIrAWisxQvaTNSA5s0DLGE4UUbr0b
+85aP+i9vDaAvM3AGpWQE0EcFRONqGd02/gG6kPYh8z2VHwE9CwwVJUG5ylPSw/3
RYpzfGLu6cOsy0pv6ODv1/kTDLVOMTE9S85G9GXQkXKLBbsadUv0JbmxfVfHssow
cGMi9xRfKSufOkS/DfxXTd9Ro/EiMh3jQZoVcV3O7R5NIPLyrmYmS3EaFOOTMfNN
0+s9WpWOrywJhCGTNr+OrOrmosWzEimB7y6WHQBJcRnI8LFoTwr84bbMj5Q2+XS1
XTeEep+hnxPbXWkADRgSuPUun0WDdfLZVeHl34RoUmDFXedZdZoS0BQK9Kk7CNSc
eAqVAgkWROqQat46/6bYaVoFbrYVwEtuLjE0ld9rhqLYLKDoGLUmYie7ksVncGwo
cOvrbCRg6V1iQhRLjIGGPJPJ5jvG1sngNFgm6QnNbSuJeSUGV2KUzyV2HDd85f7P
R/NfdKA5tGGLP++lfnpcfQ5aurl8eFo1E3YiFF9gHv7QfSJyP6rPxnhMaFOgjCdK
eh+/F3M7ECYksYO1yjqqedQPrm2oIgwrNeYKv7kxH4a87ip+JSLDpkc2bYNx1Sut
ujJ6EjwNGzg/5ZCewGQ9isTMykKYs8q7o9bzspL2OuNlQIsYwv+bGhvQqxk6Cx/K
VaUc6/QTcYpshxW7cKPm1ZqBUq429UePZ89X0xQR+aYC085siQ+fzJAm8/+DsNBv
NGRoNX574t2yb4XeDzc+VE443Z70rQ1ZIrmA/H6dLrKEEDfTDZTNUNfRZfDZzOn1
H7kPwbiW0b0RBNywRXfIUmNtZInlyOUAYmk0KUhhx5fSvDTsDetsE2rkqwrKzVPY
ihyd07Mr/aVVI6ljO0IiFvfV2Sn8jJZ0IIsCfZRZxhS++y0HWhn4XJx68nVVOFhV
NJqroSo9WVNcPPWOgTV13nD+pZPBpU+50lNM1MOnN48+O3fABZvn7aNmkL9OV3a2
PF4qlYm1Q+tfu/dXPYjeEAX3H1F5rGZdYkADFthT3JQWnJVWzkjD/10X3BBKMMxx
H6Qs20jV3FFUp3rB69d9BD2WuHGTaLsdRj/+dmQVHrQzCBrTy+exzCMPhp/mNClK
Tu5WjjvrizzQQ9tNHfUVqFNyMaHZ6/tIBapwZPcgdNfG4qR10Lm5UgORk0QY2spM
Z2NIKa7D8trL3kdEVwza8Skys6d1e+LHOalthmeCRDd93Vew84Q+ltbMbQdDSrBS
hbnsnpA5oOyt2sb9JXD7qlR/g/TJl3QaQDa/PzbS2Wg+21KdQX/5kh+2yn95RTjb
rqC0RILY9k5H1RzSVe64d+llIxwxGOd3YBt1aRgUtz1f6L4uoEumlcqyGkm2d2PK
eYsctiTtCq874oiKdBpQuDKLPQOQx4C5D/LieRIYaFwsM4NPYkiOA8jA3Wy5K5Ro
6382EptcosVhBt00m+u64mzSI9T+nrdUFHVGkSjFSQwEYfhnkBL1AVx5nlKzVH1c
rZavkJ1vM/ueaxAR/ohNVXY0s/LA0SqY0w/kh0ne6RcRUA3EJOv3JBRlWUQK74LR
cRCBB8lzAhqOx1lvBuSOr/GWmR79eTBubRcrq4sBRoDoVQqTCl5mqrPEfI8uF0l5
2vvG0Sq/muIVWcoRe7fHtdqYS0TGIrEtUgOv/1eiL4OLK2pm5tQ3NgC7iTV5QWt5
L3WosTWkdszoxd4GEihkbxt4K+g0Y0WNxK7/QyiIMwk9yTCI3bYe5eLugdqNhHZt
U3S1gxNs23cCf3yLBfeDWNv2wEUkdso6cC40kr00fibyIRVNx1qHuUwZD7mqxKdd
zn7gHvPYmTNjnVVPtpp3o9T21GatBZsT3b8ypSHj6pdI3hizKK9fmSceZeUiN17N
HgIHn1TUDbtjZQqr+bri23+JCY8RmrDDElG0FSpkNx0nAeBJBuJFb6TKK2Dwr6pr
fYgAbNsg4TVt/M0KZPpOTzA5RVhDHTy2DsBHgjFjm874QU25V1LQSFOV8X8wHnSW
1r3IZ1bIi6B4FKZaCWHo7WDfxTl8AYKmM29neqK04U22MM4mC4G3BZ46+s/WzYUp
/TNK3IEjtrQnNobCH0r2qde1GsLcTy2XxcbtI/EGZLDweULd1ixFlPllF4V6IxBl
aW5s/UqGWtEVEtLYIWQ1YubjW+7SBNeVenijwRnkBkcBWo39PnJ4yJzbFgmgdfnV
/3s+UrMhY4K7EjogbugIEbqlDEhmO29cfHWEd1VM9zEm3ULsQL0aOB+kP6k88uCK
jlmp0mmBYOK4fmMupY7HNAZqlEu2tIsXjNx8jePlkOyPST257Q928hgZC//FtiFm
4laJs5l7iwN8YVyAtVpgj/uGc8bidI8nrJmuvfrW/e/GGuAgtSO+JJ41ZHejA/il
ubwqM+Y0AO6A7RtIiI3GgFYaXC/zQICloGC/sozYVRoLiS3rLrBThl3RbFlyUyvC
g3V6mPcfkoxOWi4cCLPmtJjI2gFMK+Y+caV9YvynZxppd5lnKhxRCN3R/NSnGaYd
rnLQTls5aGT4UiV7Xeyai9BxuA59aGfnsb7voFZoF2/tbo8kTGeEp+yHY5wsWJ9p
Td0VJYawVtbTs3SuTNa+oPKcRu4qtktPLuZ3wdDuPKZ1aLrHpuI7hWwumT5JKzpq
X7B/hPVMUl+5QXLpUlu3a73Qr11QttCuKd3Xnp/8dnPW101gNQ77OcD4zWq9kFHk
3r1kVAeMVsb/lLCfVTRHRzDNk2/sp4I4UO8mp8nulcDA6gloEE/uqAMoK2n4ZULx
vIdhV/AhaPYVwdY2RJqg2V+CLyTc0gceoKUA2yF8AxQ3ruaNNTgwu4yYB7gNPgdf
joRK0q+yAWiPWeq9dMlTKLLB4lLOwsgJLgorLKtHYGh+keoIaZQyB5WQEzZZattH
sLtASZDuQ1owjpzqFubHcbAk+qgmLNI7JPu/XatHSkj67iJh3fRFPWmixBhpls0y
urkdGPtfN0IiEu10TrbxhQhc/gjgRjT/K83eNA8SmZXL7DyIFYHfgJ7TJPndRhdD
tYXZDsyrKQWjMbiQP11y+2hwRDejrBoAvHMT49MrzrGmhrhHiKcXgFfa9W5FHF4h
LaJZdbCnUI0s6D2jdQaC7gSumgjh/kFFBh+Fk/cqLSLc6aWIkKr7woxfA07Qk0gg
8q8zq+zJFw/9ZecmYnG8LlRbtUzvbnFE1HjhefcWUIQK6GP4ciIVGn/nWCg0f6fE
OvHDwTrGlXQuWCe5zz8dkEUywtqD2R0TacTjBmSVuMTd8tXcmaLvo89zVtRfZGRH
0KL7P3t7FImIWNUqntyUi+mpr27LlzwweYp8+FBOKx83PtoKdObQLiZs641RH9qe
6CX8BWXsrwu6pioy8hfO3kTCdl0CGmAp6N4qRC70mdu2R899WHbtXJbkIJD6oCB/
28qgololMexY7SuTvq3q/9M0tn9FZGQYNaSSTBP5s49a/Y1qxAeZx3HIs4KKYXxA
pOgpZdrqqyZGjXifoXhExP40wG4hMXK52KvfoNMXdACD3Uv0IMuiihIAVyQ4iamr
yOcLNaFUYU1NAf3BmIamEf0EEYAig/ioUCDH2uPYq8bve2dyWgx40MV4XHkwV//j
PNqu/I5aQRQLspj06svCaZgdMlMaGwHHRjbDQe3wlRVijdkKrDsGwJunqRJFEKXf
GnLa5Do3N7+4ud8LTMTs4/pIPIcNEhSpVX2kv6TnQoedBD+30DfkUtCCskbC/Q2f
yABBxz/YPZVosfWOzN984/bkRJFNnal1BZMFcCSybTSqL+m4zXwKLqSBhkvTjg7l
W+HFfwn7dG/F2cQkbpFc9VM/HvABTiHYDlOcIgrkHCS3uRNXyCZBrZKS4a4gQvxY
1DMdQFyXY1yqoRauLXedQZgEv7YJcEY2x+y2ScbMDDrwV+g4JCDppTh3F0m6IQY4
QeGiZ6ZvSoPDzpCZlnUmtql7R6wD0VZu6muy8axWZLgzmHZ4YOysNZa8EUhhAhnN
gvA0e4pTul7JKpq6UTBjVR/V+OasR4A2A+mvDDFGABzKNjXUfu3wN4Y7YKOQUx78
BLOk7acNPGw9JjV4E8JGVhM/hcKRxsK0vwT08/ebZ6PL/OVMTr2/li/1hhwnSN8U
crp99Dflfz1/NtyiiegVVxygPdvKfFRtXBshRZXAqgj0EXyknxopPJFYL/KulsR2
R/oEXeJtN5EsZnFrWQ+F8kLExZPadOo3in8Dv8IyV3THYNWikbuadIS46lpSEfVm
s7zhdrgk9SUNFeH1cV6KMoDRA8E/4wWKxHd16PRZ9YVbw+EbR96YLjB4+F69KyZC
sJB+RdZzuWFHgicAheG75KSuplgP0jHaP7vKJPiwmeTo9GWUPLC8CKof98B2Y8jV
VKCFgUrFhBn3qkyNe5B6KifvUyOuf1jLS7ADq3Nny2zIYb2Ezb+/yFIoPiceOtks
YplWvwF+4DYzb7mm2IF7QmLKqmXTlViS2gEG4/uai6/KbZE9v7l2CW3Mle4153IM
qMvOBZBSgtqorU94mE8oa6fUOt3MDgFrxQP1qwf0BUJU6tiQviWJid0zgXwoNVOA
c6x0QXh2+5ydkcPSpKaRZ39fpdZ+fJzLeX7cIn0Pfb8RM3ofppYyotu+r0bK3spg
PyYrx+8bonre+qy56VSfss/6R6dH2Y4VYjpfeDquyIQUjoQFIJCMLIKLw21VCvzY
0IioB3akBYP2gVlkgC7Jur71mwhoXQAo6IwTg91lRj37ncMeuj3lxGvNb5B8w7/n
wLPUmcs0hgk0TnrFjlAIhcKdSDkpwCXmhe/1Cpb/gM9SR7kGnSMamGzikwcN7aS9
AMmQ/DJ7nknwjmkqNyKCqmFlgiGt0GMGxkGPOlpsuzLAkQ+Cid7Mq4G/KLXhXtEj
RoRkbEMQOzGoa/lNTKFsUUUfgvKgHGJOgWcj11MuOsDx31tVdjUuYeXOboKa9hRI
hdJvARZkRCq+qh3e8wJ5609BsgcJmqbimRDdODdGl/pMYRFnXa3VowMSC7Hkn5Oj
pPdSbxUgBncXlR8cWh4tzhG1hPFtxEsc+Oqu9CMBN8B8egD4Y2w6ykUWH1rUc3JL
KvYn0MsS/lxyUptnzZbJFOHexzkvC2Y65TLIZCv4Yj3wK8+Zwk8jw7l+4oR6/5mo
s1qCL/JYTxkQW7wu+BC8imBrnijuPVlKH9JqFf5hVyWH8b7V6z4EnMp4S+9ufUKU
YsZ+JRtjcUhyzCIwPdHq7+HqLu+05wKo8rwFgG+RsGXNJ9Xerr2gPJQWx46dXO5q
EAXztdbB/tFeiskhPlBY765BBJCBSvXT0e5yLs0/xR3hod1uy9ifULojNnn1wDNp
jXNSroyklwFvQOZ5/5z4FTzCe2F8LhfoisVj9F3in9KMh6pPrWYbyCcip2BiqGcC
G0MZTT6gWe+5VMbDM66jqgrq7OlSAtaJqaNZvSMQb10zTd7ZjC7lNAnBpvyGpltM
a673VVQ2/RfWfkKX9cn/EWQ9NMq5RPyiLbWeUXmGlsY+TmrDbRhZBo8UhX1dL7pi
EBvmBpYIAbad+ur+9v/MGXbtZQa1FTTQc9Z7UcBAuWw0RfZGMdOgaVwUMNigIjip
V05eC3wMAWrVnoxT702KXuysJDai/k+dLucPokbG1WupdvG1l0VUbmSdnGEjmNNo
kTAPAtiLy25BlCDVjTGNTIvrvCWb6g8zxOG/zU6EhvPs5m1dxm5IpGamJp6wzYex
bHkY+V0ItAv76D7vzoECrC0VQqbG6Q3UwLAyjWgnNo35KZNoQoXAC9vO1lEuOZoW
w2I7jJtzZeR31OvfhutEikBpJpZGY3Hgn4xlK1HdfdpfMM8unaXIGU3D4/q4zMWJ
+DMUGIAsoQXAwJ3y+baSiuB9sN21bKqeWc9YDZhejXIv0W1i1BvWBmGZ2rMSGVPX
aWFAw5Bi9VpArpG+3jGSNeZBDa/ZD7vyYa7eqP7cGCvbrSw0x4tKix/ECZPYJmIm
YTZxfILs3n6JV11Spk1kCqxAQ1cPjOw7rM3qmGe/7ss3jbJaZA9SaIUjR/NiRi3U
91gR61H828YKT6zIqnJce4RpBwdJWCDPpycSi2xvqsr7uaClMGXkDgFE88PcypGx
/eFENhtPIlOyQO1scsyMR9jXSXbIulm8cOwHYd0nZp+e0hH7DQsxJe6T5CyqPA62
gIa0lQO7n0lTJBWIRWOz3cVFu7JXd56Sr16eZCKG+jnvLXlE0DjkFQcciupVO8CB
PVm4zCzHzsU5bVi6YOB+9UTkn+1riYnsPCLOFJptnUfmv32eTTfoN+eZFWOJHwsQ
NmjkHfQrY7HgW9V4Fxe292LvfmdbbMb3PxkDNrJPPrpjiCCE8j4/4Ja55xbZvLRJ
TYZ+OvlgtF9amEae7ufTBo/IpZZh8YBRLB+5YbfvUjMNhKmY8CafxTAVO6mH/Zl5
30rySqK9iT96Th7hfX9wjM/5eBDSLU/7V2BAcsADwaW9OLL45PhbUf47D9YNKMq6
7taZBJ5V2F1nPYFhSU0NiaOKeYsQ/zCLlfJfObOp9veCIIyMihgiNcIOByJLMAIK
ILgp5EkAmeOvMHdo/t4PHMtDpQPqdetvFEK3J1dagIjgzcSMZDlSKM70Z0Bhgzha
4ujcCemhKZoQgwgIbv5YG9K9TYYIkdgd/MEXpAw0gxuG3qFzmSAEmoRWB6X9Tq/8
qqQhVON1d24FfiO8mzZ1AOGIBkBm92yZBukrD/MDymvxlTf9NS6VPXMmKhUxnu1C
VxusYJVkkw3B58pOKrWoxLKOEFh53zy8uSOCK1+/iiJo0242jVECgu3kZR0cSNdC
N/xuN8eDtqvvPz8BoSnIgR0y2QYuKnxLpV1Q3Ynr33T844XYWoc5uvoiZwEO26Vd
yddysa/PfiCZCzKLpvU8m7gDu/WAvGX3mJE3URk/FLGwiezPzDQmbLSC+K3Ya2Qg
U1Eb1E6IyFxnSNdeRxYq07upC19OXcCbV9SsW40zy7HMTQ3I514rebyAwcLyl0Ih
Hi60nzzRaDyBlUCQt/VxRubZbnaQVWfZAXc9FELKGrOOyNC4QjgAfCyygsQLTYSd
gpMteghU/vcSe+0kltWfiyovkLTBNLHztb6R+j700x56fr6bp/zdyIMWt4RQyCFN
ABHnqwhZRpeSaY+T0rt17Hx0goZJE4uZ94ULHu5SyM29yImwOI6Q2zjEGu9hLFuy
+Md4TTf7G3EUq0b5M/DFAyBDMRG5RMXYe+R0HtygLjdP3Snw3dy1VpCt+RJlE4vY
+lqonJumQspLGibcsZH3802LLY6welj3AFIoN+l2B/S/Yd6z9vYymGzsaU/qtiB2
+jTBAZD+us2HGKrBYqjmc6N2R2xaNb/+F2vwEMWxAAhI9q7Q6KyTPaiVqOntZEVN
S6IauZ15SO0gnBD6SVCMbg6h+O4+6xsBIgDf5IICxVTSKxtmG0RJ99Rl/U0zHZS1
69EMdz2xN3QDtTHDlREyv5E5FQJ1uLoJHBFMI+NAXuKBTfnTseYn97RQT8GWSXx1
Yo4DWzDdrDHNemDwat5H3QtnxL7FkFN4/x66Xa8SXTE1apvn5nwAsXlljg39u0dD
Bq6bPDFirOG+ZQz93PqvufGe0yZ95PkVBkewuNAnOkK3UMKCpQTbv7lnyu3SfSR0
yjIlGQgV0+ga+Zkngkirfc7iAIqADAybqtacA2K+t3WqnJtKaFplHGrjs3S/Q3nw
FI3rCul9X3i2tJ9rWriPm9BGB2YTzmkChRJGCZqR4u0ai2vcK/YQyAJIhmaV5shS
xRBBzeJd8oXO05wefqHpR+zLLQU+xsI2g0pr3m/RzH0WxMQn0axsJMAxGKpKfhz2
UHOEGYRpPhmv4Bcyx1SwfxhHej7OXFXgA+XObRT4BamVUF59snjejd4oU3k2IcjG
BAtk+v5GMajRew/vlu0bbqPPK9FvCvovQAts1lbiiUdN/YsLfQNeNdmAc5KvyAcx
3/F3QtcGAgdTjbLlUXwHL6CEOO1CcoV7WLru+2lA0SbGJhfEAVQkv7tlk6ngGyeM
uzhA2WOsa8i16igatXCq40zMLJwlzZaMAjxNjiR4dnd3Kw5slvZA5HXwhi1eNvkN
/6WDP3ne7hSYhZSZrhuBTCTqJYFSCHIcEWA8oJ8SFBVzr34tlgR9KoIKEFfos+zk
UngtbskSYC8A/OMmChqQywJtGJN+4BGv9CmP/MnMVs5s9SAV2C6KEfGS6VfjVdUc
QFlgvU6tGElNguhJ6BpUGQTJ/qdDppXkkvQiDr4eJqMBgpQZHzleACWuQdYqLYY9
q4zEezG42cRqoQaryZZ8r2wmMU5OpEFOQe5IwUXn016m9eNds8PrBeiUHsiZMrNA
PFCIVsg7IykuHx8ymB9PuuSJ2gO3h5gM/aSoOB/whR0QFWzEZ5RYhgaaVECG0QAD
iUNhFhJNZyjeY7Uj69dQyna3FGVGxuMZ7r5JolaJ53NZnZt7c0i9F8JZBnZTSQFI
R/fg98BpfCCPo4O7kJJLl6mwlbpRLfaaHJUm4l/yokwIPJ17xEXMcsjJrnoMJY+3
jU9JzAISR+o0kPCQaA2cZrQ/rzegyk7MMgo43RoMD+Zrfaiad99ZquRYmIAp4pmk
XO6bloBEaTWf5dLQhy2qFx6iiVfu0oujZbM2ROcU8ohnT5ADu97mE9Jr7q3ztg4q
z8tHRnsYZ9BLJ0ST5QNhK7abOl6niyZ7etp145yANWewZIJurbKjmId+iI7dJCeb
l9f78R4zwJcc7RAkY4wKcN4h2TisDVT5d+qzrpL9Pi0A7kT6KjxHRifmwoBDRxkz
DTT+v3tHTVmukKurdEdyQW+RTxPIJSBIahyzocAyn0C9DlmvfQs8xy5/d6EzG3SQ
i7cRbgc7XJ3+yTTyga4HWJHk74QeaC6J//pK+iQ4OlbkVpzPtAGiRv+Uah+aKHoP
JBb6BIPFUM3dGHLKSbBD9QaGHIGRzVOyZzu3pOWFehUn9eiV/6WiJGKBKSpWmZMj
lvjgdWPDtJNj7W7CONnR3iEFa0cpYb0ZSIU3+IJjUnftBKd/zBTFzq36UiaMuN00
H1UVU8JgtX7CBLtRymeXFgSxxneFkSYj5LGcI7N6vR2rCkDgPPFVLFntNy0xSEkk
Z3uM50lRBW3ssqKC6FrupeIOKU0Yt4CI6XEcoC4LU/FqvSGaJQUb4Nvx+VgtNdoQ
2+Dfs3cprKwZv+GumxYsOBfQpOa0JxAFAJcxIx50xTmFd7UhNFMLACkJhnNEwZ6z
gMX1/eCSbdrN2MIpj9pmkZ45EJsdMp8NmFBYPGtQZCt2i3+ZgKXSV1lyzziNlqzd
DohK+55J9wO5qQePBNb0Dc0iDhxrJUkbC0pMCAxU31r7dgJFRBie0ok+w4DPs05d
k4+XrPeGSMOSpH/KXyxwWjAxeL98Oz3kqOAXTrDo2p46faZpMZMAjRkMAoG7JjT1
eejbZlNW/q6vpNLXjrgB96bR+XieV9bQ0OfA1qF5vFu6uSSsNvrBHLxSXc/6k2EL
DGfsqu6Ktyy70+qSR16HMtTGlu5mN35bkcNN81mUdIq/SZUqkwnmf4dSIPKaT86i
mtgIOyIptvAMWLLoDmSxudVtowAg4wJ8aTmFSziVmk6VxMH/xL5q4xs2rQ5SSnab
iPi96S0x05vY6nwTDYahVvaEFwB99NXdPP5V0vePS5Jjf6t/xLn7rGqk8myS82wl
fOrIYGw5TiVgXOrP6AwlLsH9EgI2vOt44q9EKOvolgWfeArUs1ekUEPaTfRqoDNg
Kp60pGr9nRBVKaX4y/zDAGzMyyYK1/vATNTyrpDoGnA4PS3zEdVYWMLj2iF4Jjbc
h1rGfYn5ggwe/3SUZgccyST2a7NS0biG5LGSmqboPlVLrEmdOHLOlK5jQqkjHfdt
mflZWCX+mkhwCToPShZT3xt7+TK/Xvam89+GOWk4ck0XsQrXJJXCM/S66Ar1Woef
V2M9Wt1lhuykoTJzW7t3dO46CS3wP02q5QfsCSX6EVkaHdE+3woUkd+HX6MiP1LV
ReWsWG9mhkbhbOdS2t2gSMpxq/BLHDhADgl+9621uG2tiMx0VFGFK30x9GPAL7sZ
bLUYeY9qwojywEBSC7Unps6BJv/7Dq7pCoFeteszP6doRZxR6sW0JihpPdwNL62p
TNExHLcfxiwTsDxWR/XHmdJ19Szgoa30YaP+b+JY4c8RjiQlaZDQ5t68LP/J8IfN
Hm9aBPUbQEYsmgLVDuap9CF2wy6XbcVDcAXagtrL2oCq3UiKLyH2yL+Ljh7N3fbX
wOEpYxjzmGEOQzT+yw4BVAcItx8Y9J7aFLoiV8y21GeEPlSFWeeKBlNf5UL2CqhR
8XCl0wOsa20YyHHgrJo5d+xs9fdS1sdBNSsQusC/d7S1FKfWxxy6EUYX6cT+MZdJ
o9eDkkFUANIJfITiAjxzZqnehp16DG1ZUAP4N0gyGaLKZs3YRnFpwqU9crjNdYjm
hlgiJo8Vku1OzMVCiRSUcsfad9a+Wyet1NaRzQ8wsLeZryRGnv7t7L4SkO8krzzh
A7DO7tP7K27i2c0Eb3dJIdK16xTplMChxxYEapwdFil9Yl91Lg2rZW0NDhWFGiEs
+CFTBE7AD5qpyrPrlqdaezhneIJrCbo48CjwjgdLMLSX/OSMU+TAveXwxlA4In6o
Ktxn2Gix/qwNQZX4t6px0pihG2ArDGapVaYP95mpQR59bG97btVanVW9VrPFmyYW
FfP4VTEkVGb838Pwc3RWqShxl0Ww+0/VejdHyzk2WwQ4KJUxFPLl6tgFJqKr4cgJ
+g2ILbQXbSp23xN9EQ3NkKZN426JMM05+B23jJLcHjZ/Z165+VbguWUxJZzTPRAx
lgBNbBYZzRn7TC76ee1yWIWC+oYYJD38KX8Tzjf2mUAcgUHcyeT//fgGyVDd4yf1
3yFsXbp8JoK7WuatPXNTJFuWmZBkHitVVXcECjpHZcoOiFMLjLm1m+5rObgLZQvz
eS12HQaC1K0ZUsYY9oXIFA2zpCMjBNj0hd7kw62YSB82LwVNpCUwfoGQHAqHcvL2
JEb2uEL5QIKE2TahEkWBXy/Btr4TCAOBw89/C3sUPLhOz8NiCdf2sQ/ReB81pyOQ
A4ggy5UJId0G6wXEaAx5Crk3FrUu7t+A/mGOr9G6IT/HMwxYwK+uzIjdONwPydP0
emZGBzyfKofxGo2fDYkDEr2tkTEIo711OMSpOA8lySW+fjr5d+h9a3o3K4mKroLK
R0+LBQnA9CyImPXNkCwvqbMGLj4z9TQZuGaNMOluW2yPzA5tHL3EVA/m17/+w39H
QCe0Ugt44d/ju3q1ztAPS68ns4NfqvT1KFaOZZj1fVMUhQRarePyb2I14NYFaMKO
A4Qrvc37lzNjEKgAqMlbgiMDR2nAVLLmEQI52ReYUeGskbkrYVj3VfUuLAkh+2xS
y29Xy12J8n10Jvp7p5/BRW4soCHixycGnHaBLIL5wKGUFAWCRKGkyRiw3rF3MKao
bjBqQ35tGgV4fHuUkZsWGvGCzDpZG0FnVbbstO4HbDO9r/Xm/KX5ZTnwdkTkB/ci
Qbq7YPsovr/+pxqJ2LJVe+q4pqu30Y1hJqL6CYfsnbiYEQqLq5umUVLF9f/7GFQ3
lvzVf0RXFMbSZambN8x4rg8FPoyXWEEo0yOLYNtS+8gP52W3UEL8cHbwLxtsAAo4
t5ZPbz/OyJX79+UGuLnnq1zG5pouGG39Z2lHMdFRwCJJwN5nkc+zWH8RjDIDGd4K
5kZt/AIqnW+aBoBLEOrMcoj9qXkj2qLG2T8HtHfNs9v/Xl6xYUtnvht0/lnXA/Yo
llIr4Z/YsfUIpz0VBJTCHVWTIQCMvpMbVWd8AHrWqZSc49B3q9Els7tODhe+QTh6
Pt2Ozl8bOtdvDQ3KxZMm6hOG/IDj7o7HfiZKwzxQnDIld/KKcI9ClFCmE6bYuEKF
t1Jtq8UItntUYFzln+8tmwg4UU75I3Slx2cNYFLoYjqTOWOEO8rfzHuS/awppcab
Kto5OsvqETN3qfKZZQD0H+TeATrK1aCMbO1cDQ0hzzi4gkQEugMbrsQgosDE9g1E
oStkEtbvdRTjQtcjTaVRdDP2Po2wp3O8v5WUGRI3UnhhH4CyPLTDx+LtlwowCZWC
eX8t9Lv6XxA5YxLLPJSQuURIBAZADY/6nBSPB/3oMNAsSRk11vQj03HxAyAPQWAH
3OE+XsDT0HLkirZ8CgpPcF1YghMcaoslmtD0OAhHTaBtjVPFiWOkzVBsRD2iQKhe
gNmCssPrq1bhUifrUSi7k65cb+QgXafCYHW7RZa8bDPvhKNG/i8zB0J9L9zWtqNi
KDRkbOJ1KVeoOiZXDDXoxNiBnfc7lIodG+bFsB3FgrxkuFY0DTch4rZnAO0BTYcv
fNOZUrTTQUUD/2+slum5PmBF1jniYSAnntMsaiAsCbcdHs8mBGWJubP7TcAf0jWf
PIPola3lGTrYJOCwhG/ic053FkOjJYWTK0MMBB1nQIaEIId9cRV8r35cgWgRJtdf
BdALjHOn1DLbDyXt2ZtTtX+J7hsWIsk1WprzeYt0/nDTH1Cr/M0dUPHlE82spFiP
gcQpCvaTeOJaJ7t0aFWziCyjDa1XsdVnmjusMiz2OGIpA849/6x+N2FN/70N//GN
qq0TD4gqczVrzwC6CdAhfyMj3zhvVWQmvKtAEW1wGPRj5aDHxIAuCJ9w2r0QdXDx
8oeUz9Sld244BG+v7F28/11zMbm25baZejNhFnhcga+vkraWbmZBt3PZ1u/WpUk3
BR9HSUR7o9RK57Qw1ycbb7hO0ceOysggkcKfxDCnmz9wSYrqRXW/A/vKeF6HB+H0
Ss6bCkFJ3l+4rt5GIZdnKoUjWT4HBA078tH1uwzFwEQhInCrpFC47qjfkYxY6VZt
HvytXyD5SkOpAiLwYDxVmWTeCWVo7WUfToPfAEeczY3ENhct4p66Dzw/BbYU/B8D
aYYSL7WsLLf0VpmAifpuoNOsbgO476ApYBdGV9ST7GfD6PtWZJB+GaTzLCB0u514
Cc83/hxdpCyJ9v67qyi2vpM+D2nYn8Rp0iMi6dNcKIcpQkav11FJhC6cIMcI6Uqo
KRdBsE+yFi//d2eIDc44VVXoS1BaLOSylmKmUUdMHMwYfO2VhcyImoxa8ZkiN5R7
wR/KMv+ukrPnD2p8Icg8dQXHpgJ7af0kPh0lIAVmIfF9uMMFhKgWmHBmNqtULNnz
QF0wWAQFJ78OWZheaVTiMcG/7kPAAPUaz2FPMCe0y+HUgEY1TDwexLSR8DZxfU3x
Ce64aXUQ4BhplYmgGMaPkRWxSAL3Z+KH1NfGJFEbF1neK77dA/v0wME58Bs4h0lF
+h6M3qSduFQRETiQtgr0O9UeMuVwUkiS7grpVjvaJXg5xA30Ewp3h/f2Sx7ERvr+
0CcYdiPS2ZbD4aamcDReIl6pyMwUSuqwC1PzEAIi1nWxB73OPfgxEo8qbyUhaWhS
edOJxE3n5KXDs3aNVIwdV6StEH0MkQlhlrRWbVyh2ALHnpufZ4P75EL6bug+1Upo
HN8AphaFsgg0D34DscxnrG13oeN9TXhkU6uCxToLzk6vpxv8y/FK+Foqm2BJc1n6
qPlZdOYXXjONZYtqP8da2gd/oJuWYnNah+0Y81cFkACePIusCe6pC2NQfsFvkx6b
cnxytmL32tI1LkrGm0U3klBGR4QaDjGwa+L7CUhfX2P6KeyAywsYWi94LJgY37Z8
Zciba9nCUo/PDVFYZ8+0J6TnLPFgfRvC+1eXvlqvmClEl+iLAF+i87/zn4FjryOU
ZFt1VTBEp0LZoKWdM0vWDesZS+L2nGnZKNxaH/IrkPSr4kKClGIiSwgyeSGX7W6L
GyFRj7E8hpuVb0hIyzW0OwuyPoWKsXJWClSgD1CJpX0QcusLCfh12inysC/xIgNK
VPWrLVYDL+dWPfsQKTZtDyLvpVpZnsL2/Bpor5im1FE8o57sruE16rpDay4heZII
cZdjgx27Br1EErvsqmHZ2WzPFwD6DhZoDtTBiDn9Phr7JIlASAQ3hXv5sWJb5H0C
pbNYgQeeClXwi0YSy87rRC7Ii0aWBDYAyVkrDLoEq/lt3Z0sNYB0luyXd5Zs6XC+
/IhP0s0fEr9PNLxHwX8u+Z8McP6/u1v+bxgKW5P5bjKSGiGpN2kcojODIl0/NEil
KkZOn6q0Hlem0PKgw1DcGo7ZB/GiNcN2/bkE4r+GEIQik3EAxPuFqjt5ycW08Cty
XGLWVMCL3xC0ErEcI5Qe/NQHRTaIkbRPCTn1IIvdkohsotpcX3xwouN7WawzFsMe
TDJuqJPbcpyeQhRBTbG27ylfGmI722UKzFUhV2Q2yFsobEbtLQTOq+e407tkl9HS
3XRaXYhCSs6E9HsRYlfjWLoH940T69WtAC0m/zbOgHChdDDUyTMC5jjoSWWhmAnY
LsW+AZO7bOLNiUyeHhrINpRd518BlPrA56a/K1VuGHCEXH+GuJuOSTzMjTiP078S
HKzFSI3zQ5q16gsZLjYtqloBaIK7oNKKju/J09yxr+/AiAV6q2IzgbB7JlLWu3E0
crZdLwGu9gMBewWpTMczjsajXBRIZ78JJjvrKlwrxIquGABiwP0K/+V9Qyvnvi11
NODI5Wh9HWtS7o6wRwJfW0d7983lDHpTb+JR+L9qn2dHUW6R1YupXNp8PBBv9Ryc
/GwLZ9IHNVyCXzzH6AlZEBszQs9VWeR1SwStuRQlt5E=
`protect END_PROTECTED
