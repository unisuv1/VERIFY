`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M6a2He9ADQ6+hWlG5uQ9wLLTf1T0Fz7yYYOBHGs8r6w94+QGr0pITCR7SHXV49l7
616NGWSrF3WeXg+7MHbTqVT/lpw7iQ/Lw2HLCLYn8Dw0ScuXnydoYZs0foHZ9+Xl
JLR5NC/87svnHHRAhQRA39PIVnEi4hjmwfiQb3nEb8s/cLGL5c16tpNzMB9ka2l2
17tMm9fpDHpIAg1YHVryzzAwvDgCxafdD4oo9E9XJyhLS6y5sFyip7+e8psKejxw
9UVZBKekn0Jx0mKTlE+0CAJ6ox1BsvzUQpV9m/Vi/+SnleA6Qev2D7qJbubRxgMb
yaaO0N1Tu+v+7B9cGbAbmD9jfEurnGclg6P/5j8rk8YTTtBmCdSamtjp1HAd/coR
sprqdnHuIyMbjevJEOZLbYdNRbiNyhRsr/RGWsWrk0hMI9ws3YjhP6NVx/ndGBZy
vdW4OhGcMIu1H36VpA8wwAJuofBUE6PQV6vuVyIXUu5vGwiTZfK9qWshsH7FHpai
OuwF+RJYAWTgVxC1hBea0S2raBAnzd0bfEKSd3uqzzv/wb/JPCCTmk5LI0eujjv/
Du24AQyy8BjWRZMGZQm1D1ioBHPAXP/axmbbb+7Nc97a6ImXRia9JTbTlUAdV+7y
ypgj0m/jT75uG9lbww5xFJMRKBA1NilPHAvpaqouWyqZANmVP8IMIKlSufZtLkjO
PynU/a7mbQSrIQ6V3rLIR9iAw/R5832CvEWFCuog9FX31szK+hx+YQQmijQF1NmX
3G3dq2fw9VcNH1sBVLw30k6aQ6zkfXFAShqgpaTLTjzOV7afLjMpxIY4SzvEz5pR
MNA+MlmHiUv2ENJML2wbcoY5s1YrkVNl73MX7X7m8SLDqfKMRpDBd8Ndob4ZLCp3
BGmwPwaSofHWYG4MfWivwvL3BAgU2QhbUM8nEqrpGdW1hlrosMm75DG+9uyX1UIr
/2kdcr/vLLukXD8uz4Mhdhf2ntZhUGEIG8xv1dkz+qTwthA/8BsKcysCDUjVM/Kr
z48nBRvIuhsFlBHiriLl0SkWeG9jzK4jpTxjR1LX4FQxk0HqBePQCcwTcwU0mdtp
dOJsWTyPJMZSOYDqE0XamZqC4bnDV0s7dQwSiWR9sknpKdcqT8spiXE5JkfhobtK
bykxnlqCSptCiYn5hbjk+SnlDwn5ik+c8UdcIQuoSzSf0vZN3DvbGHQM98wQVELc
wk3n539NxDtIG7NpieWz7pAu5qjfckDpM0jgaH1mhSTCzKw4cTIvoy73202zTHHc
fzwzbkBFFo4uBx4qb5hkKE5Y/GPgd0YtQJtPJHi48fFavuGBw/DzMexHuvX9kq7k
80QSf6OvTX7/arz0z2r/i82YRx3khJknbxCmJh2TLlUgIUG91cH/kMs7sw1RRpVD
Z6iFYvpJlfiBAKy98f7k5YYJjL7JoGRiEP6eyGdQ2LErC5brSOps4DKYiBwWqCEr
WYHnLqFbatbdi+O8xHNiim5B7EfYNtpRbwa2hvR6SU2Q/1qpCwIMnnlr+C7Ica1y
nAuPL2Jno/WmjO1S/TzJbavGEjSm2AJZopZ+LsD+qUwxnib9dIUb6Jns4KkNTWJU
sW74Zhol9yuoJruW2zLgrSVVZIh9H4wKgEPs09UFVNxmAyRnD/m1KbHxyx22h3eC
2LC9sY6lQL7FdwbmLXGJS4RBmkw0lhur0wvIuNrE6xRvH0NVkEvqPnRdnmyntuGi
QaVrYowUH8sWwCYfpdy8yFY8h8DmoNZRmYSq/TX4gt26GiJ6Z384cWEsavZOuejc
TUsfB7WhOmTUAOFBelyS4wOEmHQiD9zw/7h3Rs86RQAaXpE6lQYQ1entT33SYNpN
8v/kLJM+5i/71oBmfILG63+Ns5sSrS7e6jtPKk1cNTOnJvKKuAttoPUN1KeNI2oH
I3tZvuKYRWbhJZZBXzu45FWbijikxG/+oiU2cShy9T+sdp80n6+2r39Oo4cUfV4z
AYXh8EVcjcfVZrbLdHIDFipc2xJUtnztiRU+XV4tAIlA3mYHv0iBLc3WZ/I2GxLp
0xDLRAAeyBM88Z7W/kazNuN8cIyi+mRoGO5uSmhVNUaLd/x9Bswa0ebZ2IabEErf
4N6hrjpgxohEXs+ihGYr5Q==
`protect END_PROTECTED
