`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
cL2MnNIiGzoWlT3dPpBm+OkscQTitKA0uci9blIRbN39h+wxzH9eiptMfDpIkwYN
zlJ5qcRNB3LDbAnwDC5TKv4L0W7gncj3nTp2UI011QfdN8Oa3n6kh0WkKEYQr7Pa
yJdjHZVWQF9RThlWL8isY8tRC5IR885hSVDUTpajHAyq7egOF7R1ld6cN1Mcxx++
SiDFhaXoYxyopgx0RrOrHPOHVbwRuwPfO5dbSwoNWdjo4ETd5eY3bkO7ypWOpC3L
/0SK2O6pEsmwAjuvGM2cUoOP6ojRMuX6o1SqRAUqAoc7mQOIlT//XcbtAlnAaFy2
6gAbpKyBWF/NSLoEXybNzdru3fE8os0oZMAiX5VlKGNIa/tdjCzx6E/CtoVXUS7r
9yAhQVEsTSmq8zGQXetF4Ll5ui/vw5dOqzJ7A525xIhD9Fy73pBdfGZ5XsCyyYzx
v1E8lgHY8J4c8pqeBnwIa0Fr94OPqZfqioLFfAY425BmVDOrrjQGZUdDyLCbjsBX
iX2s+u94xUSGsrq+UsB6PvRK2ec6/4+IIJgeR4KMtt/pBvaX3apZXUyX6cGTb1N1
4gVjxPkdXnH56EcX9+Z5rtPJtVNyB4F6icy/0rjAgWWgP+ebqD/NqjostHT/8lJt
mKi6SC4nhorst/gozOo8rR6fovUJuBMfK0F7eyUzfsIeHnub5B9g22bdZDhp+s15
gQ68arZcqp5OVVR1qBgaJL3+Zj85cYdtzUPsS2apbeUH0TImYnZTG3MKwGDSr2ko
1EaY7cxKrHHcF0Tl0zA+6DK35UbGX8GSVeG1Fm6kp63UOTgFgo06FdWhFCr3DAYp
JTOKJDddrhy6Qej3lLf2UB65wYDz/M8lS3ewfvZGOqrhGPRH2/N/CjclBQWsn2X/
2qhmUq9EEnjJqgXBLi/5pSMo4OaNL7RTHX4RnSzOMkNC0OLqZhNeX2odkkVe7IAy
swK2JWkYsT/oyTDhY/7aF68+RH0UYSKGSZGEAxGArMKWAyBlwLzgmhIK08SOzvP7
LWLO33l6U8BCPJG+S0uGZExnPkCIXtmhK0Ext/38daN4OQ7GiwuctXEXU+YI2adK
qcwjFjt68shaUGyyQOBFXIP3kveyNLkoM0g3syQlLnixizhyA/w92/rci8vRmGEB
b658EBz9hN8oBGhKN94IBhBgmAlLd8/esA8vYPFAd23zYoM/aGg2VKkVbtnf7tBJ
ascgFL/5/nRcm2uyXIrqQ5IguNYFPuVT0bOJ28yZ6pBspOSNNl/451oRBGtJb9jq
ff7kt3eIq4AQLRg7UKZARPYUWfqHHEjZwdtCsq8NciU4uFe46k9oTM9J15T5rUjb
iMHxG4CN/+iO99dJ+7jF0CGFbz32Nsm2w0f2a7v7xs25n0ZPAXva+IT+2lVrOU5e
QEwUKLixIkN/gGp5p83ZIRJsMUZlNy1UPr+vyoEymGvFStwV1TtGWKTG7SV60qBh
SdDkvoI7/NGlGjyLFMMOpQBtBt1Qd8mOPVDzXppeKNChDSOoe1OtcblHrmyZmY5D
Wx3p/6mR3zL72Ew4QgAoL3Q1LxYotqYBV29L6UZLT0GICj1B+CDd0T7UMBfrbEcR
AimebFOluNfQpi27mQXY+mEVs4bhZFx3iT9NS+tJ9MJkABPMJbmjgkEQDGTNDc33
R5m50n5Yw9VkIHIUH7x2OeQNawHAIB1Lwh8YYFIeLw3UOnnirvUaAeviYc0MY8ap
Y6nLRXEB6VXCaxKX3Iu0icMkObHTyygEbvHMYZZFKFNUW2I4x4Fif8x9bovZTaPc
ngUJFmExq7ndcsmhD+IUgruU/UY6nYn2JI9Mift9e5lsA93XNncNsPs47THtXpD1
zR9ZUgivyCsF8/qLJuaq66Um3FkPC+yVCWrgXGsx7625nqDKl40dF6LBa5ZcP8x7
gZFutSqEHfpSTnsCfNDHDGbLrVcPTxAuUqFRWWlaIB4e4ytFdhP3+lt1c5VR3PnG
ET9n2kTyBP/IKghYQc3CiSplramyQfB0gEqopgNnTEVdFP6F1WBAMhyHiz9Ey8rm
4DL0zZoCw5bAB+xrZlt5RiwXVPbigvH5bTKgw67uwVTU8XySRLPC3LZQ3rHYLu0p
N567Qi52W+8YFWqy7tpYuVkvw/A//fWk8dWlis1xArHJdIiG8vvrBUXAtY+4chzM
syFzikHACt0tcul++62SqXKh6T3jokZ8O7WGW/2Hu+DcDBNYr5IbG2dFlRocYvKQ
K2+ClavELCFdtyqsw657k5Qc48FxSw7Ti69ayUyOOeV2Pivzc3oAdBVPZuVsRYQT
rLiR+uz6AJc4/Euni07crWCOrN4+kL3vskkAESv+D1GRVOYV1HmuXt3OsJtvtAy1
ZT9BXfF+tTFOYvLGlcz0b1LigBOIv3AbEfY54j/dg9fPcma8l+Xr0MWa3ieP5SJI
aZhQPYUfScIbGv8HI7LevDBh3WlzkUF0THfHCq335scS4zQ7FjT+Sscv4lVBdlIR
5tOcZn3uwJDnNASZRrfUTBr636ZniptKazoGOdMEyaKtGDnorioG+nqsefS/Jed/
Jyrm20Nbi3a/akFetcp+Oox0RHw1ELw0Ohc+MxG8RLAUaDAPBn6V95d8OBX5YbZM
MSVy3A1HoTk9KViR5G400Rw2y8K0nLBdVmGARcg+5BFV0EtBIZgPwxO/+rdaiEeJ
cLtM9UDptz7/j3LXHyJud3o7BT+RWHvQW/FAXdglslEHPC6gLWFcg0I25P7UbPHv
XVWZToO+U6B4WNCspqGAejLi7LQuu6PikPgGnRhqe9GJcM4KJZ9INL5Xbzm2Xx5d
oHcINdYrF0yUcl3KK7ORevvTH+f3rSiMELvO7mAkEVXvddMyvrSwsjmg0JEqzr0X
PtfriWDq/vHSX3ngWZs+VUrEiKfQFzbTPq60X+pkytuz1F0EqZooWlBkY/XWDvnh
vHFlsBf8wWKgpshvLEoDrf6kZcRscaRxGq9gxggOCsoH0lLItKclqbpvVLUjBQow
kwDIn1GHc48HQ6fzBNoDUEFpF8hYvA3Fl5J2WGOvCj4xu+7tBJHtR3/w7en+U5bP
bgY6X1TWNyQX4ffiP1R15frTGkFuP28AkL1GIIH8VSisXGzCpq2YongQzTU+bl1Y
A8SwCYiniyeolZKkF1qxxNIxeazK+ehsgIMSCcpVCqv6xUl3I7C9GWsjIbDg4Pv4
7OBnBUseJlT5cE2nlUy7lI9e3AwtJxRL0T1Di6HArvtVmutvmUHA7wtUlRiFdbtP
HJDfc3jS5s7QBARrbmzgNj/jEIJJltgnyoufEyf53lqwu2z9rLDHsDjI5w9qIVP0
5Ej5YoFpaz7REIocM9Iqa1t+JN3QzrQr/qchspVYphTscjVSOluf9OepZqRxXtEg
OheGKXpfu+amfTaMJwoHu60RnP2jIcA4ld9uPCHxMEOE93cytg22TAYKWx9aNTFA
T/rf5Vdt+09qhymAtoftlwJMcI8BUmPbgngmF/7x4V4bJXhKuOjBOJmAqEhAy5Ss
794SbWWfO4agmt+OEdADTKH18Rzf58Z1NW+h6P6f9zWhTj+QYwuoHYE34wchSxwq
+JZ1YjIXi6j22omCq2dKkBYeucHlzGUo8xdd/h3+4l37UyzIzMarrprd7nUypqYp
4RSk9wF5hWVdgluMf6p7RGqysrhCASKNczQ2Bng+dRmw251sTXA1tYhg2WwOn3GF
4DrKba17G78AYTWvUhNpcRK/aE/b4q+QJDOAm/OX6ouEHQduWaTM6CtV0dM1zzB+
1uzoO1Hu+ik2BtHiNucpPNSNtLxBb8YQwTTrogttW8toJ7q/+/26vri2QLv9nype
AoWsoIYVs1FVa/N7Yng6koW280hCmM7V3nk+TmsLoZ3Jl8ak8ldWDBFmG9BIkgGZ
U9sBalLvTLXGlmJeJphrtp7Ll2GYz53D7Gi3JyRJQIQc5crwbIg5wadCYfe0IXj/
ur1hIAECYV3tL6VUkk7/jGZABE8t8VPhbrVFPvPCOgwyo9uqRp6FVDkhRdd3+/71
a9hQrkvHvHW3k2StiuIzJKmvT43jrN5JVg8K0GWQe/bUNPe/AmEIvgP2SPPRstlA
6YIj7Xln5SBKTkAhV9x+fbIaWCrzaUaPWDfmlwGXFnybB75Q3N3wyQ6uKt1bp5GL
PARIIn7mGhyXZivBMOM4rfMoe/gKM5FUHTfm4tZD0ARG8UnONpSqIvCu+CPykzuY
qMgdw/Q4IQbraj2ieItAykjQG1Z5agSEb9bi4rZ1iykBTaA7PTaSeEyTpAbv2EZL
UGZRK16TGOMpeerUq5U1rL7mEDBkVvF5TbTmcRcHXVC6Nqry2FmKnhBBJ2vsXuFL
I4op71fRCyjBQU3kcdYEV8iudCAtUjbQm2pgWFhUtta5T1a8QK6MlGGHv+TF0Nem
gmMNf6939bqhlXKW3xdp9o33PSdmcsch5xZeDbaIjP4jNqPjkME0aeUa/1ZN063k
I5IPeJRX0ODvFE2EFJfTr0Rbogfgl/28J8fpGYb/pNi/UCJpDFKVrT60Q5sSbgLp
fJj2QP3llRTAL4reYbVFWBMNODzNEpus1vQ/rxMS3wTcjM8UYTZyNBz9Uiz/NqHf
JvCpP9xUJCk13RRaUJDNEtLZ3AUPXZGoEjP+TkGNyEMr0I4upWXeSVR3FFiBy7XV
r5SzTXfeBF0LhmPobWNZCEPk34usPmapbpvDwuuhluBP3bssaL3ekPL2h2Ci6q6w
igiYoCw+vfq9x6NEEilWzDS6wkajIvRJk/Ck1ppdJ68ntnUZ/NSku+ePz6gE8Ls6
/gWoq9vIo2/mjbmmXknxXAw7K7DZU64kluYnmbZeZn9paux68oCKrM0Y2ubwb4vD
jGvVlXYx6qkGuaM7cdHcCmf3TQfO5wMRK98eIOtz/OOj9hSxWZfLg4R30brysDKv
MIjV4wtS1/U2EiSjAKG/knEWbqU2/fEZP6QviLVGZKlcmclpJHuwTRNwPiPkPwAR
5PoC1BbqYAhkNxenDpcDkXcJyFVXRA4HYBFYIJekvOZJWoB9bNJuhIPWmdwCmq+N
AWxXMcE7MUtq8Vpvtm8WZUblRdxuL6G+2/mMuVqUlJnuKjM6zZAdTv9EIipCpLzY
8yXkvl/wdBcKCk5QWmdViP4ItDkJlfNU9ul+xu7NVTR8BZ4EgD+gwITNhimthxXk
Y++nMesnkDUbQev11Eg1ksdVxNYMXIF+cn2YULyHW8EChLkP+ZaVrTft88TrMwzH
xdL7Qcxf2LeT28/VEqwlepQXDR4q5Sr90BHSveUSkJpmR5DjzCCvTWGAY6uLf/rW
UuZ56fq9r2kcBwYw0g/TuyVmDdhK+G8b7L42eKTceXwkB2eBsMuxlS6hmWExTvP7
PVPnYwQWRB22u9G4ZgZi0zjBIVjXc1Psh1AlNQ1dzNCjcpI+FeWSGOPiwTQSdgtc
3u1znBhRtNjwGfWR2oRawyioqBu+sG89eiO50nZQPHe+kL2ajJ7f0oi1tPNEzPde
wYpXX7I7eiawjON0XCLVyDeiXFZD2MprVgK10rRLxdqLlKYxZrlyEG8Vu8dRa0Pb
eqbtIvKNtbSABvjH6Gj4/RutE9LedQf/Jy++jrGnjHhuS347GVcdhrCXrBjTn9i0
/q2gmfZB88IVniitjwwKOAom8d9NFJwfDFsQnd9wUUt36zvDekfcuIQUPZ1iXrKD
c/p6vT1TccIAH6Tnwvs4JpDzQvGHdwnvTp7kdgsJiVECjDVqZXze1MieSsY1F9F/
Vh2EnNM3o4B0wQgl8KwPvhMt2vru0bxwscxXe6Ymo9RVoTiT7+OSoIgwPIN2uPGs
+cQn5OzQDW4/fTzbjAs7lSLNoyD7XJ5zciIRgpBKD9T0UmxmzWI/lP22fzCtFRr6
RLvw/gvukn5y8DTMkgSIotS2uRp0SuMSw4xLgfog8C6tJ18QRTVveg/QerPOCJRG
jk/afXXNRifE1CN5E3gCF6oIN0zUuaxSxET0lYR5SrE4OP5XdJx1lFbQEJws2CaZ
1LVpNNknT+5l+cOl4/9z3sPyQ2OFCxUCYjBSH+/ggb+NQUZ5KNIkc2bfJL+WlyFm
8tZaLuPGxUr8Jrg1VltwJnaZkpwp4m8wPECP4+ouj03AtEO77TZUQjdpTP9U9uDN
+icyj0bjKcfUvc5GAmDHze4tAUjztwmbzlVlUTKAMSiN/Wb/8dKkzVotU0jYtgvo
qKqqWdhf/6qIWx0f7qotkwELx7XV50/eGiTOh07+MK1xrj9iqD5YxcOUxzDknuPC
sLTQy+Nml/ptkYIiS6tnAp7lSqW5C3CGHcRVCFn1f3eZ1JdakHDz8vX20vOtqjhA
HZSJ4daSVyETT1sxtMChxzVc7eiWV/oZFF7Efzik26Js1UpuX+SvaKJD8cKnUgVF
5oRAkUhjhRH1uglwr+qvsm610WytT2NlAoJ5g4yamSE8vBT5PYyyWsz1Ab5PRvye
KUzAp+JH2SxcPbiu2IRaDXEW+3LeO68DSHb4OeZ4DELyWt1m6VzdAC3K56o7xcQp
bunfu3CTzhglo0Gd6Q8vD1X4KbIsCCvDAwDLOdUqc0oxzDMW1XlJdWxGLq74Etdd
7GNpRl0c3nlNc3Lpyj1tZcpCtuny/8tiiK1NU7fA33FpeZr0+2XRW3o/IAOFW/B7
WlGE54sd4CB5cR/tI7R6OoRdLivek486TnWKvioZFubHR1nbrgp840JB0J5EZvz+
g8AlWSJNLjU75NqB4ZN/klsBJmlUhSuy6IFDoOhIzwy0Y2mK5aenJYDBi0+123LF
iKyj+d1wvWCk9hlU3Ab3upbazuBMXM3bDJtQr8Tx5t5OWOvYWbO+DK5Af4wV1NNN
F86vVFNE/7KqupWBGgz5XLZ7Afs6J30bq0AEVHegdEnjPzCDAe9GxdrPIsHhknyV
rY4Wlyn8bigPMpqiuWH1SOooCVml0a80a0JH1tSBvcGSfm0lL+oLrkhnnU5pghGU
rrwpNLkKIt4TO4gNykQWb70X/tNdzzPsfVOrOCRXAxw7g3Kt9JkSWt4O0NBI7CBj
vB/YkXDS2/qL2a0wP/k0X6zjZ2dbSe5cYVNsuNUk1iS0a+5I6eqH6/SMsOpSymyM
wPEL9lhOYYs2PBAMeb/63FZ9S1FeXvFbSqUb9jQL4CdVXCIwuyocq+2FcD+E49GI
kgvmzugKdEE+jVuHkgOpWi81Wyvn3noJ7Cdvk43wWR5iZZWM+uvLyqoFiVTIRyh7
X34cqgBQmz9HL5hzR8sQ9MdVyoiF8/p7T/5aixHRpDyF6cqVqYHf6+2FhXGrtX8P
NHRM/NzYm1R5tfshidAbkn83uCAh/YdZtAK/9MDVKZZO6Jk4cHDp+2RieaAcqtxW
61W41WXXM9YbXptl7BEAvjyXYDX1BZKe1YoeN7bHTCT6UUyhvHrCbFZ1yZNLTmVS
n+ksjzFyOGi0dNb0AshTS80WAhCQ0RZbGjoCRNACBw/pwBv0IHZfVC+FiaowBXsP
jOHWSEH6yy33Unmu2i9XWfwDiAcsDlGFvuZeCfYjbuJlSZQzPY8aszQxoxu37TpV
goqu8sYYSemnQWDDCNmizxKyEttOq1gL99DEA+T4cuqjy2iE6VHLvEUQ1/UrzRIo
QrgqYV7I+Wey8peDLuPWywwqHrsn6HRmyj9bCHuAGXPKQmnQqNvXVEh7NzIGg2Tt
zBkQllmo3fHdPdC5zCms4IVfiRskQFOy8/Y49wdnElm22EQ0CCp1ruGcMb0Ufggu
zmXyeT3ko9xE2WDnnUAsogyNpsxFDW400E2zpxH1DGFiepgyDtKESAB+ma1ZguZ/
QKg+M71dbGN/XlGf1gPj7421AdOBhP9kOzmMW03wph2WrvbHxd08sSEZbGOohAs2
cT8N4HStTsdwhlCU9lXILtP235s8dYZkj9X8P1vBZXlEwZX15BezL1G6UAtoF+yy
Bp9ZLJuRnvMygYcOIBkE8RJto5QHeMALWNmY614/AF2b2QY1DraSNnotZw+rXNcM
53plpOEtyhrVHED3+JZkjc3x6HZkjzqgbPqGDS38HbtJPHv96Wt759ZpluGIBOl8
AEXYBReWDYI9+hVm2LOjvDE2LmM+F3x8oZZQVInh9uGVgMHTPRd8NeqVSAYk3feC
KyjZ+Ok5NmvGaGzWgEkG8HOurZ97r+pKAvbYqlLPeYv3ZtCteMOQb1K/iZRYb9rO
rCCJW2SFjVAb1JQW4vx8OUyLbaZPsnrtb83oG4VAPgQhhiBPFOjRnIrH2B9EtLsn
Tvz+Wl3l4OEmxx0RPiWZb9tepVNKOklA1N4Yxf1ggejYM3u4Bo8QJZpkZFaJ1AAw
/JQBUOpZD3hHWFxq1jfyYGaW4GnPS2/kuSa2XEdaDRX1n1RRNbnE7yXwGgAKORB6
kB+i/iEstYqnZN3DaRtXHw4abSrpwjWPX4f5lzFg+Rwsp7+ynHQuAb9ntB+Ynt+u
6Zf98R3A9iMYLHPg6TcVoaawObd9uUSfPbNJyNgJYCRLmB+shO/eqd0yEposgNjb
9muoJaKAtjIbVrlGaEuEaTMAe0ys3SkL9a50sBycoxKPE+RMXhj6Ge0SCvTrKin5
gd/SHLJbqf08a5vXLDmhKowbjDXNlyLHGpK68QDM1r9xNI4/4m+6tx1wDs6Ug9WF
+aTvhKZcus3Lcp6JJhA7K5Sy4Z7A5z4NkWu/8qx0QJMTBPTZDbSbikFxGyN0VACM
3RXBOiIqQmuyYgyIRq4LO6I7qGnk7wTeuKrnIsCxgPWjSZNAUsVf5vs40AQAOnxD
eFCleXRKWhaVgFLfwoE4Et1FBtC/65Ld80kH7kLhNnkw7/TTWcmzOehXXNvZRCln
nq4ecC9pLdurgfc/3b9lyMhgEX/FCm1DH+Jw4drT82aAtr0x8tb4MTJ8fptOsfXX
IXWc5weCnEs/Odh5Qmzd1sUJFJfh9+ZEpijJ1cLKbANRjKbKNap6+U0Ty+xSqowI
Ggrjp2LH620tPB5u7LW16RHYGowAxPo5xb8IMCFe+E5d/A0m9SXGeIS1GVJ6HA/9
nN8i0qwwmD73qudaY84N/i6gXOJXLQs1dRzS0ZrpWqQDP35LGwrf8a5IkpWBmidT
svCqdnpUjloecsHp/aWanS05g1aXxsMZuOcDOhp92J3OXGRTYqSeH+6CQtBxRDaY
I2z/Ced0GmVhCgKy6T5LuQ6JpqAfIQ79+tZocmcAfUkIVhf1vR5pXAAWx0gh3qdJ
0LjNz+1ltLGgsKsVDJMnsDn53PdFnlc83MTIBlZma5c9KB53GShNDiwbN6neBL/S
BbzeiamVC+crJlHbi+f/kPuWpcr7/5nwyXvf0B508zvfAV6tOz6TAjO5ZstLAYUW
piw8LG20cuQu8ZUdRy8JjxGlJCx3nhF0xvVs6Q/1fSNGRg4vr0mcVAfe+zz6dBvh
g30Yz/KRWvK2OdSlMwgSsDi/rgCBbb06EIQvKjoXcnetzkhILixlecP6TloJBfqr
ErmX0y3uHdHsk+ju4+lgJzmHbk8AKA0CsqwWyikbAdAq+OD7drEQ11aPsLXb9qss
/gEefE85eubnaA0p/lEhx6miiXKo9sDvHMNg93hGbcfTgZb0WDLnTZPpNyeCL4D9
zhongQAmKuSmydPYcv9cqmgIDREYRA31KZa33z7bmJhc+SfEIv4UL57H/ZaJPZjG
YzKEmw6MVGMN8wCPJEZYC2NOsE3UEM99maAEU3re5lZd1zAYTTYNnpqCp+PT7nU6
md45salA3f6bHPIB3Xm/J/JPuupmaam2eRIJntGM9Zh29YRHv6nU6hVEuJqruu93
iWQ1hzdAvH6oESdZlLsd+Sv967KJEolyOCiyXEHkAMNC8ZeKyulNKJNaz/C7zaHu
PBthYajTI4KXxBxwhuyqF+/TItdxm4n9daiMZChwGg63fqZO8ROk5VSVDCkPYwia
GzPgtsaQ/T8dz+QTpq4WS7YD9XFV5bNzIhTg8mWfkZFgmybc1fCQmQkkI/y2bcSn
C+jO0Idbh4+djssxLBWWO8YVYsNTgO0EHFqNieLXUB3o6XUxFdcYr+NBoOrh3Hc2
9Ds//SJfnlCu96LeaYdZDkXjd+pyHO3aMDcpGIny7kpwMGNvxEPTVh+zeC5xwuAN
QL+thMyLSAJ5GwydoKONVNUTWbnce/nPKz9RJ+GhF9M8T373KRdLWvuBjQXgnjBK
6BPYGrPvI1zlgoKCPlEVpiHtKBwX/qUGI+iGMe3n62fvExL1Kh2Ex9ai0WWbuRRC
bxQ0v8c7eD8AV7Ff8U6YVVTLCuBlxgqOqG8KVE2SgwZtSUc77naThYIGvnzn83dv
TPQ48JQPWAm3NFPrm3iCBJnPEjRDa27AF35Mt04PT6qn61i6AJ9us4xvlVYwo6AR
yY4sF6rfA+RxJA2lOxzqsGIMtcFiMLYOyHJCsOZZ6jqcMYQc3TjK7lAJaznmCy/O
Jwe93lqdut0nWJlE86cjYSsfbjNtoU9uzR8TUkj09WRHiez328BG0U99+Ro8WHtA
rMmGH3suc7oKLuoKptMVFWbdoLhNO+IHLK+jk8ipzHlAw1svvcPNZroeAIMuGAKA
OdlCKGAEfGMSuxhs190ELFowpzOmTCvYB2UtfHFxKL1ZdwDDIkveIGtjL0h8+cgD
m2Z//qLH8ujUdhoS+f3itliAEGOQ5s28Db1YxmimvCKffLb3sA8+8YMFvhFA3A9m
xtNaKmSbTXEQnaXJETpXCbiOVBzU56a8B6aRLNc9eVqo2Kkf2tetNywn4TiqQTd2
bXqbRlSzrjSsRfsFIMJB4kOl5/JfvE6zuG/RFTxz7KXJhUG964hdiJVc2DC5+qYo
xwehzM4l0A5+u84BcLj5XT8/2xJw6z4sZwmI45Uje1ieZpX10wAIZWRqm2ac7C5A
HdWyJbKIspmIvev6Jz0ESmEzcHUYiENow9M5v6tTcF2s3OangxRyh+Fd1gYitQ7u
lpYz9AQnR5PMVdaH8UyXvtIm2YQTT2FqBtHvOuh8n6S8N9D7QC2bacEe0pfPrgZu
o9LxhyoegY0olxjpyVZqYHoL0Fi6JgK3pTX+beXs5GeZ0YN+IanbxwbMf6+yy5kt
3EqPwSDI3RUnTKLHI93LqtaKJz/c17DzvurhAUyC3u2cKCYOh4YBqkqzZwD7FeCW
yXhut5lefP7KEFBEHmGIjoqWRkQIBeXOFmrMWN2PhAMNLxxfpcxLbfHoSnrWTZAN
UpY0+kvMwlpxw+PWuQZ/dGuUXhHu54wsDVwKmi/bfQSBSkoCktp5LDxxvfFKcH6+
IEixiNpYG1quDClQmBjIsBkZllhNUdcquru3sHXOoqfBkSEexBC7mqqtiXRHjT2o
w4W4jSl0tUkbJWv7xvpB2VAJk92NYbdr+SFsKTH7km+UVAgSGUW6b/vGhI3vY6iB
H8iIDejWHIIgQmp0pCthmx1fgzjvdIdjMJeL12f3w73LlrjaLLviaZI+wQ08qtv2
Utehehcc/iN2RMsSEVeNjV0DpU56QP19JCy9o92A3n8ayXEVX3+q5v96OBqO1rxY
whiHawFQxdhmr9SaLDleesUyxIZziCB+geBhXJ5nIL05q6xYo+TFAYRPgLwxojwe
Eu7YQ85/Fhe0NH1fXrcvTsngQz7JU0Wye+Zjc11Da25wWFEQxAlGmtCED/EvGorJ
Q7A9rG3xdsZrY+9gUsdU560So8V+wnEZTX2SORGz4bqyaNFfJwuetakz3ppGdt0o
gkI9DObW1WiIMTA+mngY1K2AtWVrKK1oa2CvUPzqx+0K4GZIHX9KprEdlBinKIQL
HQpKNh/xkBf/yIm0nHjTq1rCMoVhxVol92zICt30MALpNRn2GfUZBbaKQQq9SIuw
Ij02VFQY5aaXjSLTv4bAkhvIiOdgGIr4LYkysX38xkHcRukKJxJrNzLAoKn46v57
QtVK1lMhQyIYOdIhl07M7v0qyty1hgOieVhEAjHXuzjvJ1l9sH3j5i05gbwFpQWA
TKxFjOyVUUKLwdDpI66Tu5aiFsmMU+xZIcQf/o+rUdd9hOYGDXfkL9gULA+R4CJU
2PeGf+fh/XVK9prIto0XyYKbLNXQceQUOD4mQwa87eocxndM3JCCJKsbfYEcrP79
woNFL1OC94C8EsZs/MuMEGKzjAGP42YQQtYAQkgI2soncALL50wqF7mW4B9P7n/0
25L9xcv+h4l48mBb1Tw7w9lY6DtWMxOR7oAW/ZdDYmI1iqg5SkSwZ5FXWPMi/r8R
N0fJoKpL+t4mmeui295MwUwQHy7ztoAAauite880iJP85VKkkGKmeJzVAlYtJksR
behnRKsH0ScYAJo15BsMCG6NQtsibywgGCedaJ7f96MpJDojW8buiVMAGckx7It5
mFdvcSY2VdwOK2wsAPnhUuIC7+2GH4N+Ba5AXjXPXVexe06eOCq0W6/PqDr4eK4a
9qBe2KzbinR6ED4kJ2tOCHxSG4ojmvsMEFEO4nf8CDjAKt2otboN8zsTDZfLqDn4
mew+Afc2vbhrXHf5zfL8JUKp7cE8ytU8IU7uwTBcfmtZwy6h+0TwRpQpdFOec8+A
mYBSwvR+l/4ILIDrXUnu1CvLeXwXPQESlWW4rpipcmaRPOf9c9be/aexFIgM2niI
dIIJGCJ2qHkrErIBoLFVmXtxBGxBQX9D1lGUrHWH6gVFAcuB0wx0AUYulBp6axQR
25THxzekyqGFeX+u2+4X34DUNSDR98HWmgir682uDJSZCdg+lnujcB6sgg/ZqJB0
Pv7H8LVzK/Dr64XhlD8xfy8YO89+SVeXrHHF1GZJvnR50H6c4XmaK5aF6xRP1xcp
hgiVdxVtZmPVTXYDghPLFxELH8Pp2aVgpGnUtCi8zLIS0qAkgu5RQUYqKihR9acg
b5LX8+Ch3dj2aqX4me0+ADXaZeuw/kQ8QklSe5j6wUpVzxV879T2PxvA2zAKuNfi
LatdOttPxkPTVXmeJKjqSw7bdTiu/F3lPP3wg/h0DPRSdFS2xfddHlMTCjrbaMtN
v9bvANDpK6F79WEwtE2Z4xZFolPKb7dD+OPqXugnIalaWzTtU9LOmS/0OQrMPwR8
9pPg68GfR37jXypRMZQm67qZuKakYOgha2HTBmklT1FO9TSLM6+X9oyJpIyyqwj2
e2n/TmGem/hIrolU3jBQOVIzfk4VZDm+YgDAx+NZwaN0OkKXaRrdjlrrsyC7wdoE
aspQIWhaJV0gAyG8SyKmVyU2O8Otqp6NfWSArnJYHWymEKBCY456leR8R3ZCQIiq
VTddkeMWEcuZ4AUMZmW+AMO6oV/t8FPEmgMuDFTKpDQ/xj2tn+MUE7QrFmjT0h35
GGZwsaVWXdxQK9GqfTNXIA==
`protect END_PROTECTED
