`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y5TujXfV1W9vM7KuwpsJmOVIAAV5EuijpP62TdzcWXadxAI/lVN/9RWO+8GeZo5/
NFTmWOi+JzkVuiBFXc7GsTjkEYWHk4xVySmYEPhconxM8X2w1FyslwmR+JcODM0U
ag2wWj+sZVBZJXVLHqaZ+cXj6Vt5xWXB0qmA3yGwiOXTcqm9xpsk5wxKVuTOCOsl
EprDmGOK9o+TI9uMSYO9h9ItkAKHj7Jk8CJLNnLbgCFY4YsPUqq21fv0JG/phdkJ
3Jq0nx3ynCvPSgruJVpwvplWvoiD0ke4iUz2FzeUsiXYpAnL4Riju7SyqRpgamgb
VeGamOF4K4WfRqHdbMIDzjA/h+BVb9GZ6zw1XMpa5G8TvNmkmCxkNUsb3/IhV6Na
UgFHB5U25KMVkIC1SuRBWlhijUSaY0vQtNptY3HHjsB3iq1G42cvQS8qXZqWR10J
Qx1eHbOBs6NWZjKfpXPo4NcT4Z4MGI3HcUYo7WbbBPQXC0SG+6PE0Y+eKJcSwSWD
OxHmK9Q+/xENCYrpcxkibS8flQYh+WzwRJegM6EGYyid+ovT8kINouBnkNIeknGS
kS5FWX+Udh/9YtLmvphC8M737lOTITYmLx3QuXDmJGz8hWSkZc21VPuZhBAQ3L4v
9r4b77Up58dFtr4MAlGxbbK5f44sqjRGHbmCIbQZrd/XVX9EDvjICvm4ZDJ/BVzN
T3C22uuGYWp7tfQkQqZSWyMPCXwYbplImuGv1QkBO42hG19hjjkki2zzlHpTgZUE
uLCOgF5ZhL18K2lcXYpsAsM+My//QR4lstYaxw7zAVQ2mxF3R2xtO3+IJf7ET2mJ
6VMhiDSuc67EdjWY1DFfl+po76O1GukkEydHg+BUT5HldEiyuQ6hVl+6CpCY5/x7
BjIDwQ+323ERpvmO3ebbdE0OxSW0sF6bor8ktE2MD2YfIZckavrdXdrjYJy+h/hK
oyBvMuKMFNh1LpepaHM+KAlF3YNvuA3+KkpAnGJDF5e0XsjPV2yXAD7XIIwGlYQ6
+TbNey+OCk+ckmfwTfNXv5gh+XxEvg8YWA7sb1fBjOHs1lzsOcJyNPodHuOzxnqC
00rwwF0rmzc5XDa6PtEW78iv8K6AXolXaxVlKEStDaYNiM7dk2uSszGx77JHZc1x
GlSa1TjWM808NIbjOjDlp6tHMqWpUfVdQTJmVlNck+C1gfSuJt3rGT/sH5qPUuzO
pDuBVcAb225lOnPhftOEWMfXHnXDA+YimYBl9k1OxDngASGSnYPNVvTok5GMYIGU
ea4fpj3WWipJnP/nAKZiOiGJF90KwJdoJxLiII0rb6PIJ8v3WxS9wB1N1tiPu8Ko
p82QElMb7kmUMB/2AmUpeJE54NOcUVHbzwlKfeOcSxTZps0m02Ovs3Qk+VM/mr9y
IJXogbeMI7f3qbOQL/msCIJS26/qMNmVYe7Q7+T+JKTiYwv3GG0VIONUX1veBiDW
sDMPYAIkBh4pEaV60hODNvjFlNYtfswMWbBqTP05MrF7ctBKRc/X5ob41QMm8nEa
FqSY1UCW+wkFD9X8c2tsZtk4gqzclhWK+XnmXqJjfcRGBjDjNXZFUoaXReF+kBM8
s3SpCXZ4gjXL2dmMVFGjwccnA0xWXNgD9lzIObeQVhXqDUPe/mwzodkWYRc17olE
8tED8uMRilQ7MWFTV1qwN70lLgTF4KymwUeRObjehtNVtdlj+6odiZSVulJKIVPp
GBo85skdKUaQXsrUO78pXRAkSl/2WyTR/QuATvSfsLFPJKr9BjouwdrvSIzH3Nj6
8pZNMCuLcqkqvxbRD89ibzYjQo9dy/Doydn2FN7lGS8JTY5Eo5BnGKcyJolxHHZF
c6oK1Lo8dtUkm2vlZ3G06D+/DCeL7dd6I7PAL6zMW77lxiK0Zh6p6O870GnjAvIk
SAMMRfWy0IWsNC60WDXEbO4i63csLIaKTu4iB05pp4FdWs6/jltrgh3uuv72hktR
HAC0dzHfbY7o1ou7bAc9eOqZmH4uO+l1eio4D0oJZDjuIWSx0LsK043pQ+oQqogj
tI+FcdKfLsimQcxOphqdRuR3WanvkDZWUc7LeDfiC5j/ZwHlhCwAaH1Y8FNHrqWq
3X4/1UA87iOCZ/L9Wua8PjZ7iOaRizhG2BLPKoBdVkoNi16cIE2QZPZJA8hSyagp
QK6Oj64CI2o/Yz4lBb6NJF79BZQ/o7CxMtg8StroyKZm0IV39OKip5nfsCjROEeV
RLNK/qeNDR8llXBhMC8EdRFtYj6c9YWaBecvbM48NlXVOU/WZKbWdug8ww2w5Gwl
H9kiueb8wsIJUv0CfqllxN1Oq9/Sd1uiFPryg6OtSNcOmtBgiXO+CKPlysbw2iHP
jeoYw6i1weLZzpMIjLmKLgy5L4kxmzX6lKJqro/fvC47cvpfpqHJSsyNd6N+Ka/3
s2n9w20n+xAm9G6kdjiak+OfY5Xk7Y5mrWxl97okdCrEvYnVHZqJlETwuiHc1O/U
OzJs/C3pDVt9SND3JKi29JHXlSABnPxUiXQhU0r5DtRX7Lg0drh30cyLfddkv2bU
Qi9DcD5hH0cViP3zk8hqI1o0zTNvNMEOuGxof+yfxnxWkYVBkqWeUQReDr9hUriQ
+VgyoOIeWvTO/xzUMw14Cut2JhKu7yDOeNFNFIZqgb/6Xm9paO3KVhegqL3zNdtK
Y1D6AGfImy3UNu20Obs7RjgDI0xcvYsPsbdDXRUDdAfFRMwhkm24MBtoC3Vqjdsr
O/E4nf68PKXUYnfltqs9Na5/VEL8T5Su7DbbX6wCdFf58WWIpYSFJN/pqQzNl/cr
Be2sIodMkjQ78BPMAGjKGJUKvGLKwUHbQgU+dvs6KlgQOKTISHudsNhUr//y/YKE
o1q5sjYvQ5GZ1KaLAZ+ptQrgy+MIqLg5G9N3Ew6PxpMn+znQ/tcBUr0vDVNOyEGh
dG4tt/UP28H4m6zFOGwrjnCOwilLCkj6iZTIOlQ7hxn1Vw1S2fGipm9k5zLdo/5G
460yg5rHAwYE5ZFs3h7ZTnd93ts/43lHFzy91zt5vzMyaF+qnh5mfewq8T8fCChQ
sDx8UmNzpX4F0gaVPdCh93xXR8DMNclfQIypFgpajRSytcp8TbI0pnY9DfQMpMzP
Y/H5XN3rDTBdpmKhz7U1zWQwwaHjVmdoRDm/sRb9Q4Sudy7NDyfKzHg/EUnKohmO
6zz90L8ODHBScgyCA6O3cEFy+56axW/TE7vJ4hfudC6rLDnGoi89IxcD73og3Zrn
7A02ix49usFueh133S6CaqUd9KHtHEKnlMa95YxoucVqVV0h+jv7jOs7US2nDtpe
uXFrc6Lo/yMTZvTaRCzxhvc2OZE9iTxT2JNc1VxZTK2y7gLR4f95nsGciob8zQGA
+hpmfVP5KCCiUV8yzEkb1QjjUZHDLUTKzeqAtvK6aP3NGN3r2fqe7Vvguq5I0o7b
PXghmmC/7wDPayopr//2uCK/DuCM6IfHeg599LXYV7wwJhU6hMwbvxKOsUNxSWZU
It5b0yIyDr+mjfQCui0QFnPBv9XQL7WU1kRq2zck5g/0ELzuweRjx7G4UBQCIQT4
zN6uFxMorFGGrlfJLm9hb3j+kVz7X09LAPpcyHLwltz6ozv9J/xdKio00JwgXway
DJG2oyXy44PbpK5m2CMK/K5Mlg7Kcq7lWJmdTf0AQakM79Damd768CahxNH0v4uW
awFVYjqDq7KxsY8qHgHonEL32r1aQybw3n19soHk2IwUNyR0CtGtyY9phodiOG0R
Ie+Ta0UqbNy2WzNg7FKY0dvJQloIoTuBhTYRhgRurOKmpTjZ8C4G8GUPyvVrtHQp
+3gGUndQolznpenTqCE5yPg1lUh7y81a8tpAbOYhnW523LiWCqapwQDPqSfL96ku
l08wj8OqIKDukNVull2ZcCG0I8UaDaoY5NKEe7pmDIhcFNifxPFLSk8tkOBA3GGG
wOzqbsZnbLr6m9hbrRvaYtfX6yv+V2noQAJoXDHPN19BX6ZOlKBES01hB+Uz6LPI
meMQOg+HKbyGJIkjZjd2hcMGMiPuk3jdgoTRY2MVU657J6Bcc9enKhFOOdP/YQW9
0BZYPXC08tnQ7P9K2+nRy5Y33XMxz5VekuwR+en/9XHA43rl0btKrE8q8a/gWLg5
9pygQveJoiwqFLKIYEItyAxi8GGnkhzVlSJ15yPDR8wPLd0Qss6mcoltWtEVodIQ
w2akRMCuLurZfV2EuRTaTpjZLY8iyNb92Bqqg2eQjD4mf7qEf0uGpXv3WYMlgG9T
0c9ebbP9WweNkyUNok6401gMjMVzRJjqeEBLl3hCah6SN4+0RzKmUpT/ZCss9w9b
l0Oh8g6wtW7CZzZMfQ/n6p5Tk6k9WafAWwkNYlRufkvs//Ox8JKUI15EdB/aXfve
cfyDZKEu/gvHlhvFle6CqUtW37PQSmQXI8lxpDIr4rC1IqA18l04G+P7++AdrB9F
CzLknYbQjE0JPV5XmJfb2em3aMyuEfaXHcnakksULvkPieCrOFax5551Hhn7txfT
XtGz0Bx8cZ7TKLnThuLbOl3JANQ0Nst6aSslZSWSebXvKQ8a1upe1rLmyljZMJ7k
DD9q3ehCLMtTU+ujOb1zVh6KzHqethgZFpNYQoGO8NppNUKy96gLKiMq+s1/+sMg
bkJQiPipgE4rv5BTS/kgSkG/EbMs7kWELBQYUuxG/73p2DXx9zme5/BNE8kzzV4O
gQNY5gguYwRzSLWg7LUxCJG3Qc2y2azbNFqWDR4BRzZADW3pymR4hE6RBOTaqIrF
ImsJwncsj/QkilS9ZnWmBcVW2cy5z5BdJ3U6JuGLYiPxf4Q+A/OcNQrlqqQz6ZZv
Qm3erFke3kqGRzY3ajtbJmhzFGhkuFrJLtcO8kwbIJYen5WvMUqy8xZsy/TrPV3R
0ppg6QhTQNUzh2BdSsJQBcJFSVWaoc3G96qTNaGeap5kq23jL0gPFdHy1LcNpBnU
FpH5vIiFlilNGyLW/a46M4G7u3cx2ZDIb3aqVIUpuHaJdx5h0NFT/6cfAVHoJZH+
H+uEbtC5u5vNh13VQTHsX2/XQw3m0/ZgcA9NXQKEHTkQK1liK7M1ld3GD61AIOlC
wyaE+CCreCl6ZzckPNzZ/dcekgCG807IRp+JHEI7LKsSS3kWMdtOnjtBT1DZCi5z
y8TMUatGOwiKd0Ot5VE9/UVsqL1/RNCWr1a3FF4arCvLzU41JZ2B9WKQ57FFT3OV
L5EYqYsdDUEsVWPYdkajKZ+zanmmE0ZnIehajB6P7HEOp4TcWdAIS6qdWmk9fd0+
4Vl5DIKqmWlrzH+Ed/rag5q/Sou/th6OV336RP0bAOVcCiXusKHfZakt0FRpac6N
+kcKqhW7sGPgopPCoKUobSDKrwZIoEOAwKIn0T84PYfpGVx1vpxgeA3Uw8iQeZZ0
diOzekTUuHHCA7mgZkOYeXUWfmg+nLpN+qRull7Us23AjY4/fcbWWMjfc0elVd1j
+Rfze8ivZGo/DiZ/ZSX4aoEIpBmRgaGzc+rpNrSuEBANgL6MrlP/heqzMPj5Gaa5
HeNVvl9FDlCXAbwAQQ/G3gD8BQB6ZVUQAQNr5IfwV66RIRQ+xkE/U3ncxNoyArve
e7SusRUeqOgqtRFa3G22wTpKFSRJ43rPd78ghtbUVAO3xL7NQycfDjo/ulOkXXw+
6y1Z+h6H8KdV+hs43edLAOykicis0rlBoyMdjnwSUqt+7lAyhu1ulKiwwTlhbOR3
RIWlDQWtQFM9IaWBBe4dNQrFkB+kx+RtIlzR/IUsqVnrabs/xUJ1K8OVwpVUaZBj
eTX1Bkf3NdEkfxJh9g0Xrula9c/qf4S1TI6SMtjss5YBmnDgfvmusDjh8xH9HRt2
VwTIEMPhOTbT3kktu/4UM7TqWtP4sURv5AJlZnmPkCCqhjQ2k/rbPtVWXXoOam2Q
5NNQdXWMhaqD2tniedCI3wW7pJEgZrxzk4GKOIKdXqTnK7t/RdxehUTuQgo+6dPb
M2HXyaQJ7IxnDmqfQ2IC+Yudpy49cqoQFlRmSR3wgGKwRk6grKdQW5mm5uCry2aW
pC6hofTLA6rchjTuq8UgpT8YQrIjFR/vBydXNrQV26va7ONrjUSrZaa5vd0kw+wI
rvBM6KKhWUfggyEIyJYEO/2MTlsZSzLR2RDlzWdgSkQdvhpL/uGmf4oKU/jitnTk
ac8vV+WsdykSfWjSvbPX/IGsbDtHcsksSVAVOdPItWK9i/T0liRQ+J4BXPQ6q6pN
TSZKRujZC+d6oFpmHH7mc8Pa5HSQK0eIabMhD/GuiS84nCkxJ6NH78U5SwZ17g2P
HWzx9XC2pIpl3rwzFFTT/PZbLOcZcuF3ZYv5SqrlJgBensEGxY3iW8v9KbrwrMa+
X7TAAfdTJnEHY+wQ/+d6+jpXgPrfC5ab6bcQPti6MNoR4DjyvxeFKVCtXImt+D1t
PIV7fK3HsBuDURXiVPxnQ7vSVkNpMUajSgs4NFsWZ+xL5HjTSdbX1jjzPKBkJJzO
BwMCl0rCQIxeVfSJSQ+/LXKiM6KNDp71EnSlKim1LsWH7YLF20lnVBj5EmK8eKPZ
OS2eLWxhrmgWiWoMW2+qCnJv4w1aWEtcZD2ukO1XtvfdoBP0IsYhD1Qfcbt5nXqi
/Bjr1x9Xe81wBqIk2XoYx7gTEl8VQAdc84yBRqPDnxZWvzX6AJcCwwITzrMxVHUV
b5UlU1ze8apvwzFdRDXytYcTzQGJ4kVf/IjRQ35uM9K744hHjGolZdfn4N72rUWF
TGcg+gLWYbsS2+R1EpbUgS1WDNx0hFb9CS7mAFFLMQBPMzauLAElOHwGvW9SULLz
srx1XHN6n3qzrDd7wuLC/vyn1HzusmXuO7IW9XthhL5ibkAoQcpIaSPPRMnyASmf
rirXLPkYl5f1RwRB+RftOEq5SkK2Brb0Aja3KMt8bJWcVw5bVtgH8Bj1Mrz8VOt4
svcCOIWztoTLJ0ba4x/O4rX2cVwvACVcb6K/8xbHj0Nrdqd+LKOA+Z1d1ldxES1B
cCTxVYcQ9gyeVPjWZB2Y+es8PWAfYnvgLTb7oidNoZ03svdT92jfTnrd8DAOmJ3z
QSZC0zB+ZcrMv9u0WX9uNDIBn9GEZUYGSdIUN+o12ufzeyuSHyySwF01TjrDeedJ
B2DOV8j/OJe1jx6CqxwWJbOtTZnf6YQ5dSL8FdT4M7vaRvGfbwejIs0KkCezKSiS
jhwrprq3PO2TGVKttb5hPvq/SapGChD5p5iaA2hnxvRusPnIvPGri65gcsZNvSe0
PucUzkr0LZ5wkJAx7hfJYQ==
`protect END_PROTECTED
