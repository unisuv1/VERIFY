`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SHUR+o5bWnylThNbPV64yEnp814S6a5Zwu67cT75XEBJTwXu2s9bYMW+qERC6t/z
aJi2kbx21LDG0BE3jolSIeJyfGTFcQdukGRDbgcSXkGfZaQ00Q9hKFPhSHwp8dEr
5c0s8Kh6sI3sXZ9NrIwJGg2lQ3rZjJCp+80xfdV3BZTYB6f1x2iHRTGWTgzf/W2s
oCTyLnLferdl2jMDhJm5GIS8v3W5FYECpMtRsMQ5iwOXLqaOHG9P2P2x/jwcywye
s/nI1WFvEPAPItHA8inZXVlHdEIUmA1/Kl/Dr7UKUWniuJKS1WoBHqW+UpaG3Gu9
qfCGgqlDxeUoYU4vmn4yHSX06W1rhG7yQWBti4jY2QlW9rhQFAG3g0wG4IG9J+1Y
61A6x5U56RoAE4r1LaUpTLDNBwQ+0J8LYSSjiBPpjroSuQNJBBq1vEwbCNDAzp6z
wqJHHQPH9l/fOpCUKdlfTtgj6rsCwS5PHd6lfmpd2RCdC/JzVaM7J2KFTOOTY9nh
xlm9sTmad7v42ZcZc9HLTwiD7rMO0hoDBvmXk2fPb9q0xWnbcoWe9dY7yWDoyfe9
XRONrJ6XuWNQgsYLAMQ/YtnyXFxmT1GWMAySWD5sf2xSYv+A5X4llcth+CWL3/5s
sdQzJWYCz0YH2xj4T4x/amZQNQNK5Yn2an2hDiSQf9DjmqhtL4GGORLhvdoImXVN
MkLpTB2aGjoxoz+mfEIKzwS+xh3/ZyvgmbcgrG5c8vhy9Li1MhJO/4Y7yA8zrJ/s
g+ClQticyvk12OIGF3D0sVQhqqdCFlajqZ8fyur2WcGSEFDXfob9ywqVy2h9n+ZQ
8SP4DkXa9/tTE/Q1CYrfQ6Vul4s8X4lCLXTVyNE5gsOgVSsqBCG6dES0bxkuV6zt
i7i05gxuan7+KSwT8JwNLUP8XrXJFbg79/QWMQPvAW+3TbjdMBkpYrPAhrptQrGA
/UaL1G0+yyOBknrPIGOOSFkJPiUhndEwxpm/GN9/66dBGnGpOiHUrRQCaOsEC95I
Lw+cJNbqIN2TyDstapYgjXACIaIMyOFPZzyhwDxxuK1tIWY6GAW4MO8vY1OFSioI
PabNP4Y/WPG3zuicrr7cdfuRcjl2fFUgCeF94wnkMmET26Nhjc95yrleF1l1bzYO
7uf9LXC/rUHLwAUvhMsNJpZ/AQQLHYYECHrrkLywf95RL8zJ2J9mghdCVbB2skl1
mjKeyCZ1uO8J7cRDmjPv4sU8w+zHen8oKdZY5TgcKiFSmu+47wNkfgeOWNY/mRJi
0Mi2P9fMHubxAEo1VkW0lFmbrb5hVgF6AH1Zzm91FbKF0SghzzNRGjwbyQtNfIo9
lWARWzES8Xa2DgXcsXi7ubXPDtYK8LpLWeF0Od1hqcJv8isiIT7FWgBfHXFqYFeK
m6ZZOHpEkwfHnxNvNDPM7DN0tU9B/nWC/HoAolMjZ1yMpo16qynmLMt/uEni3QRy
Gtvn0STk9xqmtbJS6cJOXLp32vv0UHlRiotwqyNMaHU/vGnFChgwXkoljq8TbfI9
jq3B/VEQV9jv+ysykHeDx2+hheyLTBsCoITAfY2+Tol5J3Ss6EV/KekIlo5dHsrF
p+eJs3XQvJ/p6xTrVblUdiLi8RdABVmXX9xH39sbDWNZAiNdBWXaD5oid10O43RM
+mH7oop+6WprPMJhRDmUZG7InB6mrSFo7UMpQ0H3YRh4s4nrZERmJFySYvMst4qz
tvHuwjKkrFo+3yIA2xaqlGwIadSeMkYud0SzMXavJrlhs92I8of8bhCmkDOj+SKs
mEja1dehV8fqy+pVoans18YShfnXI/tUULpuIkpUCjGCEC4yuCYXPGTlp+7F0Acv
Q5xjEV5/i+MTIDzPfeQhU2C9z79wyCkOgO4/5xsSoON3hjYEE2FO062gb+KXLik3
ySKO0Q6pZPVU6Gm+kFcFHZVnBO153byipNOuv64H0DD9UFhanbTrfxCGnZ1kO4oq
cWfdsvNKhKd7Ok5Hsej3Jf6D0hLq+iM7j6/h+mReAXez0R0ePlZaU7/oUBwrZYoO
u6bcv5EmH2/6eV4KvKBM27p7NTnu55sEKUeUxVvjUsJMXGz81BETfbQSggNOVuaT
XPvM4fcMfKGHeG074nSN/Bz+yVhFzc+jstc82XtAh1c679e929F73kCfXKk1ysof
r1zIaAEyDi+2cdQHp5yDr7UFj7IM561pQGdbm6h4YPsQGQuULZItr2nalv8PyaCv
kTWxEqW8u058yEB2GANb9NE6eeJJcLbscVnYO9/9FJUIfpQCNmN5f6Mrk5Y+QMD+
z/uMDbX4bxJ9sP+dHrDXSYGeYQuefJG7p5euSlk5vRyOBifh0FLOwt5SJRH7bFVU
jVE2WIbrWrHKs4NiMhKNm4ln0R22Ml+VE591hl/jiUcTY6C4eFJTgzTuI823g6Vu
pumIlxViGdWX1d6i/wJOKYJdKvJWFAEqhTowzZzJe8FVk6p6eyyRjP0N1H8LAOFl
gIHOYAqNp2XggARMZzOsmN0HBq7UT4+e+e9WXdkyLkaUowuXkN2YEAAkkY9QMphs
CJSJNbO4aE35N9sA2tf6O3jxMwq9t+2GwKiJanHbq/tRsh1C3blST8LZBGrLllVi
DvIjXWMIpot+bRgMZQ4boJQQQ/eKi7L64M98i3H7TCT3Woe9xs1hal14E+2u3IEp
EwsqMY3rm23auiCys/EIaBmiwjXEZUW/PtslEYRU0FEA1aGKWANiKWGujv2LVApW
/k9p0BuvkJ8QxgqjJj/JNei7ot5kE8h6GUXkDymRpD8r5yeEo/TB4i1It28x+ewb
irllmK4SkL8Obe0RIgq34HftdXt6wiNz7Qj93M8fVlqF7RmBtJYxPTpGQArJjgcR
glhS1Bqbzzs5DOT14EDLSykfGkEOzK3Tn7px7DEB79F/G5IrNGCXCTEbsNkBkesN
SIDDbNb/vnrUB+IgfwJn9PP4wmWKuTtJXLz7Oqs/vyHsJu/y8VWT3zoRGAx9WuNm
EfExaP0TqPoLNHGaYgaF1KykL4KQ2VjKvYAvTDfy4LRW27NFs8pjJ1g415gZ2fDb
CHNf/fBr+6P8Vi32qxEgL/S5wYdb4Cb/jk1i4DNo4NThbcM4GXgRHfxepmHhvlMi
WIgu0osr5jGlVjBbTWRkltrcrhfcR7hVFDWiwWZnYnKqwjM/kl9JnWNTvlpw/b5u
vfSliKjynZHOV6+89IrXA3I7D7rztnhmY38vWRYJ2nJGmvIshokFAhRI/A/tVW1Z
rNbDvcm1pI/PQDNBrf/cyeoqriGfv3Jd9yApWt72+TFam7FCvsenvIWmSPOCSfjj
Sjl0vJpfX9uw7EmlLLMhXyUTaZBjO0u8HhvELQMeKxOsI+xJm0lp6VTz+JaHgB7q
atBfBG1khttkXCTYUbHa2hMsRT0wyY5m8yNWge5+n8XZLx79gA6+BQvWZK5Q3ueq
/jMhXuv0Tvx8oyGm1Ey7QRjHMRkanTtJyDAawWRoCUACyqzDMvoTjchOJsjMBzd3
UqCzWM72C87z6XYQFGgYmRppwJr7fuGjXn5oqV+KE7WgDK3BL5HA4U+nAjXp4mLX
FE1j3upDPPW9wzcHbbxmD61fIPJJ01U9kTRnuGnLE/MNTq12VU8OmDMKwPIeEj5P
phrbGfO9MHjYxItgYt/GD1gqfzdiGkpQSiQ3x07n4JalE+G7ZpzIKEuvU+e853DD
wDIX2Ju7qdTiHsBCb1ZDnNJbhRroS8Nu64IhphQ2SZ79AAl3XyQrkf7eF8u3Oeq0
qETcy7F1hOs87IpQL+JxF4lz/OZT6ndtYBC4iyS/ZKIJlzvl66bTMwPLQPAyi7Lv
5Ij/kyxWFr5XSXWN0b34sxF2xxDAsl/PWDBYjMzK+MDP1X1elK+vQXqIukEdKhlF
79Ec8rs0Q9ydziD52mRo12mua2/IvWT3pcyAmPhZyjh/0Fvh9VeTRxOy0pX+ZmJI
bO2w6VkeVmOskDyhGTwf+yJdhbs6obSjwe2F0nbK4nQonEC4YhCMlvVhzIklnS1y
GxBi2ZvTit/sHQEGmxreMW9G6voJnsYFBQoWAgvRJnXmIafhPBenEmIhMoFHG2dq
VmgUlRlNoui8s5JcvH8QFd4kfzRm37Yxw4Ip15y3AlAMP9aoUjHIiL4ol9XFnKsY
501Hh0QPDkso+qkFviosm/Bxw5tHfbj04mfe+EzH/9Kd1RIKSvpHzrrC/zNZPIGz
hsB+3KSdPEQDwVBSaINh3kTgyPZf7ApSYqXG1ZEpCYYo+qMsJckeVMHDu4e80QBG
AAuAH68P1Hg2j5e6WScwGz0Kw0SSloJ4f7ODsRBjgshStxqVDMEd7BPUj9j6SEpX
0u3EKRunQCc1Eh+t+3ksxm9Un1VZRHkkJTQoQIx55p0JO8EGHmTBF895uWjQXOmY
OgS/UgwlCFF8aGMPaGLY/PJ0WWaIKtDdP/++eG3rzwZl2wUsxYx1F4Ssf6AHavu7
t/VA2mGXTA0XbVFsrGgbwIDpluIOQ4MauP+kLO8RpTpEJsViTzCHZJgxJ/3MFlcx
HBdG8yKWafR3Wo+zD1v7wbYjDmoEDVBnHMO/TQdqd/D1Q8zejgcbh5eXSkAyF693
ujCa3SeQ6RhWiRgyEbrNJ7QYoxL/yn37OADYSKjODelJ82pwwxp/pGVdX6JCnaq+
/YqzZStJ4JT4XbojJAo8oXn1ifh0jKDrhVHSPHgTjwsmSvWQIJHY8ok7Q+SuyRDk
fR67f2WVOvxF+Cvb9d0zTsiFkAK23e3wsXoFZx1/X3YiD4K4J/roZdYrzfgJLkcX
zCquAntZOJO7hR8OvlqxVYYck1oC3tTdERhmEiypiU6SsL5/wysvcXCH1RKXQsv2
3gopcGPvGaGX6US5PfePcRKfa2xwpsQu5O19/Q8EtbWw78De6lTpu/j2SxeybEtD
aUFyzx3Ox068pdBJduFSbg==
`protect END_PROTECTED
