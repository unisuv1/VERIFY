`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HKejiW1pIT3cH3gMpqWoa0f8j1+zbHWu5upPR74MCQxHFQOCfHiN9VZs1ofkfJnY
j3gQn7wNSRxjAxSWnfJYovnypptWShi94V5aHGLqD0IN1S07q15NmFarHVUVwglP
ZKxrS+k2YbqDETB1H/uuakrmhIJ0xPzNwVQriIeDLbtHnb6uI33P9ChqHch+kBSS
3BhbAY8O0iB9Jv22ei0VOPZPGbY059jbiUXbqmAuhWaVApuF922bGqF1D/IqzYKI
MSoGCzl8rr7nQz0Nd9Fh1PFt8B1vSS6UZ6fggk1PSQFQvCTB9oHoJrC09V9+G1lP
VjQDrZQXj8sPDbPZ1vkkg2RwMV9JkX8W4jM8GP7lF5Je7It8TveV2ausy9j3YTK2
f3IijCwPRLJhMp4wGw83dxOCo5KF9jKvgv4bGvSdpj/SV0mTdFvlF7jPViVNQfLN
TIjG2F+Bn7b5jGRAWEuucZqNMECVBca9dwrpJyDRpwPIN5YmJ4uLtHvskIau6/KX
TaQAjScpyK9rRYk1/ankFvVbwV1EZHVQsy7G06HBbKXVCcd4XXUN7im60D6mJA6V
7WMqneZmX+CZAAjl2UB0nXGrzOtht0CzlmpTSfQt/pIef/nJGs56niWh7JHBeK3x
oP5YWwy3BndKXl8MccFukeiC5MpOfUBEq3A8vb4JfYshkjtuf9nrZ2cEecLiD4KS
sSHhmWWDaPByM/ICGrKs9ibsjEeGZQSFNocQN469CIaoMAV91uo9kGiyZHBozJKS
iB0Q2Z9MqBjRKxFWxJY/4vAMi2s2v+g9rVYsWXcGf+1NSljNdc8DjTeuxiegKYok
fhrtNhHXAf4ClsbGzp52fuzGFp2vZvCpf7EKVd6wjNk21o9uruSWiBRePsgjbVru
R54sqkd/RmNoqU/0IThmOqInWq6g4zLuH/D2ieRG4GzVD+c+Q6Cbvz/Vaqeg4ffu
hgzRq8jPiO0dymWiTTeMZ06jDRdSPxBctdDv/YWeGO4obYyJx3YsGljBCh38QFsx
ZSqCpc5ljPUkIWNCuUpa7NmlQmzq8qUtbXsjd1KpbMbC2ZilrOrs/ZABw6a+yb1i
GfCidoTXPLLhzbG7xnRpD8Af+1oPP2DCAQGBSTLEVLI8g9OL+n3h1J7vJKWFHLEq
WReUfS8HYpm4XHPWGoVOzD//l1ojW79ytKg10fM0K/2dc7/o2z5+Ae5PQIVMBrbv
RDD4YH2iRAy3prBZqBFEfl0nccbHPMCHKkBbFjaLkVeAquN83kuRzjE9et9fAvPh
HxrnItuoMX6Xk1PmYgOIKDkvtvEhzTTieTBuXVdaOG/K4bfr/YhymsV5nGmMIBcF
n0o6tSxEjZXN02qHs7dd6bnhWwcyhLn/AnGN3JCt1tsJCixRgmlXEnRdcjST63LC
J2y294PP1vZdnGAzTGAjGsPrUbE/wCCxHQM4NO94Mu6kL6Sw2YTbByRwoYpetehC
u8TKUsotiGHSK5yTO86zZWUPjOnHQtI8v0lz0xfHzFeSvbeEbKKE0bDsf2N7xY8T
/FtJ92zLgGK1oDnvGjH+g4LDWFY500n50FcDxEJr/VGJza+OYM3OfvAmG+6NQfCL
2AZfIpzYSPd6J82YQVl2g9VS6HC7RBXE7NSR2+1kjtlHDuv81TjKwcbsVY3LuYs9
nCAjSIKRcA6yFeLWC6H3//GpTazhEBskbhLkICYwrEMyaumgSBI/24Owwq/C94kY
s4UOMwg2c2tHZnbfOxKrBj0Ba3jqiCFRPDN0+hQ+JygUirO7T+lPqoz+u2VpN3+K
StGbZa5NyLxxTY/CvUWsOHjvMIh2uQOJoRmNCae3fA3b3v21pJSUdxBnM+b7JKGf
wGXs21KJeVk7mitZKir3Cc2A+py8qeru+vuSERIViobHtB7B/4AOf+ib2sdhj6ku
ZuGm8sgK9JrF+yuSBe73n8JhvFhBuFDWJsZCBHnfDKZYDxYsxmfPI6aOGfHGw0j6
ETQkQC3No2R/78kut/uooV74ApoJqrlLwoOMoAx5t3F3+Z1FYXPD3DIby3L4zh1+
2EnRTDm/LceXJVuYJ+2OC8i6R8RefXOHCxKi6Ks70veUG/5YPkIn8xjzK8xIxwCK
EdfunOCveRss7HA3YumO1NzgkkHzOvxxx17K1kgvwBEcAZfOhnp8FALyMkzlKCsF
0LAnO5prYL/FRnTGM4TFCAKV7yU6AtGRBWAfOL/1VHvsOBTvc9l3CHiCfi6h66Ui
caVD5zCTAUVG8dJXLsK35kCq3vT3coKejZY7CrApazn85JDUZBlUc6GJ7t7YEUpw
bp+I7C4P+jwZrtGJM/+fkIJXkETx08zusB197EcEEloy2/LiO4jSF1Xn8fscLwsV
DUziQysXLjWPhr/m9jlLxTw44UdhM/Zu/d0XU1ESjA/KbxTDz5cQhf57z71ZLavC
zQ58NOeNZYZ41LULSCDsdoYewSf8tGTT29IHwYp2dPTlFz1YskbhFEszI1TMnxQ2
VP//WQNq0cf/pLnH+64+qldWQdZXDUq2VfOdfC/Lfem7dM6MMyj3g7UIql7eQ3Yg
m692NhOWdKanoLSQdiBQs4X4VTm4IM/NcQ4gFX5Dvg5zSKkCVeli3SU6w52bqyns
F2NA7g8qPkhDl2ShrZWjp6gybiuAmCk6ViRQe8SNTt5sv02NymKu/suXFXTobGs9
rPkRrUMFdA3iF3CKbEx0tueWqgsIag24EQmkUBRk6ob3VCHWw03y7M6TpF11+3SF
VYc15Ib16bUmaDWduH0FdGbiAzeWZ4aXtW9gl5HhF7n8YiMIJirkIlQsmmT/dF4k
CrG7soQQiipj+pHDiPfzDNe8K2PCp9Glyu7Vk57sTa2yiN4AZ8qHvtVEOiTAlcY3
wX09cUrm6upk6AJum7OvAcvxUxTyM16JxPYBp2XJjCm10NQeqPfk7emiesgjWIY7
lrw+FkIbBLcXBrbbIYhYQnhfyjlhbySFLLiUjJfvtXEw44a1b8zEugfNQu3xB1y7
bQjLwOPYAH4tPqqE9J94MrhqKTb3Is1a3WVmN8UHdItBYPSeF8nrdvtRdoicbmLY
B2WgRUEIl8Qxxzevmw6/L0hEGS0ASoghivFNPgPbUBxIgUm8iDrItaQlpCzHNF7P
Uy2lQDB/bKujSTrZdU23cO1j/BxhXSj3vdmicRIHfDbNkS1+1cSLo9DLsSNoJOhK
k2gHY2Ga0je1GtCHrclGHQpgzWREAD2uz9dVr6pnXgWc0OL9PNerCyf6O+Y3X7wL
MATk7FBbbx4GORz+tuxR7Li+cR9y6rZApN5YE3OpTFkPXDO2fqDJ8SpkBlurZfiX
mnXXvXEFhMZOB3tWlTIr49lwXXKEbVJaE23ecq5Rasc3e1zLaXS3p9ZSWbZMNMRA
hCgpY7ZoiVGy/rN+Mf5tgHPl9Q6zaYzViTjf4aEg9P71FbVB1PLsSonAVvrtnR6I
c7zFG2snINXpEV/a07PcH9OgFwLXtwEw/vQ7wcPsMGXxpU4i7cK5EcTJvdZIjfWZ
9S16hiPiU1qHqJPytV0AmsPX0f3BORkFshc9RSAayQHjnnKp3nUUiYwMoIuaXw/t
61YspHPyxwt5kclIC571ZH88ehSmXiOJ/QswOK8ipJqdnXRNAHIDstho598s5L32
+SjzhV62RV8UYZp+qIW3DQ2gaQ2XbJhFRo33ZMzLmyHOaP7DyNcA5YgCQPtDBtxW
BVgM7CkxX6p2xEEN8oxMgKsTGpXFzW9XwUWtdIO54NIeYRTF7n1+XIDhZ78fGYkH
LBC4LLNEd9tBYGfzSGf4CElIWRs4WOCJ7DIm1+2VFx06cTIOOMVO4srLsaihjbPO
j0R2Ipj7L33JdAhRrUeUo+R1m8Aqpinwq4pLqsQvcgKY/J1bojyGVQP5T4ZaMMrb
HUmJjufi2CjuuesVsdj+uVSB5OyTOdYh/ZGCKSDeL0OYJyjkzat7qiv8e+MOY4Iv
2irLLHKSsy4sPOj0e5zNDCpOxXGapXx8hm9tzAQihB7efQSTvj5WRqkCnv9onTSZ
hhYIwNol+p2rLo1ZxGgW3Cn3wWeAlN3UiL+b/wcN8GS15s2IwEL8/k8TMNCtvrFr
pBhSNcccqIup5jmObzDzmkqt4LrHZCbSvYSKUaDsfyvjJY8rj1Wl/Kis15NLcafZ
0OPGwnhBKNltlhy/luZ4JxPOF7Jx2HM57XWUGokICmFbiHPDaseqoo1m+BbTek9f
MAJoQaTMDIHV2caIdGBRA6x0EaLdvsNPHJY+UkVWHCBcK61FDLs9knH1XhjE/gw3
VdCl5DPVMB3RCAoSOWgzs6shzXQJkUC0gbQ0f/J2ZDXCJffqc1U3zu7KE71HP2ZY
xx5T/Vs5eDOJR+ADfcFMmO3tvqZOAifayVBU1yhFys0/q0C7C+ihaaaufmr1V1wW
/FXlWpfI0KfyJcsbdyVJX5SeeocM8Rs7mEAr48GuHMxtoJQ9uxsw9TY2RN1rPQzq
TN3gqYkv5oECtL8UgOaOb/6vYS8MgWdLsojVNLvf3vyI155CbijldaKo0//F52yd
PwYp1aYbk+gfLQ+sWTUVXNkiLsynOcAmD5vioNv96KI+PwGQrjF8ifPJol6w5Z4f
smIoq72HUyozkbrRQ6XSPcV0/tZUEz89C+Kg/3JXUPEUyk/TObzex7g1Qq8TdH6t
+uH+IaSzmry3eW+UNsdZnXp4gLP4V8gX9RHbQrZxmhU4cCfFlZrYvl0rIhxhZKlB
v0bXYl2tI0zkdLezGrWXIom8gPjbiks0uIS11IvDYPAR7cnFN+rb8rODnsuL/MGX
PVhB/+5c5cnoq6LA9yE2sEKiEE8m68c9JI0zjn4ts/XxIlDMAnnaqTJF1H+aRSDK
Hana3Wfk25+AM3pVd503M8nLRNVTDO9teM+grzZhGi0/SF57ijjOnqKi99hYSkBP
m0mpl6x3Gu+EA2j+PrzotJmh+LKaSLrp2KNVFn4KCXtNTgdTEN/J1Azv78flhRm/
Xnet3FcMybqq48lwFwsdOTCPj3wP+lRKZh0E2Oh93Q/An0DkSEUjSDvIE1ArDcmT
OZvbyFcyB/90WdyFuvhcbtrV3AjSnyJ5C4dWps+XrK7v0H4l5KAbV2sPOSUpi92P
Aydu7tQhaZXO9msokC1khJSPsSLSrA/iotbCuCx//e1+melh/BhVJc85tFmhEkbx
RInW0645qS6m1KV/V2WzWPzsUyLNsMNDU7SSND6KUqg7VDUpB1K+/42EKMPTPfoO
ANSOhhCDjjZKoXuofRg4tIT1Q0g0NnKnji73pxvmw0yC1ZJc4CC6NU9TqzhOp7KZ
ObP2H0XDNiyVhMh63vzur2YtwlfRYdHBmWk2gKYSqmuxqDD+Hpqo4dSqPIVkMik6
4PsdCcSSZD/SyCWInerT03Hn1tbCTDkOG8th+cczVJmWdV9PfRTNXDWvlw8Ke7XG
209QnBOHuHALdTXv6vy17NlnmwZ0pd99zpW4OxHmXwq5ShA2QQwHzYgJ13VVVEaN
Jci9scmrS0/CnCUT9T/6cr7F/8uveAmJGHRGPaAp8E43+6Qc2sGuceUPWn7QYwt2
N8ybaoaTsr5hk0BQi48O7vA0R6rA22QtC/oQgmsE65qFqJM6fqOHpMqfb5Z9gl1Y
cvxlWn29Hv9c/jkgqQIO8++I5BpPgAFFkNGgNDZo/ndwpUOtYVOH7hP4N3Qx1+7V
Av0cp7wXHbPzaKoILxsbZBOhWTxmp2Kqhd/+hL5bc80JRqHavGfTLtz+mZnzFKDg
oy7/xd3APeRsLrs0poR6m2iQsnMYU8nDl3h3XWVwkKc6t4TpOzJwbb2tnAo+nw98
n1m0ZddSgzyWxDUBEVyzJp2kpi9zZrPKwdGsLmfuLnSc1hUpIZfNbKCdR/xNjmn7
KugyFAYlnUG6WQKmHt0orXtU1uloZU3jRUBavOE5Xy69DkVO61ClXG/0dI28yHy6
7N3XF/58waJce5s+N0N9hw==
`protect END_PROTECTED
