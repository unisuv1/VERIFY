library verilog;
use verilog.vl_types.all;
entity tb_vry_BottlePrint is
end tb_vry_BottlePrint;
