`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TSldoDPG5afSKGSAv8vkH4osMwo+mnJK/eilwrIgBJpb+vo3931OIZHk3YXmLKk0
Bw+aKQVdKe7FHzgMUU0AcVPPrM8f3nr4h5r5x7LYyE3ePfYjwOPuCFxerh6Yp3dz
5fyPvSTHqnV4TRA9YT9PWrzMMzpjUgHEPdH/sRUef60bgTqyexAt6OdTfzu0H9R0
VsJpxVvIyNy4a1D2wvF/7DzrPyS+Yx2rK0mgkoHblTdeo1LXqT6e+glSirVCfcbO
Eitd3jfc+EnGdPJW3d47aQ+83YO17nAJPenAze2wIIkZOBVJ2cgZGXm9H4miuvie
IpLv13lx+5wT6+6nbWIhB7Cnm+c4RHTzZkSwQ3Y8zGSQQQKiRlT/cdrj1+hlEZPr
U7tP6ts9Phfq9UnOBqISp2BZ18MiGe12JRGwWSIdJKeJHqJf70q5B8x0OFAskY4X
edzydpf/Gc/afBIc30BxXdS3ocsANPsq8ZQZu7pDn98hv66XsQ+lrANdB+yveoRb
cyJpE4GtoDHeMG6Ez8ptykL01t8qNwNx161b5TJiYNfdvZKkvNFy9+YRaliPKn0a
GWSzF1d5RdOhRDK69VlLdl9rrAy1qCcRuDI650FsB0/yhGznTzMR6DZSI6BdfAVk
B5BlDZSZatKSG4iAurRAwTYCT/VruzRJFvkE+pp11ssXWgz96ziyot1BODRmd76u
CO9e4mNv9oE6pu0mmSxhN8HaGIDytskhhWI6gIGkSa3PcNap6CDXXVJx/clSD7fp
uQAy9N5VGjXeZlCromfKEtzF9ldLoUq6gNo2FiLHyUOcOK00+YPtsAcibvVKc/YY
YxGm2zUJHdAGokCOKe+zmsZdI9b/GKAAWu6wOOmJrAvSZzYnUn/A+ebzgjQnNQUR
hns+r0uVAJZH7rbBOHgJ9OdNg1EjCmX9iHsPq5jiEcD32vsKd5HUbpHpSH45R24H
6zuDrJI+YMkajzQ7ywQ9RltTvuE+0hNlCXGdkbKVZJWDIcW3wY8RUTlpYJW84yno
W0mPc15JdDcKdU9UdH5rCQgVWFp8U7Wbl85em0Zo+mGNTbeQMKcrRhj1RLs9DqB0
`protect END_PROTECTED
