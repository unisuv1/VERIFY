`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mEVSlwR37ZFvRxJXI+yayvWFVYH1udCmIGvWnVUH2wyUSH3geNQPy3rbdayqEtko
2a/D3ODD+KFnsvjZiZ8JpXGW8hKDTxO1oXIPlsBQzMbGgwUaOgfMTrrvbhKEeVWH
WvBD9+Tis5ERshp+oUQ59vC0t4/ivVCEiFTx0kOYq9PJkNN88LtdBMP/G3h+QzaK
hIqYsxjmYUNp3WozuEQC1kRGmlYc1om4ug8Jgl2M+21PXaaB3eumwon8Zy3tBhVz
NyfEYiEKhaKSBkrZKJiCDZt+aQKWV4FYuszQhvDz5yiLJ4O3ztboGlaQWxG+W1Ik
9P6FCg/ACaJNezPtCc4yGyZFp9bSD3TUVhir17PVPmmjFeZyOMn3UkjRNczdPQY6
+vqSfoKUKWzNPzPkIIKT6PpUWjew8TWsj58CIdpj/mh2l9D0V9jkYjs4N+E5N1WN
e555znMutaaDWNMUF9hKa83bRJNRiq0O8sywlUNPEIwNwFU37+WCTeBwc1yo/ZQ5
tRjZBUX2AAZVyatMujNHlHJFLVVDs9EuVYvHQxKAYxWWYKUM3Ts+tp9hF1RsZe/y
QLdWb9e8Vc8obztibg2OumdJwQdRQx9P0OUIcb4jA/mjpejoErCQVGoDE6ANPWwy
Z+tHWJL0ck5QCg7ZG1IXEVNKfFddeLjU7P43TdavS0vJNmCF6Q0E8IHhL5z9xA0j
0Op2nv5JMfuX7lnBxfwPQ4Xufuv0qBgIYojwTVP+r3p211nlBj3Z/InjckHgya37
gdfT6Q/QBn65ze150S1gOuJIDp/fL9Lqtn4ms2OdQcdmt9b+2tLMKDgKm+ehB5A+
U9BjmNbaK0hKV4y2bO3isJisgFLsjATMYmN7lpqMq+O/hlcO7rXnSoeHJ7VsOgrg
W20BtghkVOtG1KM9ThPOxSUBflee6wLtAPqPY195Q7HeFyuOAfS0N51nNlyo4OD1
NJp5n3DTM3P4TvKhvDUJnDAwTNh2FcxmKNI8mJKfbmpuJgbe6bEYWw0pvARZSd3c
n+j9++7nxnR8crgbg+ttN2iVv1/jc9k/LBX+iPi8GjIy5NN0tkqryWcpnjH1SqQa
3sAnw8KN4SeenWkXTfV7L9yeigsMkyA5KobPmFYGO+UmahmRyXE63s2v1IRx069o
FNqmw9rSSqLLry6gnrBEjmdVjXwdlJw70LYKiPo764QKSj1s3iTrG4pUC+qT4rHX
zElGv0WevUpsIqFKbScuoFhsFhmE8JtF6MmVL3KccIBIuwhUYJpjdez6yE2bjLqk
YESijMHYbIG/iDzqDGsnjE+koBKETkq3OczrN0zp+wZFDoPx77vyi7yKjqRS901U
sjfj3gPlXNVULXJwBFtCvhLSGS4Ayi9wKeqiSINRwxkl8PGHLlzjd+mCNPrzTihM
SC2IBdWJvvAddNgVA8syiOoN3679nBHItfs9DC0+nikNI/zVlJ6H+pEplDMVgKUX
XFPGtLkBZF592Sq5BpLLSnTESpSthKO0VUUltV/y1QHVt+lD39Ji2eyR4tikifwV
ykeqRo3mAlbvzrWyjIiVjLrwgZ0WlBFJ25ID2moHBmILdIm2xgkYdwOzGPoYgirC
DKgOP19dk1vUVCeAIQkUXMUfozO9b5HI/lTAmoGytKPb+gq3Q2Lf042Vzsqo3xRT
lYnH1TIQk//YGOjrCiJmeT/Kno4uXLenJuKjM/Vg6qw=
`protect END_PROTECTED
