`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AFGLkDLuhM+ZW1mVMIlfU2tlXL3R2l7SoXHSiggvinqf8I1UVCstgo/HGCu7lQaj
58cKreLV1GRmnVRn7z0KDsl51REMUv/PkAaIZ9Yg7L5IEibR4g535m2emIN3JY2I
Tb0f5CDj1HVRAk4edkF/Go2l2JLCmWn8XvqwJF0UK2JxxWOOQLoWAw+nPekanSvN
LUbpDdn60yIF4CxAvz7yU1n1C4SVzftUVh1AgzvME2kPkU5E5Fhmomr3s0mgZAqX
oc0RjDODpI4SWvGDtboa1W0G3mjyMGpn+SmyAnZ9/7rRrS+RuJ1TzvBk5Apu7TTq
46lvpXonomaZH5ebblFcbymFSoSh99bRj/0PrI9Q7qKVoW2tdS+JZvmLwoOtDJjz
z2NDyMDeWOHE5lA2B6xERac8IAEL52WltIYMJze7+kuiiqPrQ2duCjRVWdeVCjRB
G4XHBSCwJpkMMn3tkVWmXU1VlOKCg7ejtpQFh2HK1ScLZklGepwvw6v6vNAFUUXC
zIiopknPqVgmFU0NoRJbw9gZ8A/z9uPIVRyiv8aY+kRk2JXN7apLXvWU3riimX57
QYjyLZFnV3Vh/0+ZLrN+Ffof+PqYY01YCSvzYnnj4/uggQNd2lendfHiSJ46+cFn
a0WmA4MlgekaDCcTVG/IldffLGlSRGSC2tuRnxGUEjhXE7czz73jtK+P3yi9RaDB
Nsa5dPqdcaIy4XO2fwC9TDDN6+lPirJ+E8aaB/JcQIApg2awil/R5vIKWU4S/G/v
2hKP9roSlnJtv0eEaOP2iDq0tlR1uZrtrwDR3cVNqdfSvakuCqgalbTmyPLmsIOy
vSGzDXx7hwyYY/YXeQtSayCO/QClwbO0v7EfeA84tm/7sJD84GA06yYdN/WqXcum
TnlzRfDOtDIUtoGb8fZ4R6G3t+STEjivZ/sTADNCVunpLBsBxFdZie1+Tqa8znr2
XnHh4gAVItweDhcHjv3G4Ok0cTvFf3EoMB8mmWtCgfU6aOLdhpOINRsD6HvziGpb
Z4MJVfYcpmdBQH+i9eiRe8UPeHoWXOQIhWglDghvR3o9tUOqbrUukfBBis8p/D3j
tP8i+VHygt6EAUcGtwxUKOLL92NC5ZcE9vZ5h7FSaQd+eUybTXbe3q1s0lrQazkJ
2zJ4dbd/pUgH5Dem9a1Y6PX0uIycwQPAetJb0RTS0urdeDQPcMWh4MjDlc5BVh/B
iqg8P1f61d986K1MLc1DL2mzPZbu+gfcNfcuAUSTYucGlD8Jv55UGhBJPYZuJ/fi
7OiRNuDxf1wQ21LqtC7DTdSKx+JSHLvHNGfMmAA3CodOd0u1TYHpoDz36cvyA4eN
amO63FKvGlqFe2TyFWu0Le3Cj78hEmq9WtV8iB+mLrYKE/Zuru+9qPCbTsOWgneM
bdo87TgwomOL7Znka0KY4jh1FlrGHOMO/WjY3dy39HnZbWBAqhcKgWyVfIdeSbXQ
yA9aXZyPvJoXWMNeEfSnHbqvMC5ypN0RMDPoH5y7kD6FUss728m1DuLBViO7UczI
hmf8q87fdNb5KK+bubPL85OppBSJ3wUddFgTRl14CEZcApQgRQqgX4Ew8SMD6UmW
Y92Y54v/eb4bIioT8O/++h8bQbhGkHkkYHDI5ne8ajXy7LD2UmPVqDay7Y8zPAfs
Cp6tg4OeMlL6j/ZkUAuuys3QkFsbIamnmJKHf/kZMhCnq05c437J8Z4fWOgOiJE0
KGo6hCGdebu7dU9x95WpqWgE7vUqSXJEIcvDIPTsxGEkWVrMbWFkACEduMzdcOPR
GvaKfezQD+N+yloYKE4vf9O9sHASJhSruI7W2GGRvXj/D/jmTRRUAwWHthIfvMFn
sCnFc2EZasPDlqAYYonc0/naMQmBpF8oi9tP7ptacmhhvCgQ/dwzxkHzRJl7Yt6x
bDfGELSp4hwYxMHTfQlL7CnmNLRgP8rpDN2lyfp6TgHWZyZwhPpSbkxrEKIxuge4
okAatrLY3W0mqcznPJK0f3a/qShjPZqU1bWtqTraED/7YS2nDYTLjjX4m/s3jVkI
KppXcGg9w4+4r7/7cq1AZq9zh1aJVkSIEd7j/6O7MUHxPqlorIdJZGP07taxwZPb
Zu+ju+iNJbmOYaQGlelAh8zqcbnxWD2E5KZMP7NVSRwApOzjdMDyzKOzoOMMSQkF
wNHs18YfGEn0RUnZfxNYuCuNjN2TT5D6/1GEWm4L82/eaPKAMaH2PhklWt8vApHk
aPkrgzIYMfZ67R+BDqBfmHFZLVtiPk9gw2oA6mFnqaanU7tB7yK+0uYnjRsabsjI
bEasSQmGFbJsxgIau+LMQw34mYP8cLFY7EoQn8otSyD+I6iVREhRBuO6Jypc2jjf
aL+/k1TLhSrOfzDV/MRHomBkwQ2PDKRWoChHnUgbYaEL5oqda80eqcDBNrLzYlPq
drSx8R80AI1CG15/quf93tLz6sp5f8FMDw4Tzk603AGdVOWCzBrxbXe7R7U3AMmG
RRcWo8TS96FKpsZjtIxSIljYUILAdSsKmZC0bVQqsTiZ32A/xIUuKoleeiB4Hvgd
JZhA9u+sYI0GnF9tGfoNQiLTXE/KVRZH7LkDap0OGPi/V0K9VPmm2fegP7DwYInY
DRU4zanewz/1nYI+ymr2hZQxLnIlbemWeh4CUrfeQ7Hbc5vHVyX9o8TjK36qTBoV
2tvUmalBpZJSmIgvLDaMVd293J2NP4zP06zL1BgiIgBrlDTwsWlzV/AMeDdAbvHR
vBjQesoxLkyjtsUFce0S84ew9kUBHs2yPWLpn0EZzhzjRaxsCzBX3m+u3TfpUg4C
aw73q/DBKlx+YBXcoQ+tYnmHj3ZrXwkA2nRtTwTWwV1pcuNQrdDqSCaicft+oFvI
HhzaOeNiJq5qUeKp316NLDcOcef8tDct7/2H/SaGIlrOLXWKibs0nrlWr68SeGp/
miwGiVMRbdAcuySW1sYj1uurDPiXavQpa377M/Mohr3J6qvlwgzS/5+blqJayp+M
SDB1zyBB9ciH1vDl0kiRbt4kbXp2+nfbxh45XTrOXUo/gAXLzrE/eJBR8QQYSHF1
93JblFbUgdBiRX3pD418uICL6/mIfpYmEQlNo8/Z4oKmlXwCrNbjRlgMw6pIkR/6
IOezhDWmQLkofq0r1D5miQn3+6YqixO33GEHObbNZqDmD4No0prES+0UgilNvJZ2
JA0BDSobeDajJ6j5elh6Aw4R2J1rOiRFs9kmV1Nstbx8e8OsBIOHlrnxb+GQ3jR8
htMA/jN7OIKEFscCZGYEU+zgJlAbHjvBJFVXMteVMBgcOOHh2KdpE7+KOLTwewTQ
OOJSXauLU5Iz4C756mbFo2PJiXR2cH1IxmAR7IA0MUXV8cp2DP2oVu4lBMDe898G
M89rY7wvXXdYYVoAk+AapgIAvApfL+jAlcOUWvVWZ0KTOJ6r3h7ouYJXFUSQhsSz
KIUHGdCBSUiFXw0zxcpcP0OHOsucb2ax17HFOchLOuApdOgQ/NC86Rp5wrWXoB3s
79ccvj/NKWK0ssiXRGwBZ8pSOYE/zJZGQlMQw2HgdCpG9X1vlnup0axiPPZ8A7hq
+jx9uhA9u3n9JS0Ri80w0t6fthfNQGWU+S/LPJ3ZTHiHCk/GRHU4kvAVRbaAmDhN
5bfj/fqTa/pxCTGI5R4KnK3IEKMoT71lCMkuHICQWcsPhrFc2Eh4I/tY8B5QGg9M
uZtSsii2puvyzoGy9SL/ueOydIuglKKeuGGEI89xO0/Bxr9UtkTkndIO3vBP6Pfy
6mJ5mJHzhoqk4zLwun4kRPsdIvN2ZnrJTGe64KDQgXdHMICnPjK87TmQWNixnHDN
LfSPvUaU3P7ZoSTUqKy1SCrF1WLJDYAtwa/iRIdACKwEgICqVwdVX/G3vhycGP7q
t9UGnZnTX5v3k0zZ680wwDp1hKt3ndaQbbIjOFO8KB5MXdbUPf3ji2DZqpJxBveJ
EnN8MG78YsYqGrgxpDEVCcbcHickTzU2Av3ZO/9mpVoQEyhaXmpY97iRsJLee9MS
yi/vipglqRX6hC7jsGbOlCSGjXIwbFSmZ5TX56fGfYPXU/gBKwKep6As28BPnKRv
Up1IC/r4ORugdYTugKv/W6yjE+YEZZmM5b7SeBnRFxW7Y9w00ViymzSZaZG87jSR
0uNhrh9y32xQXgk6xTJQEsXW//zuMH9/zWGvt+N2erymDU5zvAosMqNQTQ6dIdkh
GUi6xe1IeoHhMlHeNWtxXlOjdY6/5+HKasrEhLsAzgVgfOl5HVGRUzEOXCYbMoj2
n2lOwhqHwlZrKeczMdCCJObX2Bi3J9mPwl/m1f2Hxwtb0TnteEv5tOTn3cMwTp+N
oDitvZTehmoRgIa8wRiAsfBY4QSdIaw5KQpMkvzN6oo53nGm2iONQw186Sxxl/5Y
d8slKU+kN+tYdXf4ZmOqCUKpWVPs6MvYrLzzuiLpY69t27vtPTPKXkZYwqflP5w0
I8PGh7PRGTSOLb1PB8z0ry6ccMJ06qsSGVMjUVlWptF1T+P9eQsMdSGE4eoA7Akf
c1I2p7eASQ46L9mUkt24WpVFOlOYtpOU7+nur/5CwSWCgJMfhZ3jmIRN+hI9t2OZ
bPOxyBqLd4vGcljL1iEJ/qFqQQrO7fsosmA44VVhj8L55XJ06PDvaVjcqvr/vh1V
EZxgiA2cW6oc3QIWMWwef5iVsZ4+iXmJ2VcatMPPcLdse+jzsZE2FmkqKxzZpF3u
0ibnhStxIHo1BF8XhZlP2Oy6oQBsLbNlBixugzSktdppMtBTugFx8nZNkRAVk0eC
lsaPDU/QVR3us7DFCOdWUFuwL1AFqCy0NhM8Peo0WrstpJqxAOru8ghzPUxvQn9H
Wls/iiXB6C3kQnvQu+K97OVbCF1/DJTRCDqR3JXzupEIO/b1WRaod4vaqdstsUVC
aArPkPf41dgs22mzoUCscnzMEDp2mvjKDNq7MBp9nCSvQY0SGqkLrZMkK6aPQEAI
FU7UmgzAE2tPtpY5DdoOjkZatRNlkDQfqXmyGCmU5eqbGYKRDTTyINXHHlX2ol2t
d1b9CYggK3zdOixaA4sVqh9mqZP5FZH+NdENB0+D6967+4yI04a7520PFAT9Sc2m
cVHymATTPMSAlAs9fPwcGl3m9rPez6v+RTKIjabeNCbNw2LvGPUgO71E56WuwrAW
agsY/RdB7pQ4m0N5RdZXrccEJ8qk70DX5VMVq1IHEhySTssS5LbEIC5F+i6u0CuM
36dt4AeFe0uoOF5VMvtFFL3pgTMAkOFr/cv2fPUDNek1XqDd5pfwLglpLYlPIRHu
kgjZmMUCEi706WLI1wv3gpdIctNCPJpl90FAU5rUFcxkz4F7EFzQ4Bpr7SQSCMG3
y+y46Pli5pnQZyubG11JD8WG5AFkvdKnDLylMfsOoqC1ZSZhQVY2gvhlbJSPQroj
MGhnWirp8/tks8HQPKP/wyj4VD3euTYz7/6eZHmpLJ2dd4Zgedx1dlzDhB/C0rQl
4eJS2YjCyivTtW4SRykYUTbDYzEgKbEh+wuZgypMbT+UGUOMIoH62+i2HlAsGu5R
yP3DtraVMTdDoHrLaaVAHuWK19+G+ZqKJIcHnwPkhUpA4khJVtR+aAE0qnfN4c+l
hnOKgHkjitYUBMSO3p9CWmpY4akXgC4OExQW3IssX36GozuKBP2mbgzLajZ/MumU
D13tO9kqhrFsYMdMi9exS9Ary0aN+Le0VJ0P7Z666PBjGSNTcQ4dk+0eJphtSU6u
fMuD4K5tu9U95PT+xcA7IGybAnZlOcovWcwNw2i4NEjV+kgbBoMQLDoHbnUu9pQO
ox0rdB+OnMaCeloPb+zMp9kxDHjyIn/t7XIqguETd+2kEQBP5kYsOjOF5WyFrT6s
507EPS+SulIwvMTHtiDLye4ZbZ7eEufmwEV9AiDUUHVk3gBFHfvGR52T87HIp2eZ
AjGSiKghi87R0NgE08hjqGlfsu14t6UIXSvW6hZLvveRgYApXB8fIovHo2kpyH3Q
1JuORhI9roBZEeBIw5o876y4LsQd7sa/0Hu3MZzgKrZUsiNakC9Vg0IAEaKxoeMh
Cw6titjEkDfJzkiQZDzPpGoUtJg4VHJA1NBcu7tdX4/TRgnpuIEb8mnNlELAlChG
88kupCrOvmlgt/NYmzBTLrKMMPXQkfR7PciUjWrZNURbs8Pnb7a/bjtTz0CKkUW2
yBEgAQp22wb+BViC75t2Gc+zsn7b8KkwUjCHWJrweUuujZumSNvRXCsn5BCBVT2p
VysSpM1Rs0/3iQbY9NQvdquvA6IpIcr+bv91vKka7tLShQisCGBih8SqxlQ5z2BG
tpnTSRQhyf4grdgiyWKmhEeo/AP8ut4V/7yIR3Z6xLOrHfzm2Or7/tOT0Gd6oEO+
yDuqNju/EW2Iapw6th8ZdwJHOF/FKCSAdZNJxuHjWH+RHuvg0FKUp+/qvQiMWZgQ
N+NzSThr9KXNTzakeGdecGv0se8Xq6vOGkG9rmxsORK7SVTeO5W4P37ceHBePBVo
OadTAiPK9syMItrOZM45Bz7tfk4FKZnRxQmg2bsjw8v/8vAw2sbPQ75KRYGHTAx8
ExFJ+FQZB9lejrFITE76U6Mr5dYCC1KqytwgSCPaTV5TUPwTLSUpqiWFhNhDTz25
CF5PDlg0y0dz3aqx82H3uTtkiGCgXsGnwAViWsL6jMUSVVXcP0vu+JHg4NkR505t
t2OWiK5/MosejBlRtMV4u8FyGEMP/8DIi8UIwmBgly0Hm+pFbXfnsnoBS3nTVboB
+9XGAdAzNkKRxzer+fBHSk98W4etpFvMvFs2EZ12l/YUhbgnpdltGchPjvhmZrUo
MbZL4nSJoIliefelHAx1N9YWPPGpJ9ZXW5TSrBoo1flW3nB/p8lgVn1k4w1c2XpU
b7kdmibowfnVwNwnEoh94Xfwk7tx79X1ogr/MBZiLqGs4s+RVvQ56Tm/UPIu6ja9
GHPdDiXZkn+Sb7/pgTBFgtYaUqXTIWrI7gyPoyGvYto7EydbijNTTEI3hZEEuUeD
5ovWY/zAMuCPL+FNDk0QF0PAFeLt9s8MVy/iLEafnrkY6vGGWaCDjmb3l+McP/DN
dvx8lgBxwbD6gYTDIdvvN28ohQpA3CDrKj3JUYseDHOoujdaFZ7NNh7GhQaqACLK
hFzn1aQtyP+fl15tMdL2ew6EmHLgkf5/eufetIMHObGm6TDqTKhrXkmeKMI/bL74
znLNfwqe2UJ5H0GzFx5bKOzXBmi6m+mD/e0GozcicmytDTyUuscy+02c/S+KMYOt
tYhFcF0AuoV5RUmnF32LBPLDg7IU7absczhM/t7GnURrBvS/n+Ins0hcWriN3lK1
kjoIwAE1E0MwQTCmWwq9wRho1wnkXoy3J0mlwODctCikWKaM9blKQxlRs2ZIvjPX
pfSsCitt+m1BgPBJMsszxaTjX2ZfK6jG7wm3NmeanDfmoY/2LzNz70fmY1hnsPRt
1dyRQBnPHEH9gZTButCQT9Mi5NkqqNHM89Udf03/1lEQ+cIbQRGlgASGPthuXmd0
nvAjd9OuV4biZzoe1eUy8jrWZgA8jP3tdWBrr9ALtY/eyF4lH/X9YmFFpRCr7LwZ
21sKJtHHoa+0VA4tRUbtBIt14efHCa2RTy4MR5wKht4vZ8Dg26f91KW0EFLXmHnW
DCWAVQq15gJBRONf95NBdax10doBNNvEjcchr5ALYKx+5Q609i7iYZSv3xE+7xZG
TfaSF3mZbSQ4k7kL0Ndr+jjOyNLdAnUJiP17R6WAES5Qy+7ahEkkWbgZ178fgrqS
+0Y8mHqgVjRuCCd1A6OVZxtz46uXJWjZWUG4xKVp/EYpjhvZr1r2DIZ3+xn8rXBu
DCfMxNFCpHXcKtKUJjKxLexOfIXg1opOrC8a+eRPtlIlYPZQUuJa/iX2yTcMhFIZ
r9KYugh0XxirIElVFmlsYVU74wNgK11xntcxW6XWAcMDGqyUNcynnGVSxV5F2oj8
OE42O3OWwIQLcd+xHt9ufLKLMthJ004VxFJ24eaxmnNjehL8/A+v0LraDIXCTQZ9
26NwsCivL+i588/Yf/fjQ+H3NXHOWKQ1XBNdRSquNo3MJPoQtOncCXflP3UjGdPz
C98gOX3qQ74PbxtfQtimdKwDz/Q8nA9SjEHjyB8/MUJ45HZd0YpelhxEmDPtJRLe
EvfF+eKiItjlQeP8bJWrcmUI4cxWTR0TKk74qdE/i5b8JfDcsSTyD17xWAHZe3nc
u6HzhRsTN0AovtzGHAnTVHA8iVk8Pr82+CQoifEDQ7WPdDivJyus+e6u5LiZlbYj
QWXw5pPcPB+m0CsPL7baKE+liO0EBYO7TQYRo/F1QWrGz+qk0P9zOB7mTiXOOe4+
ric/oKAFFiAHKT/EjY/NHw3m03E9okRwmS5ggaJQBiOsbAyCceCV/Lwv07FhPdRC
Ku/nSnQA9c9Qw0SzS6QD9dDajg6sLhqMamshVynWDrhhqA0IanTKf5B5oCoc2E4N
axxJSKksGVALzm5COEV0dE6RNTnp/YutzyZ0kQtI0MhCNSL3l89dCJFf+lCpg+DC
1Uqn5oRDCoC0izMpe3CBBro8rXK1AiUysDTGC2RjXFjyLjgj2+zCy62Z/rJ/lZ7p
SG+RqQ1hXyr12F0pCHJG4Wz74motSRK9ZwtmTj0Gcj7R3zSrEjaNa71DFZrrQytO
K/jJxx4YrU9hG0RZ60SKMZ6C+4mCsqQti5BKPJTwoUWgbI6aJU/XzTBq1t0ETjh4
WSkhds4dpWfPZPGK3y4+4lAijVupdbBdu8bXAYX9tAYJ0slPOflLF++5LNJmd6s/
p7TqPqvqnzZmG06q08R4dGarVFAkaMK2ql4P0WkXAEbGv2pj1zzDnEUPOEBZlcXI
x9MyPjlbduybUWW7R/Lpcema14AcjcnAVlcVC3/tgrxLEv4S0PAg6lId5oWHwGTN
Si39poUmAL7pyxmvrixxa2c+PJJCmDTV7GnS2QmpPkzj4MkMtTyKIWkQIvxfToOH
BcwftwyAClOupWjpK7rIi6oNEeGTn8KzxxNELqtYM9Pd9Om07c1tjqtr2ebXGLxZ
xfaX8G4zOWEuv7aq0PqJoSySZ2blmOdQhRJKUnwgmGePAsJ/JIjGUjBwKHsn3Iil
S6Q1iaraY+BPsX4klFdG6hScqjlNxHsgggmf+OmeK5uANs+KmAVRe2bJBfNXdWhy
VWeLwdPRm4cG45kzLO6IfNqbf2zT2LTdoR5jm1oje6jjGA+8RGpXOWWcLaU2zUFP
l9oaUGFPqAHkjqUPHsw4dzMQmR5jsBmQajkg4oRlxm516xTnsqgXqryk5H2Mn7qL
E0y62vi8KotRU6M+pEvOFz5xv/BO5GQ+ZHkeKpkiKlF1U3YFqz9nxVv+trHq63/v
nPs1u2YkjxnIDE92mnPkRH2ZzN9NBTj/Al4dMTLTBClxAxs4Kv5wuV0fGaz4fuVG
4p+qnev693n5iLBKd8Vqry3oer7w/S4WiXXTm9+9FAlP3/Zn9yY7/9XQ/QIAKQ63
FhnHS0ak3+0jdpcJME85X2nAJAs4F6dkr33zoVG2/w7azS45JYeCuKJsf8ceAdbp
cRwQTQp4ytgQBNPa6CMES2NQsdh2uypisRGOmmdajBnGo5CH9hAD9V3k45bYWVFl
kmEsjlS/znkL4LdlmIP1Q2qzTwblpoC4OnpOgFy2mrObSHWU4LgTI8s1fuukMOHJ
tCjSxDPvbuKBuCLIDo0xKMpwWtHPef5JRzYM4V1Y+PY1yQewyVP5HpSnJdor3GaL
rhvC7j79cWY7KKpIuqmnu5qbL0f9+0sMEllBAXvM9NZC8dmYJBctW1j0H+eTAmne
0CgjcnIF9KiOxx2mZxiNM81Jy1PcPGoaWOMols1TqbvETsw4GrdqR1BIoSHM7lgG
dufwcohVqdmT+VbQMog3p+liosH8f/Lth60gDmJAHwV7fmykxfYHuwEGwS8xRPhR
b4xUCcXrOXd7hQasoWZF65lDl0qu1lN/hgog3Cm5QrJElVKkntB9Dp77pMr9cJG/
UKfQ/PetoTdSM/7dLH3fGl4GSbYvls3FElw4sExEUAlo2rxnFzxL7aQYC1S07Pg/
yr4t8utxI/GdpqTFLN2nCKW0ZTCdg7VIAUiptoroyPYXnU+20TaKTBVMisavqM55
sY3prdc0zjDOJgD9RMZcjrzeFzMK1o8dYdir7+CDog5tLjgsG5VYix9o9ShxhHLg
1EQWkZ+E29hYWFcIht19pR17EdOiKB09BnXCj3EDAvWg4tlB2d1J6jGI4Aidacru
tceG5Zx14Oo+dPVBtKfg0Z25LhIM/PVBZ0h30fOtEEteD8iBfGUbnYGxpgKzsttT
qRw82SDCi5wIwnY84JnxB3tJSO/TJMpKlreKXREwuoP3OwANV0o36jAL+rt9Wiv0
SYqqdAnIGseWVx0fZFWk1xDbNKUnIWjsqesDt5oBXq5/hyw1WQV2Sytu9IA1rFuE
07bMNJuFsBOL0REDA0wgCezUD47Gkq2FbHxj4dOzw/daeFbqTEhiwCnOigayfBjR
msvMjdbI69BsqK/BKf3f25BLplbqfFZOZh8xQCnt+V3PRsuEpDCPEL0SWptjx1Et
aPxp5wNTOF0KlLf4t5oYUyhUFyXWetHVMicFJt7Bgxq1bHtkx3Hm62gf6a/yNPqu
M7wCgL4sxy+rH/pG8U9sARN6+/P687rnxT9s0e682K1qaJNIbFqrCaNVvDEhIVb/
9OdsBLDepbr9w/zgEA4MCRSxrJtInWSBYXT5ITpslATETcvXhSoKBk0rU8EJH+Zx
UsM2Vt6AfX4gUyVAxMa/RAZOfo6jC3wuQvXfZ26KT/mNoG2t2Z+zWzti6HNqzodQ
UD4PgFHV+4XraZH5bZlpm0Mv1ElD4Qn0LhTVjz/QsZxouqX5MppnvjNX3AMWiSFE
xI/dY3PtJG96Pefq9EGBikU4Vp56LDNjeEc4Qree0s9aHx6/38nCIVakmDX37TFT
OH+TC4hZJpL3H4yyrFtdPmAtPpn0S28cKAE1/aSwXnqi6AvBdwC6JQwzCB0gtdKm
HZW4HSKJQlkZZmPgY1OuVv+vyvD+jFCQMz8fhNPikY/tP4UPyjmkzNcdjhO2pvCJ
tz476kDgq5JdNGm1Nkb22ramcEemg9wyMCb2vzTrJWqBTS1YvpsMfEFmLJFTfrbR
gmrRjK9uTkVivAwPP7Bkn6k6lvEoWtVX8hTp3nDsAR5I26Wk5m5ftRich51SPVeM
rjG51jkN1vwk4xJHhTa8pKZs0J6bjkcnM3KRYcEwhvj30wEWSTFcZNWqbdCEAX+t
4gHSQLdGW2YkWHgaDm4avPdY9sUcHlBg2KsxNjCO+z1BWn9/0mgJLEgqWvgInCiG
cbNbOeAZMkFiwb8LtGQslwgcNJ2PpQo4M5ei1eNrsbc0ak94S0UZZd2NJIEOrYot
1gferSgLavaNQcwVJaNAK3+5rglWTvVt7JE3oXSKpViFTcSGUCX7GxI1GkIyXQrM
BhqVOXXk21s4PD8cVscICbHc9uRbFsDDamXVu79WvobJ4zlQifcpCV+LG3QCCbmX
bpovOXjkuK8UGg6j/u28wvrF7L34JTo6wph0EVfi8f10+LLVrNcgu9cJIoqYJhFy
voJ765p8vi92M+vxjFr5/KKbif9TT8U7g7spvEiLq4UtqvlqiGNo0asVfL90mP6t
wQxR1xC1R5F8/p4m1QJGjdXRZmKEujxVAV4kzKfAUy77EjCiGD/qrPEO/3Ckv9OF
9cb5PHTOsVwR12cP5vXsqfqblzgRAnuwsDi3Ha/6iSONm5Ynwz9Y73mrOkfAN42A
OmN89TiIEEhC/B5u4zSRne6r5h29GcHpCzOZiKeWVy1yZ0xpwfi5O7WSFcJEHNrz
y4D4+MYrBjqIIZowk8UaQsERbj566JtgnmZgCmX7tI/VC5znCgYwG0mogks4DzmW
sP3hcJFL7oOx2cuBR7eUHzaSM56tV0PGTSeg68dg4ozX//1olzlwDPiYLwUBBaUt
tkNKOGS19JLZYeqOcJzJzUdNRfTxOBFwOnRWNAXXg3pMdRYDLvOfkTfSixW1XLOT
r8C+KUYCp8MUovxdGiTLouZh6F0hv9ZlG6VX3aaqdsiow/qsN8E6/5c0qnjOeV/I
p84jky/zlN4i8ry/NJEDVFDPZ/4R+Go3IDbEMhhBeDXkYMmdK1N7Fy4DyVUkmf5t
chFo4eVtkitjGURGi59FyqUPFuhDZYMJiP7VgIv0vr0MJesHoicEzJCIXEIx+m/T
rAMEyULapKecIh7oqZia62Zby2hjY4REDfK2w+TyQTog7d/C8cnHFAOT/fhDRLHw
RxTYCl2DfNFz6VXcQXxruN1pXoUrOZr3H+Lsjgl9lC56svMSFZJvz0fwUGR84Wa3
PrK1Tcr9j07IzB8/q8yn8IgpgoA3ouJOrt4hH0U5asp1eiZ1WydS+nNKn6P58nvG
Yuzh7ciel/RLuEC26Oi5gHeTv1nD0cF4u9ly5YDTst/4vO1YUrel3CPQ/+oUVKRW
iTlxs7P08LnEPg+2jqsjUHEVwAmYyHJgQWH+lacgwLx2ZmsSKywFdNpDxAfLP6V4
h0O0qxR79wuVcK+dtzp2PC+Hzez5QZE1E23aJPxaQUgziQ+uEA+0BcJOx9oxs/fJ
XCGFWDsOnw2vnuA1nODBGuhUcx+WF3EB5sVH3xjT4IAQ1wl+Sta/3iAuTk9o0Ce4
Kqst8NF/NrLRqAferii3pRWQpiZd55EWlmWedOd68yuvURLAiUZayEtH4WNTlfuc
811RrN6FaDWNlFLto0r68RL1e+LP5vZEYSdM+WO6poxPzZw15gEtV1fagihMf/x8
7+joKkfjuKJRCC17uCtPiod1z5DzYrP7ulFSqVLJW9hchmlXtH118ebAqmDE1DU0
DoABdTIZBkuQCOHewQLhYKGWb8gY33PEUqQ/DDYsISDvQc9m2QW3hMfLevXN86HI
Zj5HaG1NyZkCbVgLhLCTd9swoNVAxcLJ4bNNlUKCATXyFtdrP4d4Tc5Wgx+s5jhx
FDhueeWac5qiE89I0LDkeYvrmkULPAjxgb38M7WiWynKwAvh1qb/Fn+mk3fkb/Gv
MYRCszkUNtz417MpFIwyuCC4FtfJtGtg+j5ZbGhX7tdXtgj+WzGQvyVKehk2U1X+
v7QXUfkPfDyPnakxaxmyuwxz2JD/MgN8pIUI9TxxCq7ImD4Gn897zW+Q3v+gDCPs
P0SJtdgNINHTme63TQyokYkXe/Ec6rxYuvMJDa9YbzIQyETklIqmC5yjTifNAm23
qovY9HcJx7LrxQfZmpKHbs6wHuqDaJFQ4b/Ym+jUZB4WV2Ht7OhRUYXSdRcwB1uN
hBIUjQX4ndaccGIxJxB9BE4aIy4/ajU4OzrtGCEge5tLkOsPbxG46BihHxgOs8Vv
4Xcyh3XHa0PU15hqwirZ25EQvznU5oh1hsWAqV1uOw6cRuOpeeiukGD7/3ziKAQz
B7aDqM+HZ/Z1mMk6g4WWlV/Tq6gKY+ozWl6DPLSD7rUn5NGiDHfxS9BQOltSxDY0
aCS0mTDblj3zpC3cnntBQ8XKdNEY/bPWyh+DCBnfsjZuOocWb+DzYoo8Pg7Yv1Bv
5NFUYpm2Ok2WWtySUtPSDL8knZi/YKMJBi/LEX+1WlZvoMlnpLlwalBGyKhnmYQ2
0KeFE8t+wh4Jul8cVWR9D88JUs6Oafk70LK0TS6bt7wOhtzxg+832vyE+NXfvgN2
pCIAJdvh9Jy8sPqwVHtO1K/2Cazu3fFo36ZEkSDsHgeLqmITxQ9NRMkRSWBj62E+
ApfzDviMz45FBKij4M5JsH17rUDn2L6352tQnfrSz7Pf2EBCD6JOuANg2edXUEIq
wWK9f048SEtbhtwJNbh583cYaHTy/ZHlOLZlhdbuRe8qiylmMYOBQM5+g2S0xgNo
Z8+/XBXeVs4u4RIhuZmpqdbEcHwv0UPJ7If7gtbJrejtNKIxDYP2CCbBtorg5SNa
TqgnqDpuNqw3gunEA0+ioL14ixQ+Lx6JiSaM0gUgH5WUlp2tXwYmVKi4yHmWK04f
klMXCMnc0aLBtjkQnn7ppwXrU02p0QLcl6t5P3PicxZ9cUYsIzc1TZ3SYCNioi6W
wxpKFWBH9MZeyjSo4KRXTZza4sd2WxSHFboCm9ZaZ+dQ6pwGGDE4Q/ti2DdmLHNW
lXKVPvWjyTbKjNC6mxpNGE0rbMsK078xOxeWqcFq1z/5OLtDQRDSYwgaNMtODSWG
p478qRmBHw4flzpfy7z5w0zn1jML3X+2OJaWU5zqYNE4zFBObg3O6hBozS2DatTt
4fyTIVxNz0vyXk6R4SluezNakqfdxFb0yRua75dk2QuDZFpelJTpsfhDjdJ6hxkQ
D61sLHz6cY06SWG1kIjlt/JC1CyoSXDQlWXYEJnFRWOLb3IIgjVujt0qHPu1S6ty
C0zJUFzISbD2+C7Rk+/IUPFZUnsbbEEegrjfjD4tq0vN09VsTBcSuGAVP8waWgsy
Amwlf20hL/nNLsU08Tgy8wHNC1/1ho05fiRyEfpE5igjqBw8iUP2l+n+SAZ6r69c
XXRrWSsA5ZRA07xDk6dbUFhICcFt2kcNjRuFehN44uPNs427e+Qugp4ELHgxLKJd
7ie7QFKoM9d2M6lZP4TAWBW4RCe48MMXBVwEMwok3r8AIveDQuVIjVxz2Fjf7Yeo
erStMweMvcUow2l1PeeZcYn9lMtX7a0xf1q0SlFT/9E70LLL6lhEZoFl742tgo4+
FiS3ri6avQcQySMSDQIgY6f0aQTxGMma6UDbQRiFbo5pVdK18O7/L0wQjwrXCA/Z
2Lt9r4Y0j92t5kpc51hpe3YdRvf7UBtghK5FmzqCrHEjzeEYKahbQFYu8oCf/NMl
X906KdhpU3vRiJt2mhcmod0dbXt34E7xGP133UzDZgkvaoPN+JR1+gpqxSd2Wzed
VBeQqC+CzoRUP27gStQkP80CFaPlKADpqIE9qa1i47ItU5ZGrLGgma6XSm+pELHb
xt7tPzFQZ5IGlDP+Rd4zhIErxhjyezJ9QmQv2DLGorNlNpCgnH5XC5wouiz5bkTA
IAaGSn/vUd6zqXpkXqQvfPEq19FnIXQF4Lo5DrCsWmbv2UgzmP/1VCFa4vZ9MrZf
4XOXEFg+VqiHKI6Nc0v49W4ZmHnN7iKv4GRc8Cns4NB6Qw9IeewS+M1tJ7nYR74I
zioRdoLmXP787AXe8dBjrvydZ2p/HVPefRn1L83lcVAl7sIEXNT5VsztHpdPktnu
Nsjn43bk5aB3VxumygK9PvEHraqTODXWsbIfLbKTBVOfQQbMW7czaVVQxYScMPH6
7i6IZNll/wdZ2pcmYdGZ+qCPWnpjZ1YuL/JSBbA/PjRyUqj3i/ruPu4eEUV74XkB
8G9Qf8ffEW9N+UPi1ImGPdGu66dd4f0T7mCcql46RldSuYOvbpIKMTax+wyoA9r8
JrXrgeKWxIc2so6Yh//Zxi4cke4kOBeQ6zKMqb4cFRcru6dB5KF2NNcG7njR4FLf
SqA9wp84sF6ZfQlH6io6To8L2VnkybfLMvWgfn8Gmun7hPfzdrPypHDxT7elh+Kx
c6wJwGNwiFz+c8qNhsVqEbqGTdDwg3x6JWa0F4AAzBuu8CtZ0Yzr/d45FEhQd5qE
OOa4Yybc+23e2afpqmK1st3sajPPQ+icvEMxVq1SB1Gyau22JLxky+9q2O54TZ6y
reUQ2xFUGY20/teDTzRdglu2eVM6BuKEsoTuAL1NpWhebSmJR2cBbsDB14YCkX0b
rmjfxxHhXeFpBdOc+5CcsYlTDoebOzLIY54uJjexCIY4goyOJj4oSbxJDfYa7kb+
8w+giMSdMX1xESnY3jl4ke9RtUR/tPj09j4Uo0s4gSYU6r3sFUhGj0632dEX4VIO
MvTov2pJ1qFbMFQXr0mly+NLuLtVLYI9AoCdOK4KnnRrzmYsU1ZmewyhT4Wt3reO
5wFEWQtRFkDngDcDBlYWCm+rAWy24LG95ody1iKY+th5xKQwxW26/fjS0CWKStHW
taw40+q3Skv+M3yQ3reRr1/CwFcvw59GtSg4trDdoApxlqMEa9cVoBTwyN3eAtNY
/plm0D4meXtOXjSkflXlmd000NtaOGycr2DL6a0f9JzTOs6rKLePWsyInsNR5M2f
arWWPSLhm/sv2iGQTWwtyGm8hPrzshHBjj/EX4cmOc1xCO/dlaOGhYr3DJ+zk+FZ
8KPcDgATq0RJe7U03xyngz3cRpzpKIXnZhA2WyDusL29ua9P5iLChu0buxi2XciF
ifw4jXENwqZvrR36cj1mwc82DerjF/hsIhNwj7xUKBaNpFJBkrFmenE80dQleUtq
EoF+VokJSgFJBkVYER3/z+q82V8dKnfam7a7B5DTn+hEtLH53iFeJ05S4RTKUKRI
AHqh1LRCljhsoy+tpJlkIGm+4AN27BgsC9KAdk5ce5xOMM+o5zoDglTidR+nQix1
mAa9VHrqq9BNezIwwe0IRxnh5aJ82rb2m+pw+qtfKvJU9IofGLPniaOOT+BcrDR0
1pdruKXbXPRH3lCJJRb8JaWcReKAGHX+UU8kGFNkVJEe/uEYXkhlodEaOvLrD2ks
fWh5UudF1z/GX+NJu2pQUetI2h8ueRzy9Azy9qsZuObPyHCiMkV4taAhaKH1nxhw
/AYU2fq4zz8/LaRQ9W4Q1kzZAzXShfEZm8YgDfR48W2iwfV0cp0RsT7S5aLgX8yc
UAuBEKHzubYrpcB7ZJG9MsshyJ5MytoD3UhFTKb8GD9vfzTzUyRluMVrm9DdQREc
tTRq0RRzdlkLMjPJ3s/fCa+Jiknes+99gymqc7t/t2Ra7UbwNSvVlj1S2lGDjziC
t+4fPx5lNHZQhqt5N6j0Nmz/02B0orMrP4CAmLWc869xC7OP7Tp99Za8NtDI+2Ql
WF2VGUK4Qc+n4PQ4hFzxTvaQ+CA1XmcFgiWMxe64T5Tnq6g+h7hxej1nWTAkxqGs
IWSBTRYWnv1XPYwSozX1UtVGfSIWQnHkYSp2uEsKSn7NA9hF/oQeATlpe7aPlAq+
RrM0d4MNDdVOz6n4yv3Pg2pX94XpvvYVK1OCq7wtHld+TiAxj46X+MTpe9uxkPsK
j9/T8ZEUoqHBLe61ukGmLqomD3mXts/O8xdx4H1luXfau0wa/qJGQsXW0jY8ogMr
Xj+Rm0OiEsRLUYi/1vRTOEZ6VLyPX1QsyMptfsE+iGpjiH8Z6a6tRtWQ9lHA/2Zz
bSTwiOJpWu/sEeLU5TruPBg4I/Q4QyHk3Ug70blCB1Fjx23IpDU+MxfpG8Dxb+H8
yXesCEoL2JQCa51FJMAb1qGHkloL1Q/kodCcANDHKu5hvlqZTCnwTandW1cmkH0W
kQw1TV5aANGa4Z7n1vnZObEs6gLL9rN82s6ImQe9mtdcYBFYE4EYNvHpKSdRiQ10
SJa79/RlMepaBcvhThjBa6zJeCg+BRCVidihIF5i8zk+0pNVloAAGj0gCfkv0PG0
ht8rnitRm9n3JQMayibB8Eh5YmRbkzo5pZM/QyVhBhXQ5wGMlr5ibfEhmhZeXbMK
AgHVlTYZs9SFOWKyyl/DqJDsJRFU2q4c1so2o4J4tNe0TXntCIU72BCxSo9Wnmhy
Ap5VHwY0slJ/cll0Z5W69EYIBDivLT4kf7rHe/wJWPULKcWk0+h9c1RE1BY/CCiu
nuoLzmBCyYZt7O6oK97jZZk53ncaCXrD4010cPiCWUyTwTLvyJvh185YB7aBAwEq
4r0lVpZzvjkaQMlebguduVNM2pHe1WFVyWqpPBz1lOVPwRg4knV5n0HgiQtoY0V5
hriAUzuwl/Yv6RqNTA+XKhUPXiaXH+0Coz07n3SM3FO4DxBmhcXJaNJ6fEIvCZNv
NaRHJTsF8aWRcJTIlGiRAKjKqSa8XsKxY/ssvbmj3hJJtnefjSktYsErYEzcbzMH
o9LdWcExeyUMNlaEwgbnWIvf6WrEnh7foQBmIUs0qgxwPgHFVNR6HV6OORwhiQB1
aYEqEW96qbzXcMTocEI/FmE0+yWnpDi+/WrgBK64rIWv8BaaiJ0fNa4KOlPwfGx/
3rQmmeu45hPJA9TXH0Nsd9a4u8MfFJcydoFH+RDZP+iQxmea+ESB7SVTUN8hXEBZ
XaG8iOF/Of6XUEVWMIaXTVPHcysho6uxRo8NUMjF4GA1KzBwZYTAUGHMB12oQONn
NLBKteIoCUqIMqmpV5h49OlwbzvPviYfL3m7AJ2a6Mp23bVd6UTjGFnmjaMV/lZP
ebXoKyzj7r1+E6zS9S+g/26758IYcqpob4VVnv9CUQ6a0EuGE+7KuG9auKXMrvPE
yD/wwfwezOTdSo2V5golR5On7anx7yjHuDdOv0BjDUpKieS+mYhBmdMnMSe/bjuk
qBMJZ1UmJJryRy2Ewp0Z99w7hjtooUe3xb91x1SLAaO958oVTkxlX7OioCTTgrGn
0XwGL4FTwske5tIqpmcTlILakrD0QTb/x0Yx++bnlPBy9V5L4z8dZUmQTex3KpUD
hAL7968y8jte6VEwOzueogGW53jPZbkcsMAHTyfklY/Pv6j7a4Zs/zYuGXuCjxzO
3/CAyAUisNvhnXIr5PTwG884getfqEh8wzkldhScjOdhl/BVgQUH1gLniKo9C5sA
qaBPRFcqS3OUPyFG7E20BbolvKuCgTe14riaeC2VidIEswrAwFxLVBO8oxYYcgWb
NlQuTDSeI20FksHQrUBLSObTHJi2rmpV1tyYEjhVPTDYxJQY52Mq0Cnl6/E7wfkj
My42jL1XKY13dH/YZ9vNQLa9cLn20t/NkfFaOXh6Os4mYhdIwaBiA5WwIXK7cgu4
2Chwsuc9thynuz4SwlbqLCZnZApDvUryZflmnxyGtiQ/grc923sr9TmRF+FvLyHw
Zwu68XDSi/H+Cr50H5axDSV/ReY7MBYcxgCwpOzYz7suxrG60YrwVrO+P6Yvy7ja
ajwlFTzVpQvrlTidDq+bvLomyjW8dMiitR1VHtqku8egUKjhPRoZ7T6iFd49GsH4
PE6PkpGhErxTGtyiVqLU/v3dVT7O7xSt4pv4nrAXxbG6pO5anjLuOoEL0hM3aTV9
suqVXQ18mkZIH4nlECC5yfT2qImWSWRgo2vBYgg7IFWmLW5CY/G+/wYd7n0Bo4ZB
JcpF3Yj177jpIADPx981ABPYzeHsx0333tmFkS2Dm1S452QpBdME0xkxqYv9b1R3
AV2xL054qAbP55o1bdMMAfNIURK03WltU1dkafnayO7Zo+t16qSkjxuNbouigmI4
8VDOyMJZDiFgA2JPbcJuU5sd/sv1R+c5nIXnyLav6y2ol0KlGo6jV89WVwducjiJ
kQf/AlzryfWD3LwfZvQ4LXd8t5iD9xbpbHAuSkoFUWtUuhLv1DmaFkSKdpnOfNXg
NPMORPTtLZz+9H3g04eobyTV35p0Md3Iedfpmbw8HMBP57Y+/ODtxt6yAKlkcSgy
qoyjcyGUop8EikqCWlM48aoNeMCOYan45kv1cGghYpxSmhJw5bKDDkg2cLlQffnT
yVob3VX/LI+lrxYeOefW0EreQtZ8BQJGW+bU9pQYWgDqbeITNcq5XAlbU5GOOPtD
a/ya/hNRkCYb0dqpDZjqOtct4CRUrRaPHZdYf+fnW/Zd4fjM+FFDeZ7gc6OYvJ68
Thcyusqe6uOQTUCBMw9kIxmpShlp7LgDCdeAKl6QQ9/bVh8l6Wu0JOSpYXPDvR+0
8egMazi43VDv7WpzkHb+d7WMBMPGpCekiH6NXlMdMD5Z29b3/sbhLW0VDCrfcR99
lrLiuluAPemuSRoGhlV2ldqt1I87ecTFZ5Y9mOsxA8p0uyBsffyUcZ/8HNXH0rtE
78z5gRT8Sq23GdFB4ujxg4K25XN5b8WsBwuxvkORtzvbkM+eRPOJ70e//Kb6zkMA
2p1VCqxL2EWugPNAYEfQsP5+f5A6FVYlSxvpKsWYx+SKuF43Pp3Nl0+HBhPt7ha9
q3njFM7zv2UTi7Xa0Qy0TUARKLwo1R3Otn5PPn0+gX0Zpnt5H9I343WiG44OQN9P
D7rpTdhCiTtNwjNzVfHoyQMKM4fComnk1V+aMN0YAsIickXoqCqMF9hkh7cnEVMC
XURw70qXptPd1igj2mx2pPGPjfHFNThDc6xx/5HT5RpBKv1zMVaVZbX3CNjvCqOI
FPmQT6LDhGqwouFz3oB7xUXgJz3ee723q9Pb4JKDZqbEFm5g5pu3EIGU5pJuVV3H
SlihMgOOM8Z5JRpfvKy0Mk9Ns+yCtzFhfAR9iQGvZe3yO6GEIE2L9tTOXtwt9aKj
dh5jOo28NmmkWECrY+rknieSbdcR7rNfYFruFdx/Sbg32aotfJiJ97FQIUWB3KfX
WfkCQ1sverb0Jq4nijlqPAhIZTy7bp95z5cbKj6iAEPYPVm2iwsMMDfMAB21dA7g
H82lUwWxkQC9zb+W5SklfMsRZ4/B92FAxJUVzOEIBNhjkU7O54EIEENHAkd7NDDM
lPLhbZgnr9+8GPY6lnkXQAzTR9OtpQw1evrR/1DR0s5rYh6gotsFXBor3D5qc67q
F3I+D1IAqkoLbcGTSNeCOSfYNKfSBKB4+BBOr4pkeEniOdQsUwcsaYOjTQoIH4oD
YvXdczl0EoFixkERDhwmKP9/DSqFF+tX16jbK7eXLV6LlWwY8sPFmpRbUbBhpxy5
px6whbvwKi+paSplDcQNzBSoGat0d3YGCBfVC8ASLblyEtDXY4kNMQbPfpmFUyRU
Pqka1xqq3TsOkRQ49rl7r3rUqUV9Vn11W+nRJWqp9lRXw7kO8xFPXGEQxz+tEZwV
0WWcI2hcbR3Oa0Lf4wil+bkishuCX85oqRuAFyCOxwLfDz4Alj30yXw19+FO5NyO
ZMAeZ79FawDcOrEA5rBwL/ZrK0oB39nY+qz5oa3UPjs1dhegpKsvwHtnnGjvkuZw
5B5U1CctYGMAT2T03BRsA0n8vix0Lxe7sjFfZ9BdRVRhKzl4KUP35IWp9aq1tgwe
Poe/VeCzOEyOCFtzd51zly5xwBgbzE3jov407oGU3pPudw4tmdvQdzwV0nupnEWI
ZqU1X9qhIcYdFT8O8iXRjunpJJ8Q0f+F0ClyvUhGms/F6znto+UkUzBSK8IXWZKC
gmJNZXeLq/RvBacRjuvjGo1cmlU8CqoltEIpUWWAO28xZ0amNikdtOLJqE5AeSlT
1PA++QYEN+xKPXEvJdxE0O97A0MfXdQU2ylTo6VMDeDANmKYhzcdcuERXVd45QA/
62UOO/8oUFxzkc3mcDybKZHZ1uqYXDJ07nMkzpOkIYFdrmlJpRQWjjANRCXO+fgk
HNGmrm9nyO/DkMSHinNj61Zisu1DH56z2dmKzcsjuG1o2UmUTaGcnF1+B/9p16Ep
nwBPiVvoCQPg2P3fA4XLX98rT34f6uZDlqJyQWS7zNC+5TuGukBw5WTZlX+nI7T2
6TLfJ3fXTolGQsKApJ42kYtE1eaRhVDquKKyPTxTZ3/DdJiFatS8EUb0Jd9pLeoy
lEqG1zFvAS5wtPQUzyQRuyqNf/d0/B31+WdWoYjgkLp7xhhGzESDizPZ1fz+9cgL
jvAn0FM2jtCbYHDP4SUbf12k42zety415SLkqXlnmsoRYcajvRTr0trWt0xtcbX/
Q2bQO6hyqKxJDNBDWLNh2RmLT6N8EqubKQ+ji/6YS3oRq2cruhL7+ATHKIAsR9ye
ekJah5/wExqCxBZbSwwnj2BoCFuL0ZXjODWIhn5IvEdFRJEHdQ+LvGmignlwpUf7
Tt0M6QpkRTzSHxkliSbaVlBIKaMQpCIefT3kHT2UG69LPrNam/FTaOCnCtHb+KUH
mrk1W6a9hzTfWu05ydDeO7AvmpNz4PVU/OW206uDPgXWWZFT9vSj6EXKeliB9K1Q
JhCnICPMNX5BJGdYTm0Kl0ubWesX/qnf9iOdv9wedy3e1qobpocvSUBIoaKm+MsV
EtV+LysYI24FqS0hAPaD4V8itFAxQTiqcsMVnMB7KvE02HXfhWgnD0atbtvzhoq1
bnIOiGpj/yn2BGhMj5opwEV1ligmvOd3I51ybbbsJLqezfJYMYCNgNmOmNzKsVYA
gBzbHZTud8eOfQ/wpJ0WCpp39jOU7hsKuKQbT4VIjXkN1YVGnX1X74oblLr/MNHQ
yWrb/1Z8vqEfU/+c87NJBb46DBP8H3GpOC/SHwlwo/k4Y9Gv+dkDmgQSuNYOenuF
OGYIZ5AaWGmaPL+oWy0yt/91LpBLMfPaRR1JQYDIb10N40vOlvTMjW1pGNmXa3B1
+R9ch1OLuLd2+yEjS40aTq30z+55cb2zEuPIJQ0vcCT7yy6RLQcPB1+1MSzkHEaX
5GAZKwRsadaPaTVp7mVOa0ioUvODEg0tItYl8kQXvarmGPPVCa3wXWMUwqBwWIDX
d4WNo+FGAASlxKT3QzN/YtWOCRyIOyYR8Woph5/Y6ToSMWEOcajrWSx6xPpMvGfS
lfqoUNZMwiYB25oGnxuMYdnqnL+hkM8fd7Mr1o/h6Ma5GRrsqVSRHElapyF7v/xk
Mi/icifCsLXWT7ah/RUJrSq7Yiayeie4bkwwz87ZZ3Q6YJy8XO7a/w/ICtxZl7k/
VLyRHBlt6mcEqMO0lnOHrNIVJGy2G/W4uire84lHRF6tmz85dYls1nsJhi7XjFxb
HUryyCPrcWJRWu94UrzyMsGdE1u2zcYg72XBBvO3Dqc2x1dmi51Mv+DfIf6Y3ZXX
GDMDodC0fz8ZDoXq12LtxiqFCCLecoEX5B3xT+Qbct7Llq0Mf/2L5ahzFhFknDEZ
MFvwjRl86UXBc4oE5PalwuMvxbhYs+2RaDl01knOMWSpY659yDRSSXj7C+RWlOKC
csEfP4dbf/LuZqbLx+JMjErey6WUry4MkTG9WR6jsmn1kdyhAQdgXepe2mGxJlAA
O6uH1CZJOXGwo4ntOi0VMcn3vsUwcZ4D/c6WPGl4ez8Nkak0A2OVtlBYP/TKJSmL
Y6gBPch/D2y53tMeXGiACfw71piKAB+JvDIMuYt/F5HQtqoVTjRL1BOeEC9iF1BS
8IyWddzmu0rqwM3caWAnHvHiN7TLb/AFqtrr6awkYbR3RosiusJ3JU8MNcV8IzlF
COW/QEHH39/3MEO/nmMhcZFrEwdkipbRfE7lAkMOZJ0sbrD2dc/w7oSdFFnIlOED
1ZTZScxkStsgEBjxIzFpeY4gPHG1ifXS69hRR7bREFv24bQnqKdg1WI1k5pOLNJY
43T/p+aTwqayDSMH3c7snpnSCoFGqR17oUBkVUMBHLyHVMUekh2UpkZKFicO2xMy
H29tCmLvRXBlNk8W/7pnfEQY4Rp0HOllROQVOg8vBh/+17vrOILESrWO0Zzs5iPS
lillecYn5yMLsu4bDQ1f3k+/thRETmErSrEhzeYQpHn8uEx8X6mY3OKubbKjDsYH
XDLRrg/ZPGTPqm8+KtqH56Z55KHlvn1Fld7O9fK2q1vXYPLywcSO202QdJXXQFjY
ih+C9xZRAY1FMyl0qlccxErr2gE/c5NHIH8AG1Hfd5NNyknm8PRs3nN+BeSGOHCT
zCtnFo+zpEwl5Ye5cwRASF1eTCIU0vV5XUZ9BVavVviXqeY9NWkjNNMPNjSN0isY
w9f8XTn3nrOU29DTnpERgaAQqaq9X4SmhXJeGZjeDuy7OeoLx8bpLQiLjvVRg+mU
u/H/vuZr9SvrWPGu+oCS2tihh+VYg4RaI6E3FK2u1UMdH2lscGQ8QvUu644jOyWG
+MrHTmZqs1RQ6huj91Z7W37So4BWMBsDWgmkswOoUMqel9q0cTbb6pLFBcZ0tyIs
aVcPWvr8dkhr67ie0jV+IJLr9S1gnz0zjP9RuOBoNh8Dy5maowIOjTHay/gsrp/F
OdmAG+MzHEV0Q9dZ5CsrvUp22J/EgrJ96aaapOTILWKQ7aoZDs93mG7w7r/sT+dv
k7TFDEji8rq7q1QmqeXsso/Bxvmo41TU2YFnrdhd9/ilgrohlfXSxhsFC1E4oVny
YJ2/Emis565eSyk4NKS+GF52qafz9uzLzyc3TmVOohBgzdnkRV0jP2BOz+XnV4CY
Xbga2g9JytxvPEUi827u5JOlZvS6Xljt6d188jUvOhsfKxe7zz27Eu6AUPGsvMYZ
QdDb/3gffwB3J0AuxkP5fuFBwhLKKf22vwGWof8pUJHN3Xeo+Rn9lirp/Se/hx66
WvZeZkQtQSCRMijtE4LSGXu/I7kxo2GnG+Q3KhltxV1pZFn6BseTZA4F9L413RdX
eopc0g+asWR4OFhyXexfZAP3Jd6aqASOk/PNiqexHcuKJeN5GHaGaH9ehDErOWJL
vIEEui8oSUvP0aEQAi3RZguvuPCLilE8OByq7pJyASrcEHpnhadjiP1KBVodyRzO
m91EJd/Gg5JNC/jKgl4nbYuiMe6C5UpYs/UN1pmg1MTjakvOY6hloeTJ1Cwsj043
IkajyXCMs2YpdHkGE7x/SoB0otPSbAa/9nESqRy1GaHMINVU2+71XcLOd7+SWF4h
bNcdPnPJQzXgVEOJXEsgUYUefyT+S0Pv4+Fjr2kjY5LNf3HVdBtdBEDzVX+HpsqV
w0UPUd/NHOtY4ILmxSirKnz+iWCQbLrL9xYjdIGuGezzYsqfpB1d+jhD1IuuaIij
SNkA+ok+cBMYRirgOi2YTgMpHy9zhha0mv5gTp5ZyFqe4jfrZxE24srtiuXoHX2a
A8I8/vqn57IHHMeHaIhkU54HkNjVjyd7ot20sWigWAjBmFmnaRwhzKutYJS7uoGk
u4sTueL+7lvHuH9fegF9zTRN2fTtVCHcl2QqejhQzYZs9llhj2X3F9fbK7BNbM4R
pQ7k6z3DXVhSE5P7FOY55Pv23lrUpkRh+ITnoOBXmM/f8qnBKDHTlzLX2iXdxRNX
aydaQxYRvP7dO9T/k2gK4p+oGhC/zr0g9HE5134XKmOfE/2ubawdEoXPI3n5aDPm
verqT3kSkSjqCWUY8HDqSVKGUbBYagg9iBA63v4ty2lTBE5MAApXr2+Aqh29kzSY
5Y95fXy6907Yvawkunx5ZIsV5X7yPWuF6FA2SrkppThe4TKRIK50H8MuXr8U1VJK
Q8JErM/ktgD9dMkqe1iR6nWrW3/0z+p/Kr5Yz/UVKLpSL+yR0aCK9KG+mmt60eF5
nD7d50kzZkH7mrBvREVc+iHS/2mniy3ViGr1PR8caYIxgXaWQqb4opCEK7+OeBe4
Z2f9PSXwNZu4CVrRFA0V0KVWyNT5wFlVZakjjgDYYqKUHAkhswW5nXIAYVq9LcQn
ANRiV/NdJ8Ea89PNcJBGlHCtwIUWTk6hV/mFlaEmPaTIr4J14buR9uR+TQdlInMq
3emuiql749a50cjfghFVoiEc6G6b1jEN0IfCbl/svM+8ckeNhIPm+CNWivs9jPix
q/B3JTp9YKPqZTeICPc0K5jIHqhAVJUPKCRXQnwIau/k+Ohigb1mNNRcNVmpjdGM
WkyoDenZ4CCHYnoZRohrEVg1bODECLp+ZPjP3RnHs3pb64kEEgbhEYP0t18CvRg6
/a3AtB6qDRqd3ksZHYuTj3RBwb2piVfQjbraiMYeTBSbhQTgZWatlUUW7IudlHhX
EWVg4y4GqX5PbQ9ZS4cTvmpDcrSzp4dStWQPbVWKv8yHICCUkNSRS5/Ux4E0Xbtd
WYNpySLEIp5If508igAyEHKu3k9g2+w+QPLi7TU56vOp7AObTi5BEas4+xXlSPlE
SB5B1wRXSBAJ6nLrmrdAORoCCFks5C/nnxESzqSqNya01VPwNwz2Bp70s8FBS5f7
hZvEHSNrVvmhU8OgUIijtEF4HtA1LxIAdXvM4txQEv+MeHJBl3wnettG4TcV83Br
4RBBPmHMzGMd8Xre+CbWvGPFsgglfQg0k0I7GI2MPBlNduGN4mzPlRv/gYhSznVy
Pg09XUTgCCqmyo6iBTf6/7zdZJCgwga236TDf4q8bg/2aLINWlSX9a9reAkYWYIO
YlX9jOkJzLTibEFhCzrHAoYwtbxuNbikrdUX/RtLcnwmp9o9I352TjMSWZhClHAT
0SwOS0jesXaKgL5SLX4UJThMGS+epywreb3G40sgL2pS0j8n0GGPDurToj3p1A7e
Eg5UrhFf5uNDqNNoO49WoXFuqadZuhOVhr+HYVxiLrTuQe8hB1H7W7litcPIw8af
DQXTqu8Xsl3r/8jnor/Xxvk+K0jZthbFrmmwYepF0J7pdnC0TLzwCvr9tH3vGo5V
7B89VlgcPt1utrljJJ06h//ThTMxUnGV7nCOj9dAh5X5yPvqJwXdFXxUCXtwNNJn
VK6EPt5TzcrJQL7q7pLy/IGK6SoDF5Xc/17hB9udgLI2AMBY3+cPumVKAFERGY74
LdTJXfSBY+jsVYvE4w1czuD2g37fU3Oa7ACF6hIoHZhyhgdRcoQlUkBkeWqxUCBq
b4gqkXbqwKC1UlP2ifVaDiaGXhqaGt1JXjGkyrOupD8R6isd7ml2ynK4HjywdfaC
d7JRuTI3wZzZ7AX3780taTF4fJWxw14TtRDPDsi97XDUjxyXnBzFG3nBpjaB2ect
NakfmmnhijXv+bVQYeASYuLKGIayLiSctNwZuKZE8aa92lMBXBV6e1YR2kNOWcin
sucs67p8cCYkNsFyoxUpuPU0G6Ej4+8rw6ERCenffVatJxJmHIFCLUjsPp1ximLE
ZfYcSRjocm1+lXXt6aJXK3wHn0+uFptOEtIVMRjnf63hDyNU/RutxWgU/I0JP906
tTSXskKku/zqmX3PQplBH/dPfxnz22JXuFFgSGuW0jsHwjZzkKchW7EgihdjPBUM
TwNSwoKTC3N5jl8RJSzL9NKv57c2lioJbJ3ONOeHN/uwo4nV2fTecWxVDbls0hMI
tZM3leceK0AORNiOzAv+WxizAV/jk2a4U98pal00uOxsLjAAxHdbEPQmlkQ8UIh/
+RVUJt8PCIIb4lyjdnutOLGj1N1xfpdwQ5ZzUhKlA+EcDLiKfb1I7BcDiSm+AjcS
eYPc5354xkrndAXWModyluzYxKxbwwXUNTalYBlOzhBpzGinJAKbFXYNK/XIizD8
MAsmYBM7Hq9/jJjNXspv/ft5+5+j7/73d805IDzYV6voj3YcvLhvXCsaLcRtcmFX
MJgJ/CPqc11jwbm+4dG0qisWu98iPigB6eEt/AZxddPyLVl/jJ803j+iQQyZR5h3
67+ptlDp/hFkr6UzQYhFT4lF/i+oUkcNZwt/D3IMAtbTnuo2rMK0NpNo+581Ky4Y
Enrt+N1jdcWVj/UGvyOzqzw1WsO2Ijybga9OtNl8lfqjmraZf5qRtvzeOm+qdX28
5k11IW3PC8QL2+Xlgf42yHIfFnP6R1uQf5gZPhMLMile1uGlxnc93ZjsoXTzVILE
uyUYGoIxfd8UBb1HUJQ+AthAxrCkIWIgOYOlHl7MDkIcYLqClMh4ntI+L6kKpt7k
JNxx/QNjbjG3Ow8jN9qji4xGZSlP/BwVoUt7B9qAW8JovVHVbZoCx7IKqyNPbRB1
DE31vvsbPkcyaegMSKviwAHDofxW2TgbooggIfyen8ayzikRfTEN/3Xwmi6jDx1v
aqp4JjRHbjOe+SP09MbDuZCtXQDv6LHq6GDC/ttjZVGuq6KgFsjbEnq3Gqd3jrtW
dsfm9Qc43IFFap+A9HNIIDZ0pGIxK9Jn3i1pN4arSzy6S/fIpSRso5SJrrKOOQv4
q8UaEAIYAcQqcy9khuHOhe4l4DhjuQwiQJWfETQA0VxIS5u91xIudrZk0r1Jh1pe
0YonclRMfflRN3wEbHSu/JfV9ddNY6iNy9S6UxUQAet6ZMjexNe4Ou5ecOJn5i/r
nunJzDg4C5TTuehJNvf69fieqKTvoZZTj+mMRp6VnG6KSJdm6mszoanmsjvuIx8k
LN3gklURBcwBcFfLnPd+ZatuByNRDKLXGIp0m2NVYRWAHjnuIHMpiIBsTjsPvapf
RWxaASADOfuPUqyt/PaWjHW1dKPteTDZOKQpwc93b5F8++9mos0Wki63cFCv0JEn
e5cuf7GUbsuRfMVvTYJP+/EnDSx8d2ElgCv4o3u3hEHK11vyTpi18Kz6Iuu4diPt
pZLtaTBZyytIUyt2dYMq5kDImXNmaIs57Y2WJtWAyxRov8agtM/rbt89Lh+jfZ3f
MXV9D9Ez99476tFDzpGy7s8EpE6ooprW8iuMcmPX+MsCp5RrDbxkcgMYzX/JBSUC
zHLZZwxCeTz2rji9rrc+2LLNsUr/3DN9pdd1h4vkLXgyaIiuRx4XKPiURmbNclVP
qzd7Yat0NTx2Cm1rOnx5aEUP9Eavl8/QWpGS38z8ijmWps1EI7UMUlX6/A3HznTm
G/lL5bJqCa9sFC89QNxTnPZACaD45cl4VguNpO5gSWyQKw884WMTl4hN53+ASzwT
lrZeVG44EZGBBKupUvm++In61k/L85IBihIMKtomkFiZHvv/qOPGkIS8SxOWKoLU
JbyM41agb/ZP6C6b2AOS02LF/9WsZiJ7tJJCMlYzTi+buk7yWdOWVNyDnf09KqEr
i6mxcLRuSpPGs8u5vY4SngZF873S3QWwkgc+Zq3tabL5uWhCCjdHvgOGjQ6LIc6J
hPh0QnfpRsXWHvxoSP7XKQcp3sI7LPZ2Nh/wsXFZ8FGJ7tuHsW0hPzIZmHZr9oW+
OJa/0Z4nIWJRdHvYMcU8pv6IKuPbNqa824+uLDlltOJoslh9WGWI28iHAoxnK5LX
HKxEEM5pXddp0R3WreE7G02U1DrEfOgQMItIuL5i40fTlvM5ECWPSwGKlnihzWqt
N9nqfx0x66mKCEx581R11RliSOydnbuf883fh9NDlXdFwa63Io7Z+wYO0BJZXabH
fq54z5YNibSspLe/Vi5fS6y1T2AssDif38jZAkSQF5QrBU3BufLLVitBXztmM4pS
O/j7y5aEB7z9HXL2dohcHcWv8zX4DAxh5bIUVuebSLv+3PUDAbIQmIGLvJTJsu0L
WOjRGNCqsBfaaYRNMSk67dp1hdQr9dLwhls8j+5EPl5D0O9WKQGxdcXzVExGTfcU
REt/jRYiJxgQzeTo+LtKdbSvpaiYiRzGs4L0m9JJPRMnYyg3X4Tso8mYD2v7VyUJ
CbheYXDYWLpuDn/GUc3qVH18B2UwJaBUyWXEk5+PKqOWydWXVNoHxpAjC2Qfzy/L
bdxKv5HZePbPvpMIsdz16C6bLw1BmVR6hOxx+r+IzG/IRucHUwZAmkcmgrlxwiEA
n//2YbF6o6xPIHK0+5XH/NSvJ52W8Jqgl7Q1fZEEwKJpctQH9oYhCgceeT46fDDP
P9Rs7hMCj07P1BlFgtdihdwrQ4byNOILU1Lk2INZ2P74gYkeg2DGwi5Nf6SgDPqg
0M6hl+t9O+jS6AKyWj5XOmY9nkvQTyN3X0gkrIbZAPOBoZW5vLpgfPLs7gdlMTDq
FBuF4pIW8vX/90JRo2lIsbg8YoQIGmBHHFyyKcQNc11/S0zs44scA1Lvn2GBt287
o+N8PUA36SlziOST/C6TV1iWQeTEQDI/VQ5KMbKUOkAJck91i35YsB4i2mY9eDp9
2qp605WyKa9LAhxJVWUiofoOq3lrLCdcww/N35zRdKvRfC2pFZKoI44y4qgS9MEG
sX5HHGFXU3gGxIwVYoIZqqz5yGZwbAAGxMLcFaWBEGKxpzzvJ/u4WckXup5pJ2dN
t7NHN4vqwO8Pr4n6y9erqCK+1dX0nsZ1ouvAaIurlv8SVmKeetf7byqxP6Z3BBSr
ldbsIVOYpS9UoD5lmHopgO8YdHZDiBX2SvEPeFiAc94B2eYIq/xYLWbfRytktc4V
U+qmB1QQ8eNWDkHDX0g5+1+fLQSQjWF15lVbCI9cSvzVCSGxskpaNkrkjo5iS4ng
qqISlAEgR4Q4yVxO3ct2BYPslbVvTrNWUj1bNYqstdnTNO444x29yMHqxdJu0zlZ
aihT4THmLB/zSAJuFM7FD4n9c3DfOfeUbWMcfnEWjlx9zVkgSOQlEdf7ZB7OfNhH
YtHyR9T5iKgzD6xZqUuw8g6+YXDEub1YM3EfdOuX5fIGveDVvyK3r92afN0pXJSS
KxEa1LN/ouo434uFweB5u7d1rnYfsdWcxtHd9luKnYOTbprgraal0J3A1m7l++aR
L2iR852gwIULk0hH8cftSJFuyuXAvKzpXqai9A49LFL+b2/1Rubl7os7BiwvAK3h
9K+TSUwB6/9NDreq2dCLNhNt2XVADi3s+5qKDK1uht4YqmKxYqHfB5bhIYlqMNpV
4EBZ1quX770+juUQCrAjJQ9eWp7SJI8YEbTQkapxU4vLVJILtcAu7m5uTfB6Eydw
xnA01xO6S12liX7RMY1IU2eirMwzeD16h+MFMPhT0z2aggNwiQgmoVs6zWUELsWD
kS51Vy0Jx7RWYR5fJxtkaXOQih084UeCOEIaLr41h+a9jxkRzsTzPPLXf2CQp0yA
5Ox98JbYw8TLhRMngDdQXT3DcMbF3ozapzUXFfpMb1yrkHKHjZwldfxxKnnYq0Gq
d5RGTTMVjGSF83UO6OddiPT0FCspDI3x642TqeD54YdTXjJupoKGlifH+I7ctFSH
JoERFECTliYiA5VkG/nV3/m/OP63VQAsVpYQswdh7uywwZKTxpUtJWAQPoRIsEfs
TQP2bziDmF8IPJivEID9kxOYJkMkLgPIxrnc2p08JBOHupUI7jv8rYzGXI2vfvxz
a+1NN+Fp4rWnDPD3Nry6br3wMvhbhQyjhaQjjambE9omdPrLNhxH5C8XVspuCiP3
/TieyNOdZ8KXmtJTTacjKvZpDSUGPdR9kuPkygLfnA3xIvogJC6BUuWclwWq7hOL
cRTE5rRDeyWiZKxrjxjGnb77gGbOL6bDVUn5Kb/VODde+YQ10BQnLkRO3+oZipiz
ntoVYg3HZBhWLT3D5WiZKHh1zirEK16VZrc5bxcMPEaBiPBWH8s3QCUYKKL4aXF9
RKedArMQmegmsZlmpxpZGP0o7ezM7NvE72oJUf5+xnDuV32H7VRD2LHYFGygXkrj
jsYzFbntdKZsULUCBoexq1IpB1Ua3iS8cqrVXZDtZ4AuDjUpYQ7lfWLIbgfOHnQJ
wT7QSCa7t837gbfmYz2qDhGJjIw6Wvh6oTUeznJc4SaTzbsvfJBHA35YHGYx5jaV
fwPGRQrEU6A+GbEkNROd+5HAOU9dFdtmcy8E2Jdr3DAZG+bYidlCClaRNvt0w6oz
mXIBMt/c/zcChB6melwjrNVFvrK9Hp5MZRexrofjtVuRP76TfFQDj/8bmupR6Oem
itWNRbygQtZBVeG2cMniovf1vHN1yM6sr4m2G7vyLTys1Ag3/aZNyAVRUXLM5pCV
VCf0TwNmdEay77OKQn39qXA98iwyIIg4R/XJqgfU2SW1oi9YVBP9WJ53fGtIIkKO
xjp3r7ucfwLeQilmrnAN8CxL03yhI0jVx+Yu72yS4nPPAnSXSm8Dlk7sucfS52oT
/mnDJ6y3sfD5tUYU2zLKwawj8bG8AW9iDZBvL2d27d0N4D5wwWTU1jR66ImwbspK
f1QHq8LNUz96CABPV0ZgQrHVsNbPxU1iaSg2/iHUZq84djp8QuQDujmIsesQs/uH
bj7+AJHRFVZyjMv5MpAHjqIhtr1BmDDaw4ZlH6Fyf9NWCHusuSKOGbG+3Ff7i6Nx
WzG7DVYQuP7jttRlREJGDBoWh8L6S+1ieRwDYv7+sVNk5VMEsghg3A6cRgGC6LHb
cSrwnbOw3sllhpa8MYadLgqy0W2d/rps772WkR3gayDTNUXlRevdRJ3rn7Hrj+p5
Cbsx+VW+ipyUBXSh5IAIzduMrgafMMsib5IMDAete1L2KJpjyuyc5QclXeLSFOd3
ey75g5JLkqmsoALHEKDOyQgLUCmS1X9iBi2GGx7deJrpZ2yZoS3HRPFN3lZCHyxy
mjnez0YIHvPPoxi6ejR4AP59SWClbIVgH/2lpeP3rJaQHcGaUbRMypa7CFkgejnG
axlmC3SL6qKBG4LdKPZ1axeW2+sEJLRH+jwJxTcaaQXoT8DxkQ++BFD+GyDHaQiY
TjDE2gWTkWxPEr2VGy/jGSKCRSBdmyZogoKRd7rJ03OxLHqCdfGYW7/8bIvCsOrC
nEvVfvxobkqErQ7JYlfxEr+E5Np7aaNN1Yjp+mDjS/Sewo5Mb1R5mhcsZwpq+gbw
t+anFPpPTe+La29EVw6oxaixMERHK/c4rkgIJx1e7wTrRpZnZWclY2xFQ0gmhE5H
zG1MiwZMOM+F5Rh822Xpbw7kBny//eUvB20Lg2LzN/8cyoPPgJAQd+6ew/kaHlkl
IeYkl3M4jctt9q0s6yiBeaooh76eTt4kngAgZojc7Qisb8syEIdete+eu8zJLBH/
Rl1PfKazrFU3U/7Gykz6rtAjVY7/pM/D7fsh3p/Ibm/81Np1DjJ3fKUSc6T6eAgH
oslEz8IWRCgCOgKkY2VvAeAXvMfIgkI+xuORpOgcNW1a5eRoYFtXBZ3WYOgMROxD
f8vDMjDBqz+gZIfo/C6jwM8ZhH0vc/D5wAuMVcr3xkmJyZkIvUsJEiBu2mah79hD
9c3RoflsyBaRGiyPzvcjX6vQsw8HTMG4LyNiyIQYrJpoOk+PiY/KFDWZIGr654r/
qvjrlppbjeDqKf68cMiCVGfAfqt2EpzlECn1+jsM1EwF1t1DPMqMoQyyG37Ap4m4
svUhDAM/TTRooDFYpZtIDp6F5YS1OA2TAYcyyqfiL7y2FEXP70s4+0pyUGaweG2W
9JEaS6oECG13pm+YpbiEntqtfhdw5z7tBKe3fHp3fLGLeNOBiR2trIc03iSXcbQG
buHvfqTzwFTR5upSKsvHFhjvWsSIHVSioUG0/dxCpUnkeEDlaAbiqluqVnmnz7AL
59G+QEPsDpAQQPqPhbWBHqvWZTUARc/GrzShwMoZuJbb270406hGudfPOMiiQFY7
f7J3flh+88h5Ks/nzXfdLYOQ1KrO3ruynmrvejKveHvwzki4S1wU4/WF9rcLVD7t
xuxZtSqsrfTWBrr0GLI9R2eiv+xZkCDG83QOfil7Y8xPkE0psgyXDH1EXaxHmTVl
aC8pUdm8MHDYyiLeU3FNakFp+DWrRu1Us486yFa+RBZG6qCKS6U6dGpLQdsuGUHE
V1FlmpHI5LqUPPsEqaLTzqEMFORgNX+XmgC1K0ybkhoaMAuQf1rXDoSkIY3T24Tq
v5eFgdoScG5sLaIPKGOaIGhkz5vu5oL8mFjwh1KARqvWqSS/HgoYVbhAH3L44eXP
6JB5F9uqclUQ4yvyIll785uMLo05zeu0qx7Lkjn/EENq7s4bsRtc3xO0MXU89buh
pmcuA0J5UyhAnBY1dUxPZBJKC1NCDEh/mB0AJPmIhc1z6j8I/568pASmbMR0yvMs
b3QA4uoO8zZLvpxK69IaXLNn3jiLp2DMamcr3v5hSSqE73KpGlaDN0z/80hdnjkt
g1k+IgzZc82h6XaDvURRfppTsPEJKd6VTUny/qBKTglhJufjpBNqdWDjG7CI/DJ2
G0rWhV4G82VVRXKE0GDgE5xkXj8vGRK8vc7fsqMnu8DvYwpjcslggEoMbxyxtYMP
/a7L/2GyNhaXDnY0qOlcZVYafpDpGisJemxxRjDaFSi7sIWZhuKhQ4k8Ta7pbbsd
6wrUsXqc0LD+9Y19TedUUwouov5hlwmSWH+rUEUDDCN5NzXayeh1y1197X0NIOIm
rn06VWoLggBqAV8HVYR7v31QeSDEfcPOj3w1Ip5HAD6VPCnLL7ZTVsVCnvybdeFs
WkjvHmfLfHEtX6vsjl9kh/eKnBQ/HQo8TUDDo45ng4OpHcX7qkVA/FD/mVnMHCSI
00t4mIyU/zkuR/ilPfVD7oM6Bd3YfxtZjMJquyxYctRh7zFf3r+F/twFFfR0UCpW
7UcXMcm4a/uUkwzupDZzNpMJ9RQM2VRqnEeIqD9mCeJTQzefYllh6aCT23Yfmsil
02h2WrXirgKg0HaPssyDkmiII5R7eYyVAAVyE3yoqY1gfe6uq6mMTnQrJVUIlrVm
wuGF3+CxOm68SHtTjF4ZTO/qaD7raoRWB/Kab6XuemUSheBPcT6pGdhX0KTFRshH
QUPfRJrXUZee1fnyW2iof5b2b/OjlGjZDer6P3Q/H9BAAWpoGCR/ZDVv14kGBbzX
P8jV3HQ1QqKwT82IDAlwoKpU9W9DOn1t90l5/24040J4XF/EYPyObDTLk+p5ooAX
qzyMkws06c5FELzujrGw+xBbsU3egoe9XU1NMlGS1VkuudU4V2rhsRPABScMSxGI
tsxsRwASQB0HsRtZCd9JtX2MoA7eJFmblNpiMFUQZm52EDc9rJtOzGDm0HlDArgk
wSw6BBmx2d2KJUjHwN93i38VV8yZWP7ubjQUsS5dh4D69hQ1WUPT6BV8i1BOdLiF
heojg/A+nmOxV1fHdV/7xX8yZ/6eHDMfNRWjnv4ieEDJf4gEvMbOpFDBWAzRpuCF
uMXlL7jjebXdEritkee3CJh/3pb0O91LInp8kbgF59FPFnwdPHFNtxBbkWmKTh01
P3vogaXr7EmL8baba2AAjlUlyK2ie0d4VBXlKwbtvhD3XnCIkn4T3I/zf8PmnzF4
s/sXcgOGjRRGrwIR7g4xxEacn/Q22zz6dU37jVf2Y13O91ExtSXmPTjQ2wBs22hc
7MMzvDJR/DT59rK7Q6I7bCAAJWoHfk9ZaRUDeSa1CqWJQuF6wtlsVFebb1N98fp+
Sjq5rWFRim1UKIs2mbuPkxSfF68C5hzCpIzIxD1aIuJQILb+jCaY0NFyjl5I0Opi
YtgQnQIYQqzQmt9vS4x0+nybFRWESpC3uWWKbLquS44P0VoWkk3F1AunKigmXpl/
VnfyQ/o88Ci0Fx4WTw5/xFjIPgrS/7EkPx4naoml5bUmt0SDq96RkXm0LCTS8FZ2
sI5m+knBnCXDhX9oRfIlmjUnmmLPXBM9hATN9vqP2eUs+YdS7ZH9nv4LdDqcw2Qn
pgg6BEb9fsdK9SQrTd3fOnb78naFw2XXeOgPrswqWrjIbhiiudoeSVPIqQyGC0rY
fNzCo1RDiztiDLiwOYyEmHIfR+F9/XdsJDbGQ0G914RZhhB4ZAs99NiS0e8rgTmz
VnBwf4jWCVnyXlRdB4yH1kQo4k1J7cR1g1rxQHsxVY0mo7vv8WqvrpJD553Gj4ub
cCBmfSrnK+1VVEv9yUdzRlumOy+ftV3uO7qoG2x4f6lqKnzV9ohvMS9vvAt9EYBP
sTP6wGa44nmKdTGL6LwTv19fClKBQuH+xgQ9fOhkplWH9tBC2Nalf050OlS81O//
jjYbqXBfwHdIdU/VdAcZTmj48Aj9JJZOwRki+1/ePDGhehTR+Q91FwBhZtN+T+t5
n7DEOMLGgpQ72jSS9ZNEZXXE2itiZTciPkrs0hUA15j47XB3uBLmINM3zLRXc9dN
WxvD6vLSw2y+6tTzHRK8kaGhIDKImYqWtT8m9Pq+QMOGlCMh++H1rGT7qHBWVeRh
KQ9GF6sij0hweUgzVMVnleRFge/gNzwGvGymeXY2S7g8c0j7Flldwbz8NiMx1biM
Hp0kY3ZtMQpAvYto4v36W5wwGw7bNU2J3CA7ymQH7Nf/8c6aMm/jYjX28bbD52LO
4H/SpWbswo3lG3wIx9KnrdLGBshOZ1elKUyF1dKKwSwg/mvWpjxMBv+OUP4f+MO2
6+0IJhLFbqergv/e348M28cgTub44VKxwxlPwRN+3G3a/Pkh+K+yBa5mS2PHyehF
nMCXEu3ysR9sMZUIEoyBS+tX4g68qF/wEFboFA+8UficS8Pt6ShOb/eIRXVEGhZE
utwZU6c2uVaFWlh13YISDtg5x7zqKx6XoI009BawPWuNkIFX/uw1El1Orw48KrQi
au47+3vic+c2n5yXQfci3V74SPfl7Sr+ph/M1sDK+i9uJL8X92OYVSLqP2KV748C
oTwFL61EqdOnwkO2YfRbWf+wZgl0qapcE52U+MGFTsP8hYbvvVhXtcZc/DVqjgYw
9PjWEfgGBwzbdnREm+xd9BoA+gsOENWaB0jS7MKGd7oI0FD5YIdA/zx0ZZIjntHu
FYJiiFu1FKSRsBRV3+hX24QLog39WAsW2pjGIlUlLN90sRp2+aZweFpjES8ehh++
iDYEv+7kDbRT0zZikuBMsN7+ZdAW+VF+zQuvGevXTps4hIrVL3wsXg0i/dtw6FFL
mqjST2BNqYNRD58oKyWYKZm5sDb+1B1VKQrOUsVGwm/peqtjZMvgsguzYLoXwS9K
PaFM/DBTJRVWWnZsAOLNFkHm4kW0BM3NDQ6BDw7uXMLvbBOuWxDqaA8FmCaW+o/1
lZdPy6hOHfX0EyZtjgGb26Gr1XUOlAhLPHFv07+S8GjCC9tn6iqw7kYVsda/HD0D
/UNIq/kQMkYZyO1k5WQQdkMBWnJRRvtz789rpn7k4eOcKfoHjOjljJ60+m3JlU96
jjMD4n7u8lMyuqPf06sBG6HCLJ5Jl44ye8zzGjf+CGI+mbZmt1bEt56Do5N83Cka
Cv6L4GBiBjEhdVT1C0d7CTBiJH/piNaUoODYtcQKpSmx8Y1ZsSPv6ZaBNQTUBbb2
evZIr4xS14rPGqkjFXR3qtg8SRttrypEaFSe5qh7t3cX5cpzfXcNuuov/LuTvkJp
xs4paXSRtDxK32ANuunklotbP6gcbfLFg0vtBAphR34gwMYlvzsE6NG99XcyMSGL
pDVPrqhZfiQeyGpIF2Ii7C4JRdUIEDRUxeyiixpmO9KfmILOemwY08cEjRzA5qje
ZMb/MLHymBPM4O9iOBt7XwHfrDbCT6PpwgTuYhEMbgr4jMeC5eoNSEoSR8VxyiNP
BMFpmH8F/jC2gil3gIwHchm7UzuaqBAFNPbM3XdSGEkvpRsyEQGaG70BCeCm3M+e
loX0eBy+lflwv3dnJR3lTWotfzF2AeqqHpo+6omtuxen4dMehHfB7MHd+cTJs39p
LOBXU5BUI1QNdjIu9n2d4wYwiLtFawg3CVqO6G8989A0pRagFAL7EXFgac0sNOGX
7wWNl2WW+pQMCXG1/ePrpVuH/dxV4Hy6Nmnx0K0YNrW+pa7WnBXHp1nnSEbvjabz
2AM8agsCg4eta5vgvYdrhqz59Emt6b30SK4FbUwjN8JRglb9yeTIOryfu7AFc9HO
Nzj732GCEHY48EDKMX6G+7WKHDXnyrxXC6L1+jedzAtFdzSfkZ/aoHFD6K89fXmF
JDgpTRxTORRgK/HibXbzmGWk1wS5CqlVq+UCfiJUnbxPmxymAx7YSGOeriC/+fR8
4kqCK8m5KdvW1VqEKMczxQoIbULDFiKlcdeWaqAuPvBb1614TMFQw2T2veUS32Bl
HbNeYT1d4nz/NR2emmHGyVwpRM7Zq2hq4tHFiRhb+w62GAKxgpWR7/1EDKQ4Gdog
3zeje1nzvsmyevyp1Tr3e3T2IyQb1x4SvKu+lddTrLEszXGjKOO40Nv8aWXsrbiP
6MGJS4hBYyFLqX9oijHVlUfu8J/FpS9GxsnAWbRhXU2m11vNW3PyMQDl1ebWvVfH
APz7hZRXoIcSgj5ngxGiP0tQ/Fg2/gSXsrBi0BOlsqTSP56+opjGWYaD9NiWzBMS
jE1PlweZiK+HjoVYEjxDZYBjPf2up6/R2XRz5vsuGZldrsFpmwWPKj5Rlih3F0xI
RLhfP2FkC+wVq2/SuZ84tk+cD53+/mIkhXmNdP9duCAn9b2+nZIxushCEhboApVW
fxZltJfsR0Lq8i3E6UXQPkrW2Ww7udMCsmOVvNBDwh/aZ18FWTXu1u8DEK4cUFCi
QT+XjbyQJUWmisdfT9xBXnT2C4VJvvn9RoA/uEnhE6tVu7eis20PRxmvw3xfUP1i
opmSDKtHcO0vuGrYCbfxbl2EG549sdRDJoPN/BjFcxVkNRdG0Gd221ZRYFhfWIIA
yERRi+MQqZWKqWle/l8TaU0V0zvjsP/qxRuid5UlEdCb9sSpvezJnj+vkKbyyD7q
45ZBioHCxZG6NTCpSTxgJdkCgUw6sLjOUgX48fQpdu8w/e92Wj1Dkt+Pn/e81/Fu
YNfvQkpn6dzUHSGBjCCGfnyX5b+Zl9ueS71YWlDncoWWyb7oNz+s3JYQG2IujNEW
cpOxvR5534arSRQac847z5w8otdfP9JblNbho0nmcQ8XoRbwzJPGuqQshZbfjwzB
p2fQQB+YcQ4BfuCpocHJtTBouNTWBua5g32cqFzYDGE00ZmUP68JViPjqJl6c6dh
58d6zWqtVaoRSKFuG4sOZcxSFJcilwW5tWAB7el9Ybo/I8HaYGr0LL90pmzhWGoP
q81JJyFT4HThHR2sOuML8MOC5dJbe/OdhwFds7SO2OQxMo2ljUrOEOLsSiMUN7qM
mgDTsLmm/kim7Kt16MHyAopClJDVBzj57h8P4jw7FJjm4fUh8NspT/dTYEvbO4Ye
GceS1l1Ip1ssmNtV/L+mvZY7kSEt9JaHjznVxsz5eoEancHU/O3tTs93qcyf02Vf
LOPfGQ8FyVzr/zcjCuo1lG/aprL6ZmrCtns4SWrk6Kkqb6nYdseseNBWY5JfC9/S
qDL00UITxYdJL7krSMH1HeggRcK/COpVMp13ORn3NPd1+lGyfT3CQcIf9Jybd/9U
IKt2ylHQXM+sARoRhQu90DHaKhNNJKJdlyrIbYLZoK8jyUXdR71lDu8eX4Sr2TMs
J+pbQlIIm5Bec0W8pF6SaaCBOq4IypFNsxas2H9laZM1Ud50fxOYJ7u8wRcO3gj9
eLgGukIHB2kKbPj4j/iJdsph4bip0hbRimrvS4ZIv8EwEeP3iz9aVpO6eVWMCbYe
r9RZhiMkUpinvpsBGfReAYLsy5L3foiWQpVE7eiF1QigR8F9Zbhy/tTjZuWgoz4j
RiXHu0Cn0hbl6xJulkkB1mWx8i6WFAiNwzW8Z8bxNbgITRoVgkxq6FAv1Yr/v7aW
TxrNpPhJ/aGZMSwfWc74/EfkDp6cuPVfpXHPvni3L1RaXUD0xNqvbjhg47b0boPj
EavIYa7rzgheEUXwyLUlwGhaA6CAxxyG/+XpJBKA6ozFw77j49UOdRhDZvUFApVi
NRY5Xx741S4Mzg2L+CtLp2IVGA6+DTUh33XsJieG8Yk6lZ5n/GKsmG0fDznqVKTU
xnaA4i/al1qk27AsFXLrKeqBfz+hjATlfSaw8qUt1ZBykehhonoct1tFAJYTxXtI
OAmmSyIhqnL18YATVAEOqTVpwckZqUD0LctjvjvhwAZsl3hYo/i02NpVpml659Dj
8oA0Bc/p5qTFJ1y9YNzGf4fNwhE3PFPv7PDGPx6Z8EFMI9WqRkE28eOVUhZH7RrV
7/psXPS1LDQ0Q+z67jMirtYWiQtA9GgLJb6PjOHUwZYKbqbs0VdZj6k94674TBpD
1UVsRancfC3rkB/vPV6CW0+v5xuqnjuuqIsZTh0jXIAo7xLfFIhCnTD43kUIk1QZ
m6CUzFA9K6AQRZ144cqozMEuhdr4MHyXD59h5HtevDClNGZBkUXMY9fSUW2fQ+d7
zyuVPnwhhOK/Yq/jU/My+ARWMa8U12iwLjdl5jIuhcz9TmJApXxqfCp1aeq0iT7B
FK6Kl8i+7+qUP7Inb0R8UVQzl7+S2dT+OHJX8EqbWwHFdjRpx5VXd6MUP7gQc+EW
4mkJv49ajYRMcrmCJHVMBjbyWMCLNWhHaeEPTFx2TJ9NWNBkhsaz6/JGWf6S7WZ8
z7qT6h+/uTCMrjbqo0Hsw6y9saHKepwFal13dcA4o0ghYj3Y5fVDsWAFL5xcz2Ne
7hxbaqd46+8ngORdJIxUmycXN2YIqEem1qo7SkMriB31YAj3xcwCA/YWTuj1kQRz
g18DR40S/51wweeJtfjKmYrXYCtKlxE5W937w5Zm93zOa9hCc9fzeeqGa9mJ+hsE
usxNBjSBjTR+zZmmJzrbpZlQ3lsfnZumP8ZW4R+pltsL6GQKCoA1vw3XmGXDgWwF
+QVV5d3AvcSALOoqNKL1jTqH952HGuMLbH1EFjOzBcgmPc+NADrGP+OmcYW6qlzC
59csAhOSLODUdkxpFm4HElWYez6IQgN/4vJ6jbSSnr5Mn+spSizkVtZp6wcTurSn
szRdo5ADCt5hAskYxG3UU3g/fOfPE5fiyQXMZ8qi7tdULe/D11sa2MECcRynvRYc
JkdGKf3oMPN41JMND2u74K/iNzfLs8GAnoAOdulzA+zmz1ZcE8QBJBebDuy5lDYP
lA3YqF5SCZZJvcI8Q2ryP66NK12fLH97UF35j9AV/HFIyso0jEbcmAgKxeevOceQ
Pko/aWsfiovcSltHDB1r6uEJ6nUoyWQSx9STC6XS7abvKk1p0G7tkYVbHI0Wdjm2
bT2wEH/biZAQMPCuFDQyXn21DDseOa8IxRn1WVLpB/cMTGpwklE6p+ztG9IoIUG5
fu0eCjZu3AfaiC1lnEdaffyxQ8DboTqlpuwyfKzf75ATS55IUXzIuxFD+1CXnq/I
cs+Cw7GDrfpAO+ABSBaYDOpOV+d3qU7SRw9ZEUkSMD9dhuPuo0gGy9QMHXeh+y1C
XpxaK+k6dmQR0vVHBJxe7URsaavdQp8Xj4YcXDVZyakTFEUjFXRwksIpgLC/UmYX
lgTpjaaLWZ7EIGcDbA9zJ9htk8PvqohPfgAZXK4TG7EfYTvniLw2fwEG3zXhNGS4
sEDi/f2FbrWrTmp9nvNc/Zf3FfMz3s6ZnblGt/VGVcxX83ymVnV6bv6yz7jClcwc
Fn+rhhBqHesN1w2JOycyzYtb+tgBZ9I9J6mK1NerbT14lpjsHnwxami5mpnjC0Pd
ZaJpKZkc8/LxtRgRhFDTODWr7wTWTnVxpZhd1D6ga6e10nGGiqguHdTaJAvTP3QT
9Y3AjwTXqQFF41BQmeR/oq7V1rMOwgx2aZKTB5HQfGY5vB14jHQ7bOLBRUqdVZv+
u89gGezObdH0WNCdYBChWjmhoCD2m8DhT+gt2QtyhFTnbSC3hPyC8NCTfDWVuDJH
WwyZI59vZPEzddaAoq4/waLpVr6CRTCGml2X3MGWTRf5mMEk3dd7c1ICAnX2eQ1g
6CsTTiley7vPS+E+9OAKHQnkkPWLtpBjgZ3i8ZJOYN0YnYAgSAqn937JfuojZIB1
Vdn27znbiVIC1qlWMTWAjbsGoT27nAHy3vGSeLDq/3Mu4r7fYcuVuwX/CIvgetAI
fBFxfHtEjp1vMq3/KxBg8/suUH1r+qMQjrNR3ZLLdd/gD9hPdgPfA8HfrsM3ttT8
dXgPVQvV9026EpghMez5DvKujYfUvFnK+Ei426CpNGabFshH4XkIKqVn2tsixaSu
D7Mhgm0fRTmGtcNPcoJX2SQme3c7Z68n+KBG8yOklDghfK0dMHrMl9HNZ+qC21Nj
/RFwF9asIeWwWyvZuSFt+e8sRTKHXzwSWntY6As2faTKWlV1B5fSHvar6n2R098o
G8Fk1bowZA8MiGrrWOkWN0lcQK4ApivsEk3ClHSg4fd0Peftx8xCQYd08KageoSc
LsDtxpt36RpUEdGFiXh/xW8+qeB0oAYFJwDr7J6GUaWprGc+jzW8frI9Rnda8Ntk
GcPfBtiou3n8dXYXSZqaXm+AOl4jiOwI9LZ6EChn50APDt+8TZy1JCjirrKIrIzA
lZK1ahKvDXZJmVnW0Nno7yeJqx1cxo1zGuCKEF/VbUNm3ddh2+UlxNoqV/TUU497
zj+dBKQPRUpi/itwybQGLzhIqeKxRwCgrMs0If9H45kdTXgJsJjzl2SRNOojWIGN
QuFu7Eb0qwwn1/88wszW9X51XAI1lSqi6a3ncX+1GZb7YUnJIfig9IoolqtyeD0v
UTAL+WvX8kpFrVYyK3wY4f8ak78Rqr8CoPOalO0VCbLMbTuMtlqezM+MkyjwUoVO
dz9Cd1rogZX5hGPoVZdHZcy5XxqmTKlry2PhIIdzcJzIuOS1QSEasEi3KjEvRxF4
craEwhQl0ras8bw+J5rdtI2jjHRyl6a3uTjyIWftkurPEGu7eESQU+Oyeaj6OeHJ
zwgFcK6GYRSx8ZQMfPhV5U5xjOXzeNfy8YONf9M4L/MLjLiW/ong/uSPwdr3XCIP
ms/5P8z91oS46jBkbniNqSpKj5/+wKaWzylZqFP6mC4V9bc71ieOiXElhxAtErT+
oMq+Pm1YBdb57fuJIFvr3UsQYyCaCKLTiFPpq1Co6NGdwq3mAIgI7mJxv6CvlMrs
9lyjLfj6njYuNNQrgmsticcJpaSxgY24KNhbaqleEt9t//2Zgdc1zJiVW46UFiQv
eCCEkBseR5v0UkfdY6YSAkbtKgGvAuHDbkV9hn7D026FdgbU/tmp3+y1PTHuiPkQ
+JGQA2O1m1OEv5PVqftwXSo+I54ktlQJ2n3HZ6FgitCqQxJ8qx2GwyF717wO1tO2
S+NxmmBytN9nBJ+JFri+Gfc0pcdhnAz3ehSLkadJNKaZ+YDT1Bw3zXvfSta7Dmxm
Xyf+jkO4dk9Pz18fCfL6Mz2qQR2vu6dHZ5db6R/TC107FEhkvtAnSabjTFVGAzBs
G3keRAkB3Hsz6MxOp41T/zPVlJgVXVY5Tgyg1uSH+cVTYV3/BOM1LzBvUfy0JAVx
jG1Y1G0oZRKz4vD+6IH7YlLF6yv51nHXo9KqHrlBRYmLuSpzTqlC25+2Q5WNikJX
0Hl6BmEUCCgzQtu14Yk/jvudBZRcvAxSHlCFqq7huo69HtUwY/Th7tTYS9gvcxlI
Disg1xUlDGXXQGP6q3i2TSasFTKqZQtn+yQaF68w+5wkPtbNII9VguSdT4pHHA7B
IXd7szCYE13Xgufyrs0sPdBckQQTy4pzYmuJ3VeOKT8+ppBn1gGgcNdkf8KHBKSa
y1fpx9xtOYH3BWIt1n78M+IwYZvO9x/Laef/4o3TSrki+05ZyKRvG2A4Y+qu4aFc
F2i0MERcn58WpswvSrW7jjW8AO0evuq1VzTHiEmyz87NVQNJfhHMXEgUpnKl6gXe
SP0nwC2cxwW4/3R+u3anHtqmbWvt1Rr9qzPASjGFTPL3Dt1ai606GVY5skUtiRZK
5MSB5Z5jy9JLoZxTORRWE7xawncjIeanv4+O7k/PH/SWr5XFUuswMQVXxtiYiMAl
1xG+nOKZ/BXnfa95c14pk86RuZgsrHn3GRUoPN2TbfpGzy+pU8GC4AIm5ZkKYCOE
GAPrBAZQLdw1tCZa/UYNVHl0aibfaWdYqri9XoTSRTppLJkYuIEqk8zR2bJPFRrM
eGuH2QKetAiLnLP+5xJlNN446bx3sj+gPz7b6Hzdfr/1+/sBhTlqGBYRRIWj/62B
L/p9rDEXZFT5zQmkOqfQBXsiy+pqazpo1SfkX5Pm0Ar7RPt/0mN3JryRctdpQwLs
/VTyfP844SCNlhV9cgNbCl5misXO5JInie0upI42J+4bNP7CeSQUcNvnkGiMNyYj
4fj2zdbgqCzwFxxR82La+IjI89NAnfs0W0sHoexTaEwjkXinGMAuWTOOapFZa4vO
RQilkrwT75I1VuHUDo2tH2t7v5vLhB/+06M8iALC6SKhcYd87qxVn+IkLK6mX5hM
ej9Qngh/Rx0uft/53cnIwb9P3+o1/m3HcvKwTfCoyO2o4ejtG+rz3Oamuv+tZAeC
hplXE4jZ90Q6FealNPhrUsJdLYc3s65bmo05Cw+Ykdry1KAboVllEWNiZfiQ6V9P
Ktd26sGKxHs90mgDdL75WKQGy6c9O/mOjj/mrlmk2sUQXsBNSsc6GSznnL589Fi3
CWUYQ+2PZMSNKGtY0KWmu2lN/7kd8dPdg+fhjn4P0jvICSAkwlrf21kmuJR42aZh
CC57HVsZOud4GXe8f+dVbcXMqmUX4Rj3NwQdj5DtJZPVBFIUui2UdFqfKFtTLOYV
/sXTYuCyREEyrm2pxeIBOL9qOA5MuWEQv6Ma/PIdhhh93hHeKoQ/bgvUVQQxF13P
WTUgDfzlbH293FnbTitmvkwikCds9kStRqD+2sHaSNnr8KH+oGu50AKLxq5heRnJ
qfM6gBzLfeWhv4I8fkUW/qwXFzkLqkM/VH7A1Z1cvMBmmR7mWHIBNmJZIojbXpxt
ZxrQL1q2/k+T0qplpnHe0kL7zvWvlLhdVHSaa+nHgSaAGTFzTd+lgLBgxGHuD8m4
XqDLrA7bNAJptUignVLb7aZb4pweQb8eQ7+NRx91jyQdIg3A7DPrwS1yHfMjKiTO
Tj95tY3VAJEWK2/t3wzlhGWPwvf2kH8Wrtxre6pYIgxErtfmA39egnN4QKt1G1Rv
HiD9I9fSztjed8bfHOag0o/nSAoqG5ZciUPsvRPFLvK+6n72xO3whFkLuuudoU1+
Dq0h8EPi5NZJrAM7daIXc+ozQVIbYUqA2+94vNhcn7Gh8Yfr3qJcnTB2e4oFuusU
xqp3iLcpXeTGEAZ9Lv/FpLZhpsgmGnogWIqH4b7ALlcU0YmWe9ad54tWlBOM0WFZ
eiIpvCOA1fu/03abx1uO+9nWt4iz660VL8DmgsvdD3huxC7gSntfeIjIW8jd5IBi
Le2ERox3kihxX0uckBM762sGMdro4aDng61QOAfhcujygFT7PfCUOL/DVNKRVzz9
xBTZrCUiX8RdL4tX7arC7yloLU2K4/hE+xPPrlWQVv/43bDCtzHla+PHjbbw+EiA
5XLjsyIWILNMS7HfUP7mYiYcjAAEsmGVl/OMGRD+zLnOsSuwnofnJl1GsQUsX6GU
Atf8iKKZl2IbA0c4qkBed0twcLj4xCkK+oGDg0ZFO4rE0YH2Fd5yBVB6wlWFu8J9
+COi30ju3f7jxqTDx2GD9F5N2ORjR/03PKm2bG7W23xfHIDIdNgeBxufHNjWsqps
S3GnrKhKN648UrKxvucqGaEZpIHmY9E3mKvIU+E/1wq5n4YWrQCShfo+jxrT76fA
XaIqCw2Rgb1yZHphDiUvaQ2CbNqGKUnBz9aVUXdsavr79rEVnGX6anr78jiAyFdv
tDmdrf5T9DFjR79xZWBfS//H6KBBhp3dF0gNOQKvWIUd8fMWptq7Y9gdX1nkFeT4
CvKrMjhtpgo0h+0eP0d4VHo64ldc6zkgUONKVCAQJHEBFJxHrU9FhBB6mwOTmSY8
gir0KLqatQyCE5uwUeWyT0oARhmjWH2zKfVRyckXFVO1sm8tLwTYQhshOxA2ikwI
WgG1YIlt9TmuizoKSH/j/R/Qve0O3Vafk9DTLH2TLy4sAfweS+d+fgHnl2x0uyxi
YUERf9Kv4PH7hSigAQYvh+eAHYcTzWVrwETsedqMtlL2Hh9SNzBmrTEdr4DRiufB
8vsRYWlrGCcNiARfrC8AFRHVL9pIAAtybUXLMYSsDOsW3bQ+TJO4LY/b2oEIYnMx
yzL4aIEKpmozafNEvyO7VGyiDGn3m47AycYPKrjZyVp1iIX3TVuRUHxY1xUUGOCj
CQ7mmHqxylzgUzbDfum93Q+HsGE9ismrBJLVv+jA5/v+wKMpoZE9weqbvFiPoTc/
R9B3xztm8V8EjgH7gK/0Abxdjt19l/bTqC5P4nkZR7aF8JQiT0gZP/J1QLcaLVJR
S/hF6/fjPX2ok8FW5NstwS8Qxwirw2Ms09B58b29RmJrFG51U0ES+hM2jFm3xxTD
CkFWwgqfRTohuwR4pc3rxDDqJS6je6ndvim/pXlNHZVD7lHLKQq+heHco2v/s0pB
tKDTI7enkaB3eKIv3lcbaNJCMkTY8MYW55CvhQKLNmlhgRx1uVYKgWyeT08VeMSY
8yTOCiCtOH6B3JJdg/W0QCsJkPnZBby6xWvWWJY5bQgi8bGhdPXvMRIE1ZgQxzpc
NdXWRAKrC9kNZzSaLsp1cqGm5XdKpu+be4LdtCGC+kiLLuvJoUU9RUVf3AyC7IJa
N+gykdYg6kw8TPRw8TUqAqZKIiICTU09ua9QE4jWWvsCIbHTZtuFpbaSkL1XgxPc
HG62LMkFpityBNcs9RP12BpSj6qi08ePYWdCl/L2u3J+SdsI7Q47QYS4mmLY/K6x
zXEK/IjobR5xTTKOCxJ+Eq1HPe3GtiiH3qRkzOHPKSHitaQ+8sVgOG7BoUFM/o3T
vBMU3OSGOdG2jcZlTI+6jqJI5yI8B5j0Wn4aWmQ0vAAWdX3hAbnnfUEaaIcFNyxP
bxKK88GilsnEBitwzdqBFoTzkQjhiW+C12fBKGO8K5Vmm21UWf984RwPFRnZcFil
Ro8O8jrTIeGxfX5WH1e8D+wsZPXUFbDEXOuY5VXJDCfVKrKLcNPYNv9+5xRERjVU
W3K9ix+NeVnWVScGxCIiesT/OeiGEm+KwJ7/I2cPacwwxajW1DVlZoNfQt/fhP1g
Z5KXV3nj/vopFkU3OIYsCPTqA9oglQdYvz4PPkHiF4egIIy0IjAut80ThkQKwQz6
J0XTvllqGhExWhi93Dq4fZRPTQUXThTBbXQtFemWq4h1qh7vVMNdAxrHa6M1+1fe
YWA7eIWW2qUgIxNvCBS1OTtXQdjHPfcnLj2POGRLLa2grRQp+1RmwmtWKA0L2qtu
5NpluqgNSsCorXlRVpqc0/HDSDfIcBGbKdwYHarmtGOUZ09quLcGzmHx93BgBJ5W
TaI6rU9eIKTgublWSlx2VhMHyvHiXbNqcQ+4mZfhLxUA3QidXnd++yexyZtufKS1
tpVSaawebM5qxhurH5BafqqGHmyZzmNKzDDuS8D/+UYQw9OMSvB1Fk4CgJ/vh5Pq
ZeBncJA3KrGyB5ADBYAX/iGrkmax6EGTtEgxoU/fgwUmtBZQW1TEyyuV6ulzlkr4
sDn98RgOUf67v0e6p7njbbfm75VCJKEP6+jpr+74Z+eHa/HQ8FYcJPSLVmaTPrxM
kBElubUqULwtlBvUspDyMY5Dls1cwrRG3RVmlyU/ALqnXtL1TUwHoODRIpj0f37o
SWG9xLdPJezSf0iblFf8+LQuuo3t2tF2pLORzOkX/YPwjvzpXqgj2kFoQl/hhvn3
CmE4P/5x2FuP88H5luuMFsYmu4hneD9plg83zWmb9FS23zhjX0fqyjR+NFm4aRa2
/hzgoEzADoYLSZBiQ79IauhaDVlFctiq4OhLWjMIrLG12BUGjNDgXml+OyD4f3Ua
sWBeeU9DXdNpyFTb48X9J1JwPAXF/Ekq/HW4Bv9EwlBPBIKJqiH6WuXErkU4/8+L
BtTmk64tIMhl2kBrBS6M8MZIgtFVNXMgvtANQ1qKGItGP0rxmrlUGDgn58hdIzob
1SKZ+UKKQ1eakGAF59ACIbVMTFMKBhndEW7NB1TjOER2rt6LaJnc7oqkMbNZr0oj
65I6tt18HeR4RJqPDbZyAweiHUi6gBQN+iHd9qfmFa5Z2ADuys70J6ASZWxrAAME
/nVqWxv4yfTVauE93Y3S1rgdfiKgLD22ERcfQ/hyrIntJTin7aLEKUmzpZTTaGad
vw9ItUmGn4KOs9Et86wWGRUTRwsDoH5Sfqh6YcXC33KdFcDsNAfJevhRkirgTMI9
kZJRcr1VUQbQ+3PnwUm7rP9wYa6y3R/n2GZs9KQfUsJgsgQfE6S13uqnecHpUcsk
nffLhJrhrO1b+JRPwcN2CC48q6x/bE27R8UuMr18IxT5G7UuxgZz999vF+GV/42g
nPOCTYP3px2T1otT0CKnYRSZWcjH1P9kHMmywz8PpzCAIx3trBrViGHlUNq1TJXn
H4/yApo5uFVcRnw3MLitgfSJQpf3fhVIsS2xVUXhokvljeMfd+zuAW7zWvvcbtOt
8wZDhh/xiMZoLhDVGUupEEOyH9bsHjRsJeoiAbKC6F31Wi5cFaPlF+ALBvGyl+73
ZJOCYhN2RBzqLdZyXcqrhvTiVmRDMc2d6Hqda44qpiQQmN9I9lPLOTGsegurIPsj
h6PbgxxvlGbWPF9b8v7l7Qsh0lD6Umxp/w0hscqu2Q3MDKJjxZvALmwlYLggOFO8
HRG1+6iMHSHzXa+nl1dZidmh6qG5h1PIn52SxI7+XWFLZNisF6qufBnP3orvjzQy
5+eH7aDgut1UEytldlbVKfAvktL/nJfJs+tXgn+w0JLWsKuWAj+cT3B+T+cSqzIb
Tsn75wM108JGjrezRpqF3IDPTL3u9h2WcsCULMkUBLPxQE/G2zNb4dBeKWUXZR27
GggGbXyC6RzoGJLyE7fXBhXq7Qt/zVR5onW/YOl7oSQFIuY9uVKq/1nbo0scAJ2N
jHfcnYwukRPL5Aa4tA/NGYuDs1ZzAcLEJ/0V7wac5ManxHvGN2Tm6BeKJbj5a8BA
i/2AZdfSD7gKHgoQWm9U1i9GEMRwibyP7o9trYSGkTFJ+L9qWHAwitdzjzszux7a
ZXfxeeYRkBTLkZ6XtBeIE+7gnCK7gg0U5qJ/OuYLYKvpAIbsIhf5qkGHgbc0ob6j
ZirbehYCKB7de4kMEZB89UMbafYQxZrwtfwMPJ1taaGIqCCeys0ALVDQBzjPRcsQ
5Qo1+67iPjUn06ChUOKmbeNPkm/fWTWfb82PzX6zotHOoTvfy63UwRX1kjm5lEhN
X1BI4ldIxvR52L7HuoVqmiZ4aC08l6xZj9Hjc0Wr1SzJxpAqZgscx1I7H2J0u4oS
E9ZLjj4TX3+Zoem33lJf7N6OAhizvnZO3LnFrgC42+e6O408p4+YQDJWILqn5QPb
K10lj2wW1Q9jXs4Y4o1fizwFI3n2UGxG5Jvv8uKgQjY9P1upNrn0p0wiGP0Fhag/
9X6K6uYH7QzzofjbpgSJ2LzZUCa5xnndAUhLjSiI4dVhxKUgG6Vk0en64yzdqMtL
aLJu6dHF9R7dUFfjoJFZed8bq+wbs8MK9OhYJKIdJuenG7zZQyh5aS3t3pymRuFO
/nNEhnKtznTbINVxuvEQVoLCnvmpoIWtACtK8Ev/Q0HnaqkZB9UuzfG3Wi2r/fG6
fCcRpVJlJYhVM/eBs91HquvHlmNRC8QivC/ZcGmKuhvFK57sNcdcO8PJWCGmAI54
XdSWPasE3gFA4glur+5CQ2Nwt+JAJj1H7MAhddF3t8C6P5K1DW9IARkZsZRNRmsb
9kZ1rCoHcMed3Pau8iVGYXsUom2tBcnSHz3VzdUI6O78BDIczo528/80vJsUax+W
8OaOLFxqgqMsJ7Y64ZbVHMrwffej+r+lpV2lnXQyOjGiFuKqntGE9Tt87JeR6FjT
HsgeRZZSsv54XGtGCthniamiZw46kf982XcRxNIsv5f3/L7wEMhSk8/7Sobceqqc
t3fxsHDgj1tHP0oi3O0fVxVH4bWNVB5NfrKgaZ+O71pea0cEbeyPejt39zQOV+YY
G24wvh26a2l559VXVwKUYkd7nbE2eNmjMG3yXyOrt+zuX4VYeOhpyB+pY9BAKKBJ
IZsT6GwajYBFlqegvbx5zuyatzg35b5MdWi+9oxj9MWngBrOP33xDyyjt9/MK2Df
zNcx8VWzwFires/yoMwrUsxy8RYHSwPni1NjxUePERQkpL0YSW39yGAWzb6iGlgY
BRBoK9PRXBrbbRfmZitQIfKWXbIU7tiiMUe9XMUdLhjd4JQMrHHvJ6WYCDzzNg1T
caIX874slrOMVCZ/mThT5OcmOdRSmKCgOukbDgcIWdXxPI0rPtw6Q3EeeRHeA+Jd
5PA+gMTN2mHiJe+pEpIKAa9BIyenT+fb0EXu0O6g1AP+r6SB9ytxwVcIYMTPa1T6
SYrONmGzkVzTavSHH/cwPuva2UwAjIgr8tUqEqZC+kJIUdkXkNVOq9GikLJeL2jK
MZi0i57bUBumoX+/79+AB+N6PVT/5qvUtlVY3ObDxPvawBNQw1kaI7hLKkgDcK6e
hwq4nQeoYZfifZ2NtBAJNM7TpsFbXc4UiffZvtwoVWrqjIq3rbAn9ieTTgNCapcN
fSrY3x00bHgKxmA40GlHNu0ygh0oSbXR8JQyWslQJeGqOUYvbExwO+zTw4ZWGb1q
cms6HWH7nJ+YMZLllDFU7TQZjA8wr899ZAyHyjkbl/v24ceL5eR56wXufJJKHnav
WWzu6E16gLZwHYorDAjSPlR/a2kLSUS4FzS4QKMQo6YI7aMwp++NjJqYNDiUAyn1
MCxWdW+vAKJLYVmrtC63jjrAFj8v/bJ2Koe3twLppqqxRIRfSE5y7SYDjvgB7YAJ
XH2wR3/KgKUxiHwVLny/7hk1sG7G9vwydM+xz8KyLJUgvrbOxlP7hVrcE9veqru5
a2A3jZxxgPTWv4qXkCmgKynCP+dJFNJnbPGBPvhA1yu8VXDbZHFAiAluBuvl3UFG
Oa6mbg+sDMUHVLgPXHeZYWIgS5j4Q5jNlEugzl4oUpvml6w0Yjo5unATWcUriZqi
3ZJcaDkHodf59WP1qbE/7F0hwk/IkFjChgmLphWSaNzjT+gEWsXVkxxF90Pb8Qo/
OxaFIVzVcA2wqlna9UdLPo3FsnMQ76dmlCyGCLpvQdy9LjB5IG71xna48MVdzRRs
KQV+sn1MQkh+cxMWPoimDFAgYTtVkHMYatEhNu8NCrdONSC4/+jMf/NGiw/R/RsA
4HNOhb6OKqP5fMNvRzQXWPrreuI/LhKp6awDzMeNbkZE082cDHScPZZp01l0OhM7
yFA6MiQpohnEe2auSIjMNH5Ig2lJCY8fzByvjZXMowFXFax+byrNQNxcxwiuMtUN
64jSdmTY3tBAvtzZoji1q4Qhk6endt6KZE2WudQirDbMxsl7AxAMPP5hndtRCfWe
O4H4LeIgMDsbbg5DfAj913gOelMfjefxpwF50J+RoqvXSdF7aCW/ufLRuXrN6+x3
cXl2buNJP9MlR2xYnjmDmg/+A5FLjb483mcVZkVWdtz8yDpApP61QAJM3Yomu3n8
WwZDFo6FsoH2Pn0knJ2jgFO8Bkuz9lX3fE5Ky4epWn1uRvyKAXu5p1Mg1tFrzZDI
7wt5EXnHXEXF27OI6Na8cg/JodRqAy8gCi+UzKZg3878bvmaVjG/ic9JItDhUpLm
o8dokkvsAybN+LllnNw4ykj5VSDrSFJ+oDDj/E6N1/HpPCcV1L4qJODWCx5CVupC
+wDybhRYyXYtcVkANFUDiOpKKwatN3XFxFVoGKLlVDbJM+4ZJF0P7QL5hhiG9ezO
+CtQkQGXeWOl42kNIFG64O4f2sAb7P4SO7k10Wt5qSjVTwR/xuNpBUN90yR7k8pp
JNfDGpsjzWMj8wXqKBVU2UCI83ePaaUxSu4ar451X3vGGdJirW+/KmFBa2A7IPIg
5NugY+xSlyciJhfMe/4oo03/h+lsf/SXAQyay0Z1DK+bqopDeFuMhU7t480erSpl
PuIFu5vaVP6eW60EQG/7o+5hkjzGjMW3K31JbB/k/XqbKU0jkobA3DFvRXc++GnE
8pLSueKDJHLeD0a/3vG/4DaCY7ugyp6entdxSHZaIa/GjdmBlVgiiEcujEeFmJyv
OaUMGBAie8U+W9pDs66aTEoMxGl0ms3JWJQxPcX8+q4caFOhHY2sA64S7UXZMfPa
6gS62f9GzrPGpoiYz9xw2mgthgwJ1eX2K1WAeUkpyooXqHw/FWymQyhwtStQ2WR7
RtVleRpp9eZzsMQz4vqAmsyP8jei+I3tvDyads4stuvcg8vAsWnvva3K5uM4NJjK
1ZJbdiBOzRxA+SwvpTgR/FUyTNWuepRjp5z0tTenoUYtKAGiT6KxlUA9QLQukrI6
sCkV5cK5x27OrLNI2uo1ImX8liXKXxVpkIMe1bhq3aHkNQeUvYU1dZjSrUSCHX37
J0XJFdmchWeFosuUSYH3INGt48S3rXhZ7YkLFX49ShxatppsTFhG+p1UityOxN8e
ZPqUYA4I6YfH0LftGazmH29CXuPXph6OGjs+oCi71caacpFSftVAnJXZZ52Up0lf
uwjW5F4T6WJDvQZZbKrDtlRxXz2O0C2nJ3HAL1oxKHjxWo1davAJJvOUTjaLEbTZ
Jv5uEAZ+bbwUja5eM6xssBTjk96pxMjp8/iZpo8D/PMOeLS9vt77G73VB/R38Vjq
p5jlN7lDjcoEYF3QEHRI/b8xQ409WyZBtitt8l5/2ullP/qXzkGve/prgBKKqPgN
0iCroq58hm5MANNj3UWUdEY7P2AoEev2Qm36EqmM2FguDHm1vJ99LKBMWllwRLRg
txoLZD+ESsTq7FXrAoDWw4vj2HZfVSv2KSfThuBPQa4mpFxXOnT/DATee4HInD6c
I/7o5/hXAYx49lsNk12vJvNGoqE2gMHkAx20ml0bMous8D/RXQDtLJEo/Wopra0l
MHJJ9J1o7pC9kGqzxsmdiOHh/v24YXAtKfL7crLdCbgrfCLYaoV96zV2Ygm36IYO
IIcvd/pNt6O+MSCp9FpXjpK+GWOtC1lDJH4w4eBEBudMhZwhj3yxouN+OCbzEkcx
EMKTHKgaNLKvivTS7Ktb+K2tMqEf69R0Kdp23lh0MB+wvrrs9mDXRBlTrYu29BaQ
oX4s+0PONpJLRwRGCObIWJMy0VdD4IWPXT+0yt07V39jRkMWii/95Bw0uaN5Dtfq
DAoO75030Xfd0K/EwnmjN1yC3a2m7OU1O86roiVAdKmJNBhrDfPUqLRTwCwAOskv
A8nIn93CkndIWmhEGmfY4cuURwywGb3Hsv8mi/gZNdVAev/cLd0NpvwI5yUQOz+B
jOGB2Ufel2wTlKHer8gsOHnYZPJ0QGrpSjBxddWNwokUhUtmE/BPPhxDVsvkAARf
t/JBSoS9KRN5+CSdQjtCf/3YKIpdf4zWl5eVKFOqraZt8umV+0AyQF/BOfWSfQ1J
njxaP1k/onppbnQwJxz+/NPY42QYOBaIYgxO1/ZD5Wyii9P7O4ZkEXxCuG8aGpPj
EFZcwT+pdB88Tvgq5H32Fdb/c9q6nKiINP6b4dK/AkZg3WdVIw6O1lzxvrukTDHs
c0MbOv0Fxb/FxkxU5lSkUctLVM7ydKM0OLqfpKn4d70g9z0//uLN9sbC9YpRmpK4
ngQuXfWyVaDFnOeHbilyAAbE5pDEGcMgxm6AORFHRH67SXp5WcKXfy208DnjPvGU
r5NB9ZP0BbI6wXHKhpX8PPjdM1Bv1HkzDTsG4qDIF9cPGKn58ktxh4Pn4JoOe3sJ
D7MadYljSsPv8U6T/Q6EIg6b/yC/Ewf/RxBXsGr1YNjlWrokWZRnDl0D5MS95T7t
WdRRy9l5i5k1iElHUOFzQH28EmsckCBsF/7pOFuA6pAd5LltRiAc/23kMiitFqAK
r5TT5besp46lCM3oCxO7xdgUbOrUK0MK+f+2pP9Xftl+y6MGzCExd3cedcVPXBv0
zu8/FOWuz7oH1ad+cHfzhXwiBsFKCQKVeiev3wNIKj7dq5cree6hYGt1Q+Cd93Bl
EqjPNyC9i4OdL3En+QZ95tse1bwhkXBNjhpj8I9KrkfuERpQRCAirshdkyYbQUzm
WPm/Xh6Rat51sPL9YTM1siLlwExwhxHr6WJFuTwAufjlENdxMjDC6BVm3Kq1kdS7
+KZbjBX/K3LZCm+Qg0G3SDdkIKlwNcExKef76ggwzhvjPswJEoYxDGMF9qKuUC6r
SMIHYLctnIb1ZT8YzTnmCmZ0u4xN6ioMaifjz2vLk+Lyt4urxm3u0qd5b2EuDUb+
K3pDrs45au7R/rWnnePoZxEaVSyV2fAxV5VZlho2UKJRz0KzbJqLXclOeJNQ7Zjt
u/8K1mHuwbYsunGoZ1pXMQEhCpo640a9wvV5Kb1CXszi3Q6d/aHWw76LCG04tSeo
+a5gITuNHykUUtFQoyjB1CjeKfrEwL0Rdfk1r5P9sDC+x95O5+lhdE9wqrsRmHDr
+gd83zrPr/sZ4W5ct6v0MDvNGo15MyYhEDLYUum3fjZ4IWEKFnKe5F+r8+/D8yXC
iais/FNdbfdui29jW9arQDILboAwWuLv0tEEVT+aoy+L2wMT32Bt/uU3gA8Aoj/M
Y9QJTg23KNOiFlmhkFyuBpvLp7OoD8SKc7c/Qd1ONnb19U9Bdaze9huDi4t8dZfo
v7WIdvFr4YV9cBze0DwT8vONNp1/B4cFbV/UP4QJFcZ4P9yc7PXeaxgjzrKXeFyC
vKPuaz+ZPg1xq/q+0ofpuMMf7znEH27MP5Ihq1Vo4Lo+AYwafrXwGQzXEX36eyVC
QAfftIslZ/00+xGD0Kq8uuB/NG+xYl9OmjqNb3WXDguP43zQvX514tMmIfu7J4sN
AreYnPFbUIB/eI4GoyKdyvWoOLlsygycIAkB1xePZTm28qv1h6A3XUMPMfC7/Mtu
0lzLD2aHzDjOOTef5Ge4FxW3nwmsfMVEXQlXapFpE00SQkjUvbQLnB9v9KfMq3/g
cNrqi9BDXnHVJUN9TuHY/jl1PY70/O0i7RBYAXX1t2T6EVe50LH8mVPeU1EBVyuo
Va6TQsrjMAee/khyl9rvhNJvmt+CKdoEmYrXu1K+FA2SWgLKXqvfB6dsgF/MrKjw
AmrKgdal4yDOoTnS0asxYbC9PPkoaQ8p2V5tLDLLGzha/fnYY2l8lqQYPGBJSqON
l8PS4ydlK6jOIomvQgEVGiP+qdRzmmsCdUE0cTfxBgDl8MiMKEaeRd+wk6QmPFvf
Sh2vKyboO/PcfQ31K+noJxPdfY6aZ3JFXY9SfUhnaAsd9FSmsaP2c8g9GjQVEpIV
vdD+cJ9pZoaq+A0VvDGeL2BGKnGn4k+O16WhHaAnKLfsFqsU4M8WWxaFPbFoZv3E
SunS5ysdQQOStVDK3GkCIyoRQAgNMP7D4AO1jc/NqpA6Mg7MssFd5NxILrGGXBwi
P27Rkg6rcb+vhRmCG84uDFVWVnYN+hI8+JLwCd80zOd7e4P85wcQ1CNbUNBjIPth
wk+t3fa8CU1N751El0S+n6AhbjL9ZsAFTsSSZw2a3IFLhGTAwpjxeWL3jeuTLfNR
ZCuBezsn4mwq76GbjKMBnp5b7mIrio+Pj7FT6eUu6B3x+bFWU3M9ztLLNoM9b9Rh
xbjrDhnt0/svXiyusXBsRwCGAMxJyXVUAAKr2yybmNzh5t/1d5dkDS5Hh9ufd9Kd
+gV/59O1KYglnJ+enN88RKm8091C/NJ62zh7nIHTkHhPM1FYP7FvT1qkK+QDsPqA
lhCXBvOJaVNr5QjpHVxj6w2XckjL5UC9FnWIT7PMYaMcLUExDi72jGny32qkM45M
KFlMP1dJuwf+dUO1MVIubausRm7/F9jnSp4uYV4P2bpwgj0pOkPAUI741e/xks/1
+YeaJWWcfBVc1fW/N4VW4rSO3vQYqk5uCF3gmn6CAOn/m4ZbpmZ2MOf7mkKQsIM1
MPMfGPWwkSq1RmCCQ2TXE7i9vjee4uJShNep8WDKULY2k3Rkgn3wFOb3N0C5W8vP
89WnZs+rcXGYk4DGUtetGCHoLEPMnaLt/gqjEZJt6ndt6ZqP6py0kn/2neWAa/na
AePn26lV3PyhLhkorVE1h0u50Ib0NKAc91PJmbkB1D9tCGA4D62ETwLCl3oMcOCi
Q/ClJ/V9cL5eI1bdXvhjGDtES+h4NXe8CsGOID0VTBqg/ZBjeQ/nalGAalBYNs8U
UYOR72nDJEsYle1I0+ZlYMsHAj5CqR9t331p2QAc9+SKn595KxQ0NT7iCnvtSP5H
RUKnjwJ8rf4edKj7wiUs8hjf0rg+40XK2Pv/N2ybKosWeTVOTUQgMFIRmYeIznjm
a3OOcuq8iC5ku+OANcSnwJusXN89BFu1NsARHG/pHHgkqLNRuLHCI23oalHE1msG
cdpTqcPQz0tbR70YU2cmts0A8KhFxRmYt1VQMhPzwu9UkpQGr0L1qH1e/CUv02Qb
n67sYhFm2krgr9DqxmDWpYZgbyGUfYMAbKxCBjQaykHe0S53rLv2MT93u7UQKIUN
yDAfVL3LKsba5eRV2hlGKnUo4k+uTwjvDsF+Jnj/JLBnxF+CyVBOITEaUAIB2oU5
wKBkB5IPBi33mM+zUcGJvvUUqsgpopfsloGK+PCfxjBeYGvA/GKRiYdARUEVJW8N
AkQHFgZCGed7T9IGvfQ7YI16luKBQDK7AkEr9KYHXZfrx50WYXJ4PspQVDjUNiMk
5dOiXK+xpE3dGqf2vszGaNT3ZwSTxbPdmTGE+tjcZaTsqA03nrelCvvRzTCnI7u/
s0f0VLtX5rUbFicKTU5S/uynOoJ66uipZlFUx/8GEEs/lMgSKESpXb/pAuI6tC5b
HbgvsjWCa8hVPR15Ka6y1/4C4rnvZwQZ4rsomWa6FYsldCuS/FitlCO5pLe95JXy
x+jPD/q/5ZPsZPzCY8yk9oquMY1ysgshzaAqaSi1BMxZfZgoCncDFL+1seH/dCd5
1bMdrfP0zIhXFQX92rUMcW8rO9iXNYqZQulUhkDhdBR/k/vXDDI7hFG7n48sTuT6
hMbv5+sfO6DFzgE0+Syj6rXw7l3IokNolOaW69mYDAHsM3+dCZDxr3UIFE840t1Q
p8SYf1XJSZkhp6wpxSNU1VBaHp7XwkzNO+q5tVFA+yD/GsjT2pt2QZt+/Wn+xjWO
77+5VsAtyQOqhAJ49BoPfCLvKuScu+cIMlSs3rHjixj3qXOV6ngDbIkG+6I/qPn0
O3FUOkSOPiDT+xMVm/wSi83eUZD8zcc+sIwM7+BwIVTN7VVZpXjyuwk2NscNzwxD
vCU1hj9haise0ZTANWi3DKZU3yzhIXFfyz6xNTRVxH4g4tUNtpGHT/6uPl8kYCvp
mAaiB1xf/ytNo9i2N8T1DaH6+B68B+N9GNkZZs1JKZkJ2yuJgG6glXGxN2oF0+5E
o1GVDcp+PY/S0VlKUynfIo1DSCXduCImrPSJYrZ6B74rkFkiBikK1VSr5FMedb/T
Li214M8KypDG4nhEsViO9TI03BciK80UQIC1iQWG4tyTzgnrSO4inA1UE46GYWEV
aa7XbpD+ru7lQy5Ncv4X4PfyEoLHTgYa1t+2fq3L01PKOpdrzCmqLk0zeBzasZTP
hQKd2WgNwTT6nKpexPC+jg5nuPwsRm1j8qHHyXPDQIQsLFLelSLi0f2cBIsYFKmz
Fnvxe1jn94Yza6eG7peiAE7+O+7iukjM5hid05jys5caRn68JgW88gCuEpZ5aWVh
NMkr85GOkIzqkC1FjT1CarWYW9zlLdKqWQy9sib7T8SVwQGnDy1fUsUuJ/75s+bE
GOxqL8sij5p2u3TDr4N9chVCDbL0SCnU3dN/vVXih0hHtMOBa2UokMUIC7IuRm18
1B+qwdwziI72vkD3eHeE/TJjpZWAOWg89FIwowRfXnoddh9w6Jwv0xkPYTHiLRAB
eP+Ycl53O/OnfDP6Gd8MjLoG2H4+xrOKsjJN6oOpBEYlxcQbkP4G8zV2GSO7uy6C
P2Av6/8K5+4dKO1KgRCxQSCXWLgoBi8kLcGp2nQ8HK9dbaZdsoi5yVi4J8T2J4fc
eSYuFhgLlsgvU8F1z9a1zsycCl8aEh4/La9tMGLupjJFvdsptTGsltV2TnNHh8ar
t39ChKaedPbmi5IlGgyG51uSomNvHCAzarXJ9mhdr6EsIncIWGmQhzwF/al/tK/C
k0Gs1+H0l+DdzLfA9TbF7nSVUQBqGk4LRpVqzMFSOhZxMKU82CvqRDYJxweDJ4WG
hdt/0rY9HJgGL7uukFqXBfSVS07HerSsnd6ZwlBWFgASUhBflgC6us77sQYFXvIe
wnby2sFFVLC74CRAN2OTVNpZkhZB0bIw96rIuWlml1sZmDe/x1BfUGj+QD1h2n4U
9xRNIqBAG0KptK1E9aIM7FCGhUlLh/NDmyGXkPbIizJ7wKZv+3gwLdIlVrT+Pop5
k3IRJ0NO1/MNfwhYOMO+TV488OB23i2iSzTtZhAPZE0072yG5uu3tchl0T48gvoh
scuRsBz2Txe/1+jeHEchEnHrmL/gd5yDKPNnvTQLnHptVVGo+z0XUGBV/TrFnOwt
pYbsDPbsXBM4x23vJflEOwLiK9TYwnWipK3GWyNkEbOxB3t/vXiwRzNfM8eBKZNI
gDCiiPfKLgxYOuRzn3GlnZrx91zIEE4nBcHHBQ3yM93PwiYna8p/bASxzVZFBJOg
0qMphtIfjqI9pqKu6PjBWqtOXF7mjNtRq9EEq9dHL0AmsWAqx/yw7568eY7h+y0s
Ekp4yWjrEb5LJFh4nyJkHl/yomYDOBEQFvVDRrmWq8RdTmh5ciMZshXQ2YRkMV7o
Zb2RYkruoTCMqsfjthiw7X3atF6CUScYIH5FG41P49RmblpN3pAqZ+dgfv968XyW
0dAJGaNHE0wz+QX8Z7hshwFce+TWfwyI6g9LoNQnv+tcHwB+tt5nQQIgKLHAdA5n
4RrOuO8zABTzWG0hV1g4rb43nu6LMszB5RNt0fff7HIqLQxFSL2czOXODdWcFo9G
r1isBV9dq5+Gv0kkMO0X/0sXcvYqsFOMxE3N0iYruWFQ2VjbMIpUjDWVp5FUaZzC
P1+UySFNmoegMRwmB1nTJPFy+uW7Vd6u3r/qhFgVna+PsWUC0pBJT6jSdTPsnI4Y
4+72pzoBECeW9pS4Hewv16fvJqlnekkz26yEdAU0e5KqXIyt1qIoSrO3V0Y6XhaU
Hdr/nCdZWf4pHnjqxFk76x+OqCxp+Q2gNzMUeyq88jQKjggjC+tRBtDNPn38/8Fv
rl++ZSmztQ1l6fujwxYdqyV6AjSfsH2rkY1q56wqU0fInYIAEoEperS5d7tN/yw6
h6X+im23eXPPcOeYIxaRWshmpOq92w8ZmkqF7O8AW2Oja9GWVmQVm/oTPerwABDr
IS5/Qq2VD6hUb1xIFzQ0IE2hD/SWBQoRKVSxo0EyQxlVWV+lQi7VG5wyLcQvJF3I
4WTrG+tZiRlfp/uukW1/ySaIGocAOpev03X0VNdBJCkCcjfopfLfJ5Pxk+l9Yd7b
ZysNJnhHXmwJWeTue/BSkOhROwMWpLUykz1MbPw64mFPAjC7vtl324sg+9ayEhLQ
E2vtW4D+ECo4tUnNrvZ+SdmFdPuMyUuGo3wJt2hc44LygW8etaEVb/uKALtTFMCC
YklQPxkvQ5TBxEBZT+uWY54Zt7miJ488EtmyIRSACfQzfd+59dwINVQQ4n0EdqNF
uOze3K5jEF1DPWNXingm3yMn9VYo9vFHUgzgagFewWlcOxsEb0gMBFXEay2eWfSg
hp49k7vQ5ZJirHY9Rn1diXyJsJWxpY1TzIIisqIqiVwlYHsXok9j9PpCPFE8ncnn
gBBV1s5rRbn1ubSxOwUekR1w7ij/asH0csnyKo5xPTYjuAiUP9GgJ0vTZTF3OMEh
Ufn7UXqfEuDz4YemgIcqVmAPSH7X+kSOtGcUY2GpCKdW1P/GtUYqpioUHhNtXCaU
GuW6MWQvgHFZQslBa1RN7L9bvk3XkCpCihv+RfDsnShjvorEuEanG6Xr0gf9va+c
h2XLq5JoZZIKsr2FME9lMci3mQF4++iNq0b6dUd8Mu9qbHAZeefw99hLGqN84Y7v
lwtkQzZKda37TXUzQF0sqZt0Jsj3YbpT5KR8EItbLXudN5JSHHJ2sZNtn4ZEBO5V
qMbUiSyEnBTFaGrdOongdeT+Qpbvuo1BzE/bljZiWThX6dVNGw15eazURvj8jlp/
Ec8bQklIIeXBwXw/USuIB9Vy5NkfgcGECr1C3oRgDJWdCXr6eLILqp85zlv7jH0v
Pk7CTxJAcKgAc5xd9Pmud/+O7EVl/rbSkU+rpbUSBzBRtxDLtaCq/yK6GXvRxPr9
hQNu6aL2Q+XvLChhq894KoqC6fWSdoIZ0hr4fDo1oxn9pi5b8qEd6zcho39UkWvJ
R/tDNXaXiAxTbLdz+SvPaQZz6MXFMoyJd2mZcx2C6IXWV/HDyLs2U1qj9iqsy08B
gIoRgJh64jhi5OBAiIupmH659EnCpb9zeGdyjmDyvPdVubduS2Sb+Z7ZR6/bf0DD
G3juEfgxh38nNkVv5AW/g9es7TENL6gSg0FMfkopvhw8b5jT0CzyjnaVnUwk5SC0
PNeFCwvyZ86Mkx5yQ0mHM7FsJdsn73Xoo94D/vb0ua3rxlb5guTHIfcLIUxIAkue
uUfyv9mpkQ+gtBQAc1z9V1FDo6Psux6u8hcdLQXYldEwnCjuEQoKnXioyTxRwhJA
wnpkgYbSqcDGAj/tNrrqC4gNGT+Xm7h+caUcEnECwAzYOMBiycJszGuXRfqH65iK
zIi1UnIUSRV57CFMNA6f452C1Hgi/H2hmSGXl+t5Gtgl5XR8C4swlupES/siVMP6
DJMaF29utdfTktdNqrh1BCVsPT+Cyts8br+OPrjB5VvPUq8xGnsSpu8apnwKe0ib
mUFwpz8dN3lUPthViTsoK2/uGmwYKiRMhjRx/XzAJaOdFkgfcSDZdkNRBGGpR6XC
GthnxhSXmGcQMTe3NbeoWTX9DIUNbMxa8UoR6ec1niZ9JxgmJNtgzeVdq0++bvbv
UbsxLxy+YitX4M+F92FOW/Sbh9Sha+VgGAR57fuLSyOQNYbZ8fJwS7jTM12qzeff
yzD//tr/QgPHdD/RMZOnM+jyem86g1sgMt/7A/LFP7Y1D/MBJ75qWIBEvNemxQpm
XRSnMkz+R4i8XakzhLbbCJjD3wTArGIQd2Q8622lpuo2iPx4Euf4jGQD/IOO0+g3
+TFUbxvZ+LOP7engD6f0XIxGMjRs/JgjSQ5RuvmmP5FnB0ge4PILJCxdITpahYDl
fsYxgFimlpR8gjp99zjLqbRfAa/WwunE3ceF313hd2BWPvlDb21aYLJW5TFacO5G
tmIGFzJPtOv9NmZdmYuIQ4GMQvX86RQNTNfxrdPDPHsfk1ZzZ+AdX5YOZa5sr9zA
vG97QHrz8TV80ySNPYW6HEoUaSuXYe9i0S2qi19Rg/+YubEpuFIHDIsDHJpUeq1y
qjsc68685Hzypm7Y7wOEUTVaFLFwXmLIAVVA3sAZVFaNw4+fYRFRo6NT8VFEXedH
a1eWpqR3avd6KxLWqueNCJgA+jTlQHotUsAY6sGkhm4viOljrYnjuGtfKa7NfEAI
ANVQ2BFYpteUu+inQ+4oemDA8iXe45md1srW4g18zcQjNsJe8EUpnlBJmpP6nOjH
UIJUIwa4UkZXpnZl1a9qi7Pxw5t+bYdXiRMLIqWPTrXbBOqrLa8sPbAh3Hvy6rZL
YzqIKeOGIRizR+BfG207UZy4rwD7dX/YI9bl4YRWlIc3kl0aZO2A798ObJsLrKDM
6A3ZgSt8X+qIHt7rRejUi93sN8YvaAOybr4EAuVJZnB1x9nf00AF0Cegoy3To2Nb
nlY3scjPQIUKxc4HWizBogn+Ypg7jrDjgHcGBRQ9kcMTBKr6X+pQRC0bncIkfrdh
tZTeCvDCNA97+en1IRauE1lvOARK6CMC+mUeJGHpa5vk2+qO723N1J5D6CX08kHM
CYt8tJOncj7PwRvHTzNR8LErj4PqJuwcb1kmqpja7+KERHpAgK0Eaf7Xzrg9GxXz
h+QmQ1MDLSbNUYgAeXgKcoT6fiswWVzGnbIN+SrMB5c70XAxIuZxCvZRCFuMj1jx
ER9ZjWhscOGSN73JnC+iGQ709XyElDrMioPTfbvteYeWAx20PdiC8kLRtaXztYnK
J3RlcGruZhW8QzDNquuxMiim2qPitUlcnd739vkAH0bty06kfB/Gy6cIUJMQuyUb
rqxQM47cNM3trpyJ0oKHlgo9Ahkv4YzbXRMT7LXaukvnSsSAvqTB9bZ36LXeKLKl
N5J0FY1XTh4KXt2N3AVIA8gL/6o1UZXJMdlq8+kiXjce2sg2tJWR7H0c2Jrn1n6I
NHFmo1V42aU4yPVVP7iivGx897utjlc2qAZHKnm66aIg0nMXqIPfEpp79gN33/wg
9bwjMt29kMP4cU49XKR0qQyhgzzSxNkIJHOJgNdVcwtI+kuY/vRh6n6J/kgEgY0Z
WetAjq+cL0DF18Cg7DfCLMRXgawpeb784Bk57xg0RR/ixyHU98k2WpAJMYCBWc1p
h1ava+OuBQvHyGyqj5LVoy5o9zz+3br6S4Zc3NQL14jBeD38sle0ZY0a0d4LmAD4
3/j3rj+jj/TtTcWuY0DnWtzsS5vFf9WqPviTHMsW6RY9sNATb40W/vL3+K6yc4KQ
TkzQvx0FrtSqXMz5nkTd+dymuaJnr/WNU28rrrMJBD/eoDHXjI8UNIlZJ9fROCMP
NP0ajnHCbf26UTYgwFSrRpvxyR1U6KyZlGoLeutSKEgkq0tIsW6FXm4//UA84TR8
dT+8glOdbx/B9wJU7v3DVdohVWBKuM+NhWEgvArEGGVHv0GQhqcUb/81zv/+m1BP
AFdBu5Pb3Mrafq4Uq70UiNlVOpJ88mB5LSC+KiGL4nd2UplHoyXCjj99/tJRnR6L
mwtyL/I6eb3pugxraB8vJbVTZA3QZBW7cO5LgBe+b4/GVgZt42Nlo430mODdD+fN
vY+ja4/dnIdZAN3GsjoNYXWgrzGf8GoiYJ2lkaaALSQIiZPamxREc8V9mhk0qX0x
/2NQ3vpRSAongQRCXp8L0p/cKZGsZ/mZfgdQl/cxstVCDZhdo7kzdT5+tPOOIz8D
W/1i+gR+kGAAT2+G+yQxlNvwTIa7kkkYL3oVnkuZdgKd5hpQkLZ87BFAbJaq2Mi/
LjadJ24PjmNl381D27aXJcRImBGpCo1k18RUT0+7biZdjrGlBdMeBC9R9vc7viJ+
yQaeoXoCbNG1G8Wx2wfK9mFEhN7ntL4gbTfXqh+pFzbLVC6lRmxXfBuHEs2GpvHI
SG3SXnU1LcUEm2H00qBsqiNyKS5LPENu7MENYHa/LAOQ8pCsgnPT5GJuguEDgFtA
ScNH55vCT1O1wRYN6Csn6mX1KEeMNGGBmHRPvOeMMLkSe4ml2g7AjuZo75nt+bL0
0FDPXxMP4kG8xwJ7jlNevX0v89FzuPDl6oOBEjxSc1IvfJk4u91J90kSSdXVVpAc
iruQlLJAZ5Vu5ur1pfN+WtWXlh71vY57riw72CbyaiCwKohK2sglU+iNy7lBuAuL
PH6QdT23DukW4LfJtk/wAhLEqxKJAwunk/XsdJgITB2+LDMqHnxIMsWshN3iavh+
Nk2JksAvp6PWCIDyGRyLTd3LRkenFlmh77vCI7XSThPriU9r9UKmVCFK0SMwd0wt
fk0Ee35FPFUk1W169SyZkwvx4bwrpe7cQCCaBgWcLR59PkCdfWdAF21XTP6YqRl4
RiS+YwJCEpAq+aMSHTJDtGIu5tup0Y7RHHU33UN3h6tneaailiDMEXHUtIAwtjMl
kolrT6Y2TBQC3rrknol3qnCTHe85wu5+BEtIhdgKwI8/HZSbnDdkrqlZq0Vt/ATQ
RXKeoQh+252Uk8fp8d7FYH78W2m2axQzhZGHb+QrYm9JNapbclmhu5a1rw51Ep/h
SvBVyJ12MIFK2FMUF/3kNaiWwamwOz9Jj8YeSigGlIkfaboc+pAmE1LHnZkel6HB
2UxKYQ1TZ6ss+EkwVhExU8P7a9reNc46R94oIYoPH3jg31L4TfbYkzbJPM7Aj7H7
Tgfp0y2diWJLs3tV6akIeLxBipSJnJL6wWUNegS9T9pSIKrrnhm1UOw93I3fVqTY
psjj0LCtXIM6ewn6gV+hV0ZfG/l46MQd6WuNdlMI//ytCDhmEXjr/Xk4NNooNYgh
fjFojd7I4/IpMWnZ5jSCeMtq78UKbSVcIgF+0Ccg0ztKuqqUJNs8IsMLyreDruXB
Pi3Y+6cuc9zXBsHPEuZ0oZpzXvMgHwp1KHjw9rlJpowA4nmPxKCSm9t61WmvSPNV
crdumtqByTqPaeAS5SwiawrNDHzH+nME+RsVh68/C8gjiPmCI/gLc0LB3qxD12Nu
GhspiCEiBYtnPOZoQdncaA/oD+6xXCfYKq0KQULjFLjPmZ89pkvk3kPxz1WtI2mt
kzdcK0eoqOg5TFBF62ru9NGAXXuIc87Gk+orIcmY4H1E2/TUb6+yxofISjeNePNi
uknppt3hdSEWk34EWybscSbqAp1PQzqm0ULTNSOvwTzUEoY5SXPtSWuwF0blxAoa
KQrL+u/FCOUVPFrm+tWCgNDjqpRYYAkVUmaGcpCwl/SfZvYuRwwfJXQdzgeIiumv
8ddduH7OaSiNb5wwvW03DD7LsGt1ICMJTNOAmwh1sbWtstQYi2KBdPVI3bBPPSaq
lYpjh2xbmiRhylvLcespXvhIK9oUIqtFpShUoLAJ+rSVh5c7xMPtI85hj/C0mq1L
whta/Y//6fUF66bQBdpxyUh7UWDgCdgBAAS5G06p1rEv+5VT70WvAGX9Pr8doTgn
kW6eFrkDPfvK1Evyfcb+Tjj7UZ1rTXjfzcX6nyu9EJrNnzaxgYpjUR44VGreVuza
ZjODxw2pMCbeJucqmR8ojnZ0W78e2fguUOcNFwE7a4Xp/i8mud4REToV5Z36EpA4
Qtk9u1r/xGAFONKrhbWhOdMsHLBFmQZHprGKAU6NG+jhlVtEG7uP0GQyC7D5Yejz
tzVMG4fHsjdkTm/bB2E/VcTbdoPIgf550JOOcd8PbpYCxGb64Om02uF1PjaqPbTe
97kWcZVmMxXlmRXR0nrdRw6mH+UNchCRYAmBrYwqvC9SjftjobEIDEyHNEj9IRwO
B+Gxw9CtNNtVAzRIdHO3zDiZK69dv7U2x3GG1w+EQJjNSGYHCTqDB3fEjtloSJns
qbgQbLB938IH8YR6KRPH6KxdKbWkP3yuL0ho5q+HHJL4RUOfkFkupLXvTu2fhUDB
VFi/MYao6o/0A4XHDlJTFca1c8Bw1J8QFiXX8Z9zMJZOH12HVmDdwkV4PpCu42GH
uNDFPp7FaBoMi1at7sTIKOkPFuPxMGK5xnLOcEnm48mLzIlolzqOit/5AzE5YkEn
ZRpMnvExo7CwZ290c8PJgGdAsm0c8DPgW4l2cnFwDXsnW9qxDt8oVf02Y7AwUqvI
WBXAyHWMn8paObHjvy8hp0vPpH343EeK5pZMoQfCnFdLETJs/XNsvHDggIT1Ybbs
QZ7vWTPluccQQ9IBwAPG/7RMv2ck4YLeVoN7RO4UDEVrrZvNEdng9GQk2K8q+S9/
FQOxN62APKKzyWDy8fYdn/20QXQ4zGwpH2id4+EMNtbL40ZJtKow46MnudNI1ww+
/NqtTqqCE129B4ZrocuP/LKR9uYlC3xqi5I8UrUFmhumwIEIRgChADYmnVUixi88
ydM26O/tfG1JqB9rHxlt6PApH4407xzgt0t5LwDRaSa1sDw9wwfA0MUjs3X16s78
StbeG4cinyQFUu+Zs1MURjfc7sMJTWptHXowzM8FRp21RzVLGK0HDp/suazfVL6c
PWlE922tZu5mg4D2A/AxXfVMlINNVkALOz9Kb6K36LQXv8Yc1q4NDN3nTt9eQory
YXyPpJH3J1X6sYLisHJdHGxs+ZGik9uvGVXB4jFWqDaXiWC6tGeJzGwVJ4qf7mN6
nb+IXnrNES7uHuzSTeHwhlBwCbY2j4XiAgyBE5htvBohvHsk2igscKOg7BrL+RkE
qLFr2U/0FvFLelfIqhe+AbWzQ6GS2KlPZ3o1vLFWakhLMLllBvrbXnDKGipqyuzm
ykgF+rUlpxBP9ojn2G3LB5RTGAD30mbSIqFE15JW4SdfLa/Pt4bRJgIO73K3zN3J
du8MfvrbCPpykdNB0ntEPzAkd7Qw//p7X/f90oDa19UuSMBbG4l4aemnyPGYzhrC
lGlm58asU//a+oup/91R5/b+0m2tomGyB6kUZl9Nj4riad9YpL8ZF9qxrp5LcN8r
hmgbjxqmeNlTKIjfS5zCGFj3m/yviKjlPDTBQ2hBWHCNs8j8Y8X0BIgpOXt1JplO
KH6WsfQeXJByAOTj439smc9B7Lox0ouNC5Qb9RUSAhSidmyRreskLnZ+lwypywFl
CyEZkD7SfdmCufUR5Nk9oQxRF1tZpZqRmu6GZUmytlxFQeS1NDHaiKZSOu/WDF5w
an6dIwx0ZlgEKaAJ+/3cJgPsnrcCUbNh1xBK8HPsKcSKkOf+5xFslWjSwrWC1si7
aDj5z+v0HXefTcuk65/fRzgSGG4jXw1JNNRuot/Ohhb9qcrv+EDR8SMQeNBw5PTT
UImuv/1TvCNzvC8ARgFbh1d7Mu9zVdLfWlDHncRLd+pttUPlm16N9Ahr0AxJ1iX1
Mr7WLJsGwE5cFGAgZfpRV+RK2gdPHDINTH9uEKLSy/uYY5Q/yr80nHvjdYwP1LrQ
DdwttyPKlyOpLGgubqbypck3reLUvk5bIIWr4wBomg89bFGfBnMSz6bohUUuLzkT
+rgjPNwwCgI/gq1VSU3ZnyT0rBhmUUTpgosH2+gaIj+lUhKufuRJRLobvxquA3S8
/Ci6tniJU8mpr9BHNe4LO+/KoQoh0MK0Ayg2JtQjFdI/yPNK5BI/9nKdxOv8v99y
yVyeqzVSSYz4oCDfuy+OY6v9P1IH9NUNj2zx8ZNigZYAgqPWtAoai4gMdYHlOIEh
/mzytiAPaKaEjpygzrasVgk+q2CcOZ11S0eyGzaN5rvlda7pew68AHcx01F7gyxl
7tinUccExdHOnAex1OH2a29vtytNIUwGrZ+eJYkQrPskw/rYQx8VVGGEtcPgc/Ri
l0+tfrrCGViV/6t8RNqfOE4I9Is9GsI1+F7ayq/l8w5fIVP2C/9h1SJrE4uOasSI
ck6oWkfx2UpUFzCu+BOPXuORYNj35VBsF3uRz0nDWDo2D4cTRqBRwTGfvkZjZYoY
Cg1e2P08uxbg9IoF673kyQMJcKyVrPH2lQcUKhVxl6CvZkK2/2jzUlyeHagx6ZaS
eD/HXEvEw9hMGDFVYUO0Y5bTla7yiE3FYvf9lrW6R7+lOd2E/07pfa8KzbKqZG1E
DSMz9mdOwWYkfw05k6laZCCxO/A6+etMdkKFxiAq2k/WuD48QLhE7A2Lx8Eb9C1i
Y8/fCGQJZLIuFiR/usBTKW7UXQSsqc2n1mbcmJ4ulE3JCFSI0PDfu112CmgrAUlH
Sc/9FTRKul1W0IoWmKd6TijiQg75ZySdoFJq3CC+RBzTKKkBc4mudIX0te2wphlA
/7Otv7IbNTkTGNHhxUVqSRE67sW+LxxynngVhPAhm2QtMpWLbfJNSs04HuSork9c
ZwTY2zt8mMhyrIbDW695pI/2+MkoNs1mFEmfmXRKwLIfYBqcwHlLYnfWPvPTldzh
LcXl26zBD+HKLq221p8vdHE71jt16z1kVsVUgw550OIQeNlOt7ML4b4WvAG4Nf7x
MXuTAW6/XbbQMphvDqgE+RVxbV6NmMLGUkPJroqQ4DH3NSxcBO0LN4qiB+hqCl+5
SjgdenyzvuHKBWbKXjSoZCqcp3aEKT0B3GhR1pyGhewFCM0bMCwa2uEDs5fya1el
/4hNh/EI0oqUeA9utPfFuBvGynBJz8N/pOg7Qv7tf3wcRg9y2q8PD1Si7MgAUQB0
4wfoR4i8+JPs5ZOxd6sZapgN8FliEjT5hxefn04/vhUqB5qejYiUYeJBG2O5YCRR
+16DPRx+lRCmd8AQOjJz7gkexqvoZFiNDCGPzL6eVSuw2I5qJVoFolmLAPxAHTN1
fL7ekVHHKjb+y9xrAX5J1DSmZGq2D26DiF/JCz2wAq2FiduhF+Uk4iD3OFmkyYNn
gdgWFzEdw/+bQDWUfGOXnm4AthdfZEjGTDHgck+xvTWvPKPXHQCZPmZz0wRslSmC
uElsz4NKtaaydpo/1p+NpuQ+rQxEF3VvlGMQ/hZFHI7T6E7VQA8Ez1zgfO0OYDXg
8a4Wq+XukPc1AnLqllh5Z2tLvtbk400b9IdqTY8fEvtYvb+T6vua8m56XPEgPigM
VkN25FhfKjZB+1iseFRH5pgLI5HLqUmN186H1eMQiV/qn8M+uUVFj5ZfgnMlQBzL
p9LwS68G+G7Du0d19IrGjWbMrOK2uig8hxc9DfRIxuBXBW+nEgGBimDZ5Y7DPdRN
h+BKrKue5jxnHsKwKE2QiAmMK9rKE/+pHJWi/szfuUeS627J2LMY9leWBUHJFf1f
59jRM0lUQqkLvEmLfq1YApK+xHPDOED5/yrzKf2eqOJL0NgC6GntZfMsML0vhpRC
3czLsAm+SFRVNcfgaWjKEs5+m++44+4hPrwwoDO+VkIDQf9iWT87pMCoixc2UaBU
E3FUOw+vP1rHZwfp96hvs7rxt9TO3tOdeJCXegDaufTu3CJ12G6VbrZ/AfTjS02y
8i3QHikQ7R9GHfr11f1HwA2BQ2wcXxDh6SkGNirUL7I6UWDH+Pu9bsN1YBATtVwm
sTdGlw0JqcLhzevHSYtm+iL8HqHECsx0VhJ6dE8MAGb9RcNWqPyVA1S4niCnexXo
IZhq7XBrgkBNN6XpK8CmAt7pYtitffIPLo+iJ/jrKQL/x33Sd1GZsDq86kotlD9B
GboCfEi0ESib6FSULQNoTzTlRmF6UBK0ICyf3ksDTGCrvNKVb8W1Vqltm+EUs/PY
+X51JQ162t+wCkxBNbl6fQQ0BXDx463FrtAlnX6kXfkCDdVcNgBKAT/ov4y2Z+nZ
GL4EhFqkTjzMNtXAe9zT9TUoFE077PEV14qPv28i040qNFCX+n+lkmiz4MSE1CGf
mwCUeQQZFOWYii3n5aOOoE2h6R4xKv313iF7wZbsf+QDfeWkVQfXTpHYtWFhZjgX
GKNHZZ04pzMK/i8JWwiHiENtk6qbcXP+C4KaupPrSZPr/AIeICYjTqqFJoCDC+06
3VAImbasgGDWbyf1jYxB+xJEAt5FpVoUMovwHwuMEwN9TX5S7S8M8nA4ASzR8FsZ
Q+xXhvB68a/fKJfgUwx8HyfnnbbimUUA7HUabFjOThXSywwnxi10BfXfa7rt1VFE
q2Jb44efFO1XMlSMYsrfYAZbkMuJxorCBidhVtMjmLqrROSqnsPJQkTLt8W67b+y
CThHm//2omdcnkCUjqOJpaMACvFuR9E+0rofbWwPTGA+szYTLkEyLZLCHZqRZblC
BB2na28wDuga6UX0cU7AUXAErACxrzVwq91/sFVLiicGcRXSlFIJ4pM7qEzomzOo
rp1EL0YuXQIOu/EpfhLS7YfAMksqPzhGvX9RIvARwpDpNE84n6gptd8EIaf2BGoL
Fr+a17n+7nTCdwgv1NbwXH2oloJO+FORA3kCe2qHkvNBYNZYX25Q5Tz0iyHp0VYr
F3l7j/aAQY2j6E+6IDOBbCJQBolUZOTpsg35wWUbHmxI2nq16oyPRVhK4Y+IM7HB
jqkR25IrOzxVGOvR9gc7M9BYdmJQbG/UbwXq4jh4Tib7e6gqLlZ98DL4LoTz5c2O
y2sRVmITYbixvQ45OspnGNQQ3nesUcf3eU160urdKbASo6MjoKEPWAIv9yr4lNbC
EccWoG9gT4m1ca5ehF/bQ0scg7Tr6Vk1op5Bokau4msaZCBGt0lb5NKfCGGZDDm9
UPgC2rwOhs0YPqzIP32Aqhk5f98jNnkYgAkdGdacL5kUYKYSEnxhdbMMQp1qHkEs
7eysAvDxceOhKn2E81v+dY6ZVPqq0YydGOUhB1xfTBq+JmPj4TE4DQc1/oMusatV
XioFgTKcttAwZsJblcc0Yijy/qwYJShpSD0m2EN7DfmYOqPlRK6lsjSQB5ciR/29
cxz0fqHJxL9CLFhyP1fnx3qhp5zltLbMeUL11Pw6pLdmn/Wc8+/pY8xuGlv/ObGm
lYDCTwkYxdlHUI1dfDZE7i35bKShFVfly9zl9rHCGpvZ2Y38EtP3Aidkk4rU710U
obzSI3pqtzSSmIH3vK6/80buVVt4doXbqJFuK4RP71JAhgiWR6xxPAX2dwl3kkfd
D7rtuKjSKG0tOUNdXCmBfhhHpX+kH5lDK9S6MTV7KCfnD2mFqSiI7CpkcdVXKJwv
k+RKKl2Mva+1COO6dZXvaWK7WCplPd6p9pRBK+lYO28dC59eXYbesQixPtHrrSqp
GwbBUClme3n3vIgC5dRqJnE7u0B7vLNL67eHydeEq6DOjE0uw4WdsBO/NLE+NRrU
f5mApMo+2WOShL67Q3McGQ1NSb2y7pSGyvt6EK6frRTohuR16iDbvy2jhzLBpqIY
fcPpiBLi3xGwiI92y3wrARoQJe3TCfUyQl12ehv5DlTrMkgCxgkjKwCqB0pewaEd
mOgzx3f9oFi3TGX0BYZMhy9tbQvnR/8Id4wUg7n/O1NQaqF5qtnWhQ9mpJ2HAnFQ
NmgAUktFc4eLjIFhmA45yzg9H1d/PznMx9UscT62nONt4qmRAdUkntaCF+OymTpm
uxsymaJ+Oxjqn5UiTi6MSdzSoMRMMtUzDc076fj8C6nM5uqh8fKR7qUovgOX2hdG
LOrLZfStL60phO8ttp+5vlg5PZvkQ/DW7wZ7kVKwCnbG135eUkmPYivInLvzOMgg
YEkMruzgTxX5dcRpXpRn+bayILk0KRC7ekw+0z7Pa1SSGOSvU5VE7pPqUOUJL8eg
dlVcXMQwiOBs0WR8hWxKRe8lpHyOPhTNJ/bcihzOvXiFIT5657AtD1iprNr8zeIF
HKYqQ+H6IrcGH+7LgXFmmnpnM8gR3EQn9RFbxgaYaRur5ERIRBFh5GQ3ZoGS6B92
j9hp/icv0vGI9Bcv0l4u4y0UMX78PBWFuqd23Fdw3/JSN0p0VGqlYnixDRP07CTr
3UVUyTvOPLk/bcWPotUBvzhizZ04jxUsg9kY9lxjrQgPrxDw8e27oFk7VdcxrRpB
EFYJnHOUNPBOgvXHaQPkWbUjYGPR+K3VkXfnfuxCoU2lLwZMmVa8wrsREIpYDwnG
FUGv+RrKZBhh/rWkA8cGDVrRM8lbj9cq4jCRJvHzgmFPqAHuGsBTZx2KJaAKsEhp
NsEecWzqHl58Pr1jLboYcHwGdVDrcMN2AmRS2cbFmDvxXC7XXsSqVcxOhlmwAZ/7
6aRScVnZvsp7uIApYYp1LP4HoDRRzLg59+HFrOtFaIDQ0j+stb9wKKhd3VW6e4XA
L4+WXxDjM0Drk7tw9SzCvmdU75o5LrJG/bhUiJiRjQgrF0o1pxmO76ID205zD9bQ
8kYQ0TtvMEHH0o9m3SDdh9X4reg4alm/FhXNMpwvTVGbvbNtwDt2rxANR5FDktYl
djFgwl06i2c4uDYapJ5n98LBjAM5eTLjaB6QFMTiDrDXjpiZoeTUbMFe9bBZ7u+o
xJ5zcYPATW1wIGfYkCY/CYiJUnjoGwIKnNUbrSB6R9qBuGjn8tU9zGg/wTYeQIj4
UatxdA3MTgQ/uerU4vScCjhIifCXyj40JVZspBKC7mq1Ov31VNe2e59qKjP/vlCr
VcukPxGlZvob74dPgmy/JBMPmotgXr2c1J0Xpj/kfuMpP8VjFl2/43bW9AeNftLx
qezfAloTgd6nucwhg6avHHl9/rtfKtPaCSA9JcvtQFHAOTy7ufuvh14rsucAPtPW
sDnqIw1cfEO3wR3kbSqaHCr2eA9e5bbxZzf3RbHv2gMMK6er2JM1n+MvWFAILesB
oFWozSs6ORElncHOjYrrbqqFcg+uGO1dr0Uexevg+O8u4RAgqR85v1DZKSZAKSWl
NPF+ZYBy/SMejcWATeWkW6Axq2VooH64VRSpuA98YDzy4SKnRKgAMejjj1nzO8kc
1aZ31eyNzqoBxs5hrMvtl2Umo0lTI+5HTMzAV8bQUJhRvmWnTfdpWNRSX6cyaAfw
j6QzOvnmcP/ku0lqOOX1Ezg3EpQFJXi9BUnVeGk9PqCCeGDYtMix4Hr+2xcCHkif
YzRU51ToAXF6KnN5l9Qult+Bx6yu40AGDwlsxzP8EWLGpI8KS1JlBJ8nt9sGTNk8
WHE1IfJ7vHE+3rBO6An8jOvY/lLE7K6cm4MY9e8qBaNU00NM4Z7yN1O14HmuHkAp
rnBcWbTHBCm4MGceuOXZV2AX4bXu3r96remod/36pAP2WktQL8HGGKsyvfVUtF0y
rP9hGoixzWKeOscooa0IWVgPEknolLDJ1wveJxb7i8oLDSGeKFcVyNYFp3nSCKlA
WOJCz9dD0zjtWjpnOlsuNN/pEyxrqkdDZin1Kf+nhkAMJ2KSn1uTgRamzMiGMnlY
BBJsY46EOXdGaZ9iUdyvvF8JNx1//+6rUtPe1UZCwZYLBq/ft0XZLFG1KlwwE1Zt
uImcKWRnVvG9kO3SRyNoE9ydyjyKPAXh5mAfvKRafQEFN2VxJPnuelBf3IP9W960
fKcXSh1JTueML4wlubhLFZfezQPUmBMer/7eUIfJNH2cYsUM5re8hiKau+E8P2xo
4VpSWynBvOgsSNtPKM8Ckvs/Ts4m/aTO7Wmg9S+/fjtKvhrJKY+h5hQlBgnRmPz/
5EssyIWaoRzGw9sjsFiC1Bz1JVZYo68WJ88GoB1MA5ejn/yZZao7f/3tSXMZAg/d
LoMtkNu4cYWdaEQIrEnszqRemfu3GCo58sJhVoScJ88K+6gAebrUoG1e1VFTpY8G
R1kWpVtK3mQYe5lXHpL+TaG66pVs+2P1qDlaAHGk5f9nNFHl38YOW2XCbVhehzXm
pPon8fcMKmFPtbO4Jt/TXCDvT3zdMdPEBt4h51q8qDFEwvt0b9gQLds8cfkFn/by
m85SolsI/dJOMqQGI5vZOmYWXIuuGDz/SUJ7ULaOibjRNmT1hCoivEK1MsU2QQXH
EgDkKLlA025RGWPY1EtR5zakQV+MotuURRL0pTYyVVoO4sCWjZqEQb9qOySgUXIU
OsWuyJ06FJx5zrP/AjfxpG2Xbja9/SUHhP+qKfRjMjSWuoMm9KVhHP9Xs6xXy9aS
4xwIY7SjNAmFz7kxB05JbZIKmDj3YLJCEc/5KUTkEtLQkDZCRxX+N6EGCRaivQIn
qonMuVGwK3hwIF40UNdWf7NQpGCnbM8IlNQ9tT5tpdojhHTHp/4Bh+qlx6cUabyK
gDss1a5XulJIVLYSGBZlIVk21hgIwVJKq8lS4YedQAk2KVg0xaPVVTfNYGSiZYui
5pssUI+SvVc9DQZYbm/ve+fBwKTRUsCkgRckaUycJWgXHh/Ie2gCf7SKOr/JNgQh
ALj0Q1uI35KFgK7zexEH+N/0JfadzORfIDbk26AReTIy3j/q2eyuWJbCX+SHXu3m
WuYE5PoLoOKDrIBQP7nqq/mHT1lQyibgra+NWYFusnTul7/3G/z2cpNILCVSWTY3
C0WFEhCuT7qiYT/OvDxQjCKAHeuFwXNpCz8XJYTGmfIgk0FrPSpSTCDotArwiZTO
MTRljdDKUdypbzP/jq8eSKYLrAY9BUy+ClqZDJ3NxBhlio7peec/zP/WHYVSt5np
zWD6TM7QNp1FDuPPK4xaFu+EOuLAUTfPHa645xH5NsoFCJ+X6UQDldyn+DFEIwpS
NljO8kNKwMZLnTuhxFp1upxduAVxMnRN9YQ10b6uRxrtEkuZcbREh5DOOmt3i1U6
Lz6xvcni5qGVGK7B4lydb1WXyYeviP+2BxSfFEZVse6qRVP/cJYUatv3flFsGJra
gCI1LklQySNHVZrxGjsslR6B9Cecghb7zS0X01/0XsRr8M/ja3khGIaFWr9WnE1P
r1b8IZSrddVQoTq8F3uuydngmh2UOIRVUjg0nILRCX5jevmoAspZZnTqRYydUsfj
YvXJkR9U667s6dLjzTsEpU3Brtdi+3IB7237menQ9GthiatpR3IdvN6NZxrCbNzl
pWHiqFdE28deGnMpuYLwK+Cyoyp8mMB+N3ycBfaQwHuJfHwfU8SDCdAb0DDDVqET
tjcaVdka8CnkAUuvGiezyFBmrAnfieH5sPXUiLtp4jDShfMPsd4KbRSqa/OX0vzT
59Qs2P0UDTAeippzm5anYtqBUx25DAhvwzt3N5HngSimd7z+4LWh8p45BmvNJn98
WHgbs8Q8Kpk3M72dYhvq/jLhTcKWFj+qnaT1uD1lDX6mn6ufAp8CcHJd/oUbnMwF
IiJLm3E6USaAQ0jvULu90KBhsXZZ6RceShJRQmlU6fA16vc0HgUVv8GVwziuoTna
B6EPF+abrYalMkX6sXFSzAyxpKWvsFJYDjJuci8bTSv8aWr4BdSEwkRiLobPRSqX
0WfiEY8QWWIQuLb2BhoZoeliWmS8oFFgTP74DLyCfoczAyG44ihRWjXY7fe7FWDI
qY1v8bH92jZn3D0+48RvVJiiH3PHgSm0bakTcAxAeav/J96XVQsfZB19LOishKXm
br1SPKz4F6doEI2WmopHmNzc2PgLo/k+l7MjeM+itGqjeiq7rhUhly5JbrQq9mdE
8wlA7cn04bdLE87fou2eZsBLwWm/Q8w7vKB9F8/OPeaYJF7A2Vu3BhE95uNgqc9M
BochE/zCRiXyv+QXtBfQRQ+1xlHKB9z6dV5TjwJXvSAFRViavZIah7yX3fVv2mnS
RVfPkszfp8rRF7VmVurapWGcLhQCPwUE2QudB72b099zXWU7m7w52GeCFYqloBL6
D9YPC+R5UIuhCzce6ntIrZoIzCKUjQlpKNHs1rdb8fk1VFsSUkpUGJ9Y6jO3jpfP
TBuJt6dIcx/NLh/yQKcBDzB6DzxZ9YZ10I4rD4S3qZwWu9zt2nS77zeu/jqdGM9O
ZAO9Z7U6lTiWcncAv9lfFA/gu1WbaQWRzn0o8yDgUaw1diwljIwqLBGoNTTVpz71
atBStfz3u4qfOrI46j0AGFSpjqpDuOp0LS1DM5gbwe4udjpJ5w+mdVXe0TLfn7+8
h54+SGnOKEBsEg4O+GcPFKVW+6qba4d6K4Fes6j5uBpHJGeQX2XwRceWQu9HbUpE
4HBOLuVqCpSzYimQTCe0wIFurkU3ywHHe1ujRmF9QNYNC8Tp/wWUM06XUgwFF7xD
q5B37NjiIcG/EXc4f6daT9r8mWNWkcr48m8iCfkZR9x/dGa47RkvHKHX2b8f8nin
JC0qtGUKtEYAuGsVLakA6LjISK1UOdttScLAbuODqG6qp6GV4mo9ePtJVkUDq4hC
6SE22ZIqP9NsU+wp/WEAYlhhFVsoaONNJJgjI/tW6HuMecYwnUBAAY8K3xJF2YaG
zei+1xdFOdKlLV1RDpkuSWRmQ+TeN+EaOlEWGUm79AhLFrYj5+aZ6hys2Luy+Fpb
ySpAZJLJXSr4l3YKYpYkUYeLAQ4HkV/Oa5ot8y+nYy/w9cq95kBpUPCkBFV37/aW
OO2nzUByRLDPBlrcEdcd4koxj29xgUhdCrz969KlaPSY6CIOF6tzZZeqKjvIB+/L
ZxJ2MD+OXRdlH1Sr74TEptyc3Cmc3tKWUYPo/ss6Wfa3m1oW3APaAY2n0xXz7jX4
hSOorJwbG8fqbojNuwo+pOz6/gAngWQbRU+kq3ATvG0N5AZcBZ9RGNVPE2mBu/hP
mHVc0I07BcF9iFuXCgF57d7E3NK41GcUnqQ7CegVuZIZegwdvnukb7AuVTE++For
d3/tUm173t23L5S2r5gzo06+jysg5PO/gZVXvmD75M7sY1YFLjTEQkOAs+ck7jxt
tgmeVuTbM6JycuWf4ZaPCBjj9LEoEGg2UrDmj1cvcEw2m2wYMRZdqeP0lQGOXuFi
VF+7VRaAzUbYJ2xn9YOQDKMvXvk7nxggH/gcmS2Fa22/1cI9PBSAJxfohvgZou12
ifsTnZsDDhV164cXXnxCfkB01WCjrx9D1oN46FSp3GBbNyFHRkydUcQoVbhjBeh7
yXrSoTAT+FeCswkWeGwAA1q7m8dVEqX351cxRIqlAU1TsCxTfyk210dxKCdBlbuZ
nXRXl7kHl3gVkihCRdYQV31HNLeF4yJMoxjceXxlGzdNT+MvBQoqsoW/2XqAwIXs
FpCHfp4oZa7Wu7ViMdruQ9O9QHGJJMV1SoMm+pO1C2HwKxIS3ExfmksxxbNIki/1
OMJRfSxZnOpHb8+GIQI1nrSsINogENtDRUhKlIdYWjeAnF7onM2mh+w019EL3NWC
wGS7KB6W5bJsiI8M8oOiFAeeVSmsIfNT1SC0pDS0jil4blIisEJwVrHEhKVZBds7
BpxnWEQBpnQzq4tn0HVzrVMorrNzFkKHGLIaruGPYIql1V66LOQcHy2JOniozrFD
Q/Mh2NSbGEJjkkolmxO2e1Z15gM/OajRQ4KLcciqZ5HgsX/pqmkNom77DCAIqs0h
PJ/+y+liHYvt0YD3HukgnQZvF3zAhdUvMh+A4WBNvOdIDfZm3xX/wLdghN5NOC/i
S9/sTPnqzXCI+PegavbUx7bu0QSQY5Y+P6D/qyVEsQruRpYaw9lGnc3u5sozsZWG
/a7MRIrdYvi0BSIvTeOZBQ5IJZGaOr5f1KyHpkbaCE+VFKpzMoG0WaexWop9XC1Z
wBW/jfLEPS5MrAu9Paiw1pT3jITODE3CZvVWVEuAFf7M/UPn6wYS6821poIDDcbL
4sl0kD0kc0aNLoYghr85/3XmV5zICWPK4/i91kVJkU48is8KUF+Hu9H/VeYgMyZG
+sNyZKbpyOKIxJEDnjS13LtcELu5Oy78YQ8/+fmVs93hFKKeujhRpx6AbwYxJmfK
Cv/tzeVtItfaFuZpa3m5ml3yojC1wMlT/5j3W3A33Az8n/ZRwWaMshzjFde7+fEN
s/dB9N/quArqzG90rdvb6YWw5ZMBP7eMk6zA5a0eMLVrHnCV4YlXtzLqwWQ4YwP+
UG1ztGT8kIw4z3xr91FtpQtOqHegEe1+ffbCLCtjn/dhIBcWEa+1gSSoLJAssaT3
76FTt/F+xs0Q6LrPH6k/0gCBJEvRFoWJUA4Wesd3R0zh4PhYCOmqZzwPxLkT9fI2
Sut7s1LkHvxx9KOUWf92hpimZMAb/HhbCwz7+9Tc5Mbouh/BWEKmTPwQpcJu4tpi
cqfrPqb3UQS/dfzQC+Y1B5v/DeNh9jAVdkMTOVyozBCbK149pmqTCsLLnVX3Hyoq
XIyvxag8H+E6jFWPgcNZ4yEYjn8VnnSCHvJAMFi5/HbjV/qeDhgz+5dvx/Ncch7/
qhLBfidRu9FQDKoGyIK4HubEEEVVremPjc3TxQZCh07KICLadAxI45PVLQ6PqBMp
qwfylrYWailPS0nt+CLbl7pZ3QWXuDystM5re6zf9asr1QOc/tHsBrOgVoQnqUqR
prDzYluSA/pDu4+BFma3DMvqvRAx8FI3DYjgF++UQq3bjE+k+7OvCCteMkgdFJ1i
kabDNRKv5hbbNTEIdmU9lruTPvwaKks3k8fMeCsd23tRzdS/Suu6cokB2ANc5HGo
QJkA6nancTbhf8ksv11tcjTu4IOx2O/Ua1mIdYlRx/6WK8DekSny3HKLIRSLapxJ
zSyfWJeqXw0aqzUlYPy7rYuWniDgA4yFAjRIwlTaYsBNogbQ/xnJPidACKSJ/o9H
qibY1jvqDN6PAoOiFXovEgztiopqyFlxPd8vTMBRF/UlwxyCD+QxmiAw7gXMhNqk
2ZeZWmo3Fe3/PMxVzpgDmB0b3QFVXnzga7vKSYK3P86MJ1/brDXVcUuwAK1rS9ln
7H/zipIFEhZ01dRcSFpvsA0u5v/LbD8rCwq0eVZsSFFQqyoEAuTZZOAINMmrpPHm
43NZo7wbjajXTglripQ4Z7BFMQe8hLVuU7EtgDqRcVpB22z1t1JstjgP7ogUJ6EC
00wfAha3ozPPyEvH3TT5boGuS7+sKtGggvM5c7lu7ViGQGt39kyeem58RBmCuu6A
uI8GEW5mweH4s6wmjPAAYj4OfNCnl4Okhp9JtLOAtIk/L685flYCFuO95mCzr8Ur
iNrZf2a0Mj9DUF5CFG5UE0hDix2mc57n5KzNI0z/vIMUZBN4vkml4GJjCf72EFgi
LcDB8ZeqlQ8tlyVpKfV2bGDGxKPvJm6mKTKSrCHD0cNW7RFuEULZVqqqRdrWWBsO
g5hghQ3XfaZJ9IKjUFyuLQCF4+SPvV7KGm2M6xdaobC44tCJECcJovBAV6OCbk3G
DnCaGgToOaSXynr4WGkSem1AnuW5fXuprcZFtBNUpDeZzLIJrf39TxJjsrCst7Br
sl0fVBaoWC/qm8vCGnENK4D7sZlCXVHYM+yHevyDwpEbNSCVnxF9o9cCtmi6BdZQ
oOlUY/Fi9yq+7qPmS2QffMboduJ3tZQknwZn0zUryJhLT//UbKjC+by5JXeTwXEo
xN+mN7+IAN0SI3Yhve4zP79nUkzuO1VKmhXnibr13lG9JzR/r1TA49tmGwScp7Ab
08Pzcq1Nf2hrmGJudjwvnjeV9SpK+24vcbBFzB3d17z1ffZD8J+FcAYWk/iiQRHd
zpyEXc0NRkVjfyxAFIUlSjU/BnGIhCXrgcIAd3ehgAJEnE3pZo4EOUEKoEeCrV6b
TZjm+hO+7X1mZwDUEGC7fNTAqbYpOOs8yR9HwjpviUUrOxc0UJnbBVPnh6bUoayQ
nI1YKjlf+XCSoQ/wNuk8VlJH7o+rlGmdLHuF8WcQYEBnZvsdWcQSsSfkvuDrOZnf
MpuFOmsnIV0Ej1R66QX1WwDRPzrtdOUMfrWvfXYcU3DjvhstPGPYZpp4ivh2Iei4
WLw2EZ+0thi9L+dOIx9O4f3wJPbCFxoqdA/WkYSoNOuxfsAdmiVmx+XizWk3EaFL
FVFPfmKx9W3p2tEx4fpGpkhzZU5zmu+UBgH9O0kGm1qbwzhy2UbHHBjznqtlAlK5
G8VMAA0JTC8thoPPDb6IGtzhq3CfLFOGYQFkF6NCuXQ/Ac6DdIzfKpPQQtkrKVlN
EQCX89j//ceqQGYYYyUnI3k2EIMn6ZMrhxwJYykI+F/yl7FX8TbRpBnxxTNvWdbN
oU1g8+Vm9zkhl/23wizUI679DWC7zasjD20KCSCbTOKvDoqAczZAkF6JCsp8J+bn
tt5hEm+VUhDTERGv+GnqzImlV351FNX+IZbxMp8snT6wTGt/yzuLNY5kNrpEMimG
nTtqW+RMLLA0PzplidUAIrj3PSncX26z6qLQQYlwRzDxVT23QBSN88dqrIrvrmjm
WtksfjjHLna+XPkTektIIk6QSpT17Z/Pm3dv/61GO5MMxFlPzv0e2bs6cs8IkpqF
JEqlW8KnyAqZ9nLDhR//VGJ9u3RtsBY+PIfLDPPujXs2WyOQdk/o30ly6mjkub9s
vQOp5He/jrZYi3ljmrhtLNvULqifAARsRFMxq+TcrLRDY3YN4UHVJ3/uusjdkLr3
LRVEqd3M+3GHCSHbIZfXuZYRjCWTjP3ETDiIPoMpYAxhW+/x/jpI5UtZ/r4iSDXy
sa8Nbvt7/3YxThtV9o18lFXpFK2DKQyD/aGJfi1iw9BAS39fw4QclDxIvfdL0n11
/2G9xqjWVvOy+HblN/b74AdI6kyo+1cXjrqwHW3Gwrkk4y08UUv/9XIc1XdC3wFT
vl550JPVzAMEoevxRAbXt96tlsCqIlRBUaM/AnGzctUZN+mcwTORzbfhvuZg1CqM
zQU9qHgUDgvjRLXqGsFehc22KHKXgHp33RFBkzHOWHYQxryOFnD9nyaXdW7FVeAH
hdeq2Pd3etQ9dD8KPS6qhjATdP/CNJwBISd8H/efGhbDdLl0XurH5gCYPcV5n+x5
bxfNPQyyUNJniF9DL9opGi6heg+G4zwKqoH93pCEeF9gfjgkD8KCKeY3smBAWBd4
M23nIwx2RogllbTRRdh1LEKb8M3W+xIEdJQZJ1t0TOE7xlsISK842dNZ0thUv9hM
hTyRX+r7gVuqeiIR3UHsA10/J3Moxeo4JYd3G6lnuESYVRqrIUVrUxTgatk7nCVj
5t3wkQxd3nIZVMUbExsPRgQ/IkKoUzfsWa8GHDX4TrKrdT3NK0K2w6C0ZnGkzCCS
3DruFjmhSsNjU8/68SYBTLbBEs+Nfj5sXI+6WdhjlutU6PD6LEfXn5EnNimpQ3pt
Zl1990d4e+LBDVfSx3DqUiSj71n5bTPbLgb8e4aoQHsH+2T3cGZefsuCAErOb3fk
cMX47OHPaGrY5r99tONiGddAnoYF+W+vYld/mtTMJX28OdJfSYXSt4vyaZQLfJI0
ekO2wxCq8nwN1u2Uy357dxC0R6UYlw+LNbF+1RHnHrGwMXFogAhaUe7IXbbgv88U
HF5/reuxOZMAIvCJ2nFqgbTyZdFeSCtf1TppHv1Uuf83VzyX3FyxVWb0yAuv0bQ3
3FuuH18fDQj/EZzLYOGbvwQ3vkQ+XCnx4pYfGVYBLt0tRAkEXOyAImZ1yNb2ooxK
sMZ87OJ1vO+U9dBOqnGg4prqRlJloWu3sriZok7B4o1wsiQmtPlTw/pNlOTFZDW1
+yxuRUPoA9NVxCpIoSlL1qRBp0tAQ4uI+VamphGHBIG7JRP5Ijc65sArcRVhbzgv
LZee0SvvW65cFhe3L5GbpToTtHyhTItaIbN7YUbJ9ZZ+iNkuzKJhNtqfUldFPhFZ
4xLExyE2j5bPA38vWLW1pwVHaM53QjsNgJwhfoxXiZOXTr8FQSQcnPxEWj962+PA
Q/QnfLjojzeyjEWLt278EGOu4TZdKgbQSMfDbAcbx2xkwydpjU+oWj/1Tk5gGlyO
Mt4VEy699XUvIFOdvdnRSo52Fmsxjw4d78DVg5oIZML4/QFjax80sFT/oq9+kb/T
qyvoWl2/pwygc+4B2JO9P58MxVeKSIWdhv3qCDSzRPQ7kodcwvY1ZN2ozhl9qw91
9znSjiWLb/3ckCXmZq3IKQT+2m+F+9960I8cZFJHTZDveIzsIlEE6X9BZlPT0iRE
84b633wknKBDmt52aiBEXHnXEX99LWnCTW70ITeyoDCAqnXueuvXKPlQGBe0D3nG
Hx6bKr9OGyXUi8YDFCCVXYTdI4GXFuEzhTCxeol2Put1ja8ibZjBWVC8thFc2h9/
h3nd5o3XQdKZ2xFXtK0mgAGXEgy6+MpBe+aG/liujkFb0SC2s/S8vlZYG6IQbkZ3
pdh2gOT7jFNiKgfgu3hBhHYqTjlsK41SDnE+1LHaFjUElPzXJIZOLpL0LZXFvmUy
IqFrS/7MUl6MXEjSPLQbJf1Wg7tALksDFbi5gwILpnuscRAcHaCZswCDNVhWhGZi
E2Cn+Q0Cuow++OOor2VAXy652UC/ejs2jQ6jqITZI/i2FsuREI04BLXO99nNApmR
PEe1hmrOP5t3ZqQMMv13a+rCE2MWJpfVfzLIqeKNCU4TnAsdZdeD2Uz1VviB82+w
Kj3npkX4CZ3+LNqmafPBL26kJJz+QMDY+KD9bcjv6yC8kCy14dPlibtkffbolNk4
0UhrR9O3jR4RhalspuvwHagKNXfi9+L0VL9xcNUGVjWLxwBPoNUwTbS+RaCRmC+A
TfjSfq0c5ofI63pBTSXMOQ/QK399alkcuCvWxXpLpgWQhdac/T6ZnLYP77xi20Be
jNBCHR7vvDBh+7SIvh9MedpBzyi6lDcNCdJAUZFsJ9hrXBZfLkArU09+yxjh7thC
M2pr7t5YdRGNLcPP8nDwUvyMn+nra25Fkabby80a/RL97snmNq+xkHCOA6FC5j7s
D+kJwsiOEv6oWQrKkX9kWMdEOq27dv98g19YmylKU4R7dEid8gmZLncr9ZFyoJW1
jmRtZnpMBZjFcY5iFV0UwpsP/JEqv6tp/hZRRM4bgclb7VON5vaUmncNuA0rhOx7
+l4/3SFbsHshwaF6OR4Bhz8HkQW+EN+9xgDpalIRgT6Tglp9H9noWo7OVQEtYGsO
Aj7fTBggc1W5D4SjO/J3gQrWXzCgJam2Fc8Fi1ilVrIg0qMeQIKm8pCYzUipYbM7
Nd+1KOeunmhp5D1v/eCLX7Sd6cNkLi26cs31Y9Qf7JVOwOvkO8F/f914Q7ORN0gO
4FgxYHHALbqS9xsWg6O+Y3tvW2sSSFfxvv95svFiCE/SkFclyRlTCdqyq2pmQtqg
Lkjfc/vLrXk63REEYTX3P2c9kJiJ/XHTntp0+ZEaAJVWULnpCiUXat92zIP611+z
T4mO1Abgi+FMc/Bs5BJHbTZdsJaD7SLof+yKZonG0AUtDiWStciA09BgPqEfLM6G
jyeDcjS2ueom+57C09Tvgy4iC7BPBd8FNNhFnOjisJ+ntPpgPCKucpB2BwyORath
IQsUHnqzX6+h2WkSefNOTnoXHlTjmSa8pN8qbthzh0lmwsPHy+vGWgibjkCCXuUa
aUraEeBnmIBhqMtD25HYtLVX04NQ+Ng5zd9xPDaLuAl3+mD1IuL3vDNR+5RCIBhA
yMAtnD8CUkYHM1F8JdpBizlVKFvtAgHjpCq7uSxuihdzECVBzu8VV3VMVH/Rf9PH
8rBc6M/lbjQ1GFIk6JO0XfWqXZVysVbkSO71ECvpwj9A1QBdvA+BTkh02YZizx8G
PAExkKas9lX1I6QEltgRsCMhD+1XWb9ZwaqU5HqgVWNCGA/N3lNW3OYihrNOFdE3
BaUTeLqLUnenQ9ulo2EkzGwlSnU1ZeAThPDoUbGxnyjKUimCN+5B+q2m7OaAqcyj
mHfdyJxhuhFqIpuNbe5AdKxxyr6maaw/+Kg8d8KjRm3rx8KAt/qtsM3oMub0vYIn
SZdQqD3BCTpeG4v1FGYCyKsN6aHf1/5aJCMo3sRk3S1TdjfgGXUyBb4pe/8SyzWp
FYRE0tOSjyxPn/MUvMYoBpMV81zKO2QqAsrcQEKV5AlCayAmeibxA8jFQFb8QoVI
ZEub8v70Dr3nicroZMrMMJ6mE0vrTn+SNLU8SzX+uRYSdLaXSxK+5XH3C4EainMS
Qv63Vte5GF52FCqYn+tUmI6B6wkYuuT0iOIcrP6ujwsvPfQC0O5q9giVnnwPl9Mf
uzcEu++rtqNRHV7audLTPTyqOOqe4zTnoi4SYk5VYwh8khz8OOh8gzdJNFBE54PL
bOiQRQq/0/rbMKRxJA+4s8aA5NvzG88yPeJ6RnkATcLXSYx29fX6DF2xkA32t3WH
oONPmoL+Fnvm8Vj092yfRvRrmWmjkw4/hypC9aaT4LiDxY8CtHeT+Ja1HEA3WLDX
TEnc6yDumL7HEvn8jQlYxvBteSWLX17aE5kcuFp+eH6IDqdInxzu7aCMDPcNQobC
NxUkJckAF/uifXtBkkiqVDI81RhoZnAqHtkE9W+BZiB8gBsy9zEnYyjZssYjT37T
hsDWzuRmFY8ulshnUDSdHkRu3QutGQMY2eePDQm+sFRbSfKGrJ3ZCqjrBTffPXnW
QixDwaEfqTGA835RGQkYcPAXlyThIB08yWSUIqolz8F+sg9C7DLyZCs4BhBBpRbP
659b5uWfEEWNS8e7N+MZXUN/QaOUX8Zx3DCXbqtdylpH4FAL7slXouLsrV0joUCe
MszhhfPyL5mIKzCQ/8SxPDnRIlgYmoxirwQENJYQidBop1k9TLTegTmTzxkRsZlw
BaErSXQuIIkGCEi0qm2Svqtfy+/O2u2FDVZQF5qbvvOrgMEAw5KnBMp7x208LrQx
qV7sXFCrsf5Jrd0Rrp3M30giY0C6dbq+A5z8sR1/A2vWaC25WwHNZJo6aQHOdh2b
VmhO2YMr9J0t/3orXejlESYz2pjAtC6uykVM4y62ath+wJMmtUP2muSjl8Ul0QTU
j/KM+3mbmuSc8Q3IlPUZmbhuIPazbTRypi9Tj68hMb/9z2vglfOUb0kqP+mP9q9U
gzVXizWquTrwXZrnMSR3Yzzi4UlLlUh6PPNOrjBqonMepWTmG1knVR1rD6EDtkfT
JzyJsE+n4yWw48iAZMYBx2IpPek5V5JfFamFoWyktR4hMAcHKDeYUbLZzLQCxUu8
Z/EjlpdOOCjs6hoimKd1QGr+ngwQJBdgVg56fPQMp7ymxp2tYtduwpKsbalhbvR8
OPD7oCnDjvVvDe8OFqE3IyQ6c0N8/hW8ee9zS3aIGNOSvMOJzlofQPvXu+aV7CG0
aF36Z54wa9E6rk7A4Z0+Pba73tdWbGGUP6SDLPBsCUI/mk+6h9YfkvvbLM+YmTy7
rMRk2GrEdNe+FIpqj2fgOYGMtbVaId8C+SVxuXCBLIVHf35YaPPMUoPXcEv0sm3m
OzfCu41Pj06g3xG9YFfimOqe88HDWJu+9eCVMDXKBAbU2toSlDSvjzJ0ncC5qCK8
bxbHTFl3Lu9x5dbtXTq4HCEkQbLpg4vB61uIP30jis5YjjFhKh8nQ2C0LnkY9Pyr
QpxxZBCdZPNZ7rrhPo50tQFcR2O5nCOtL4HmyC54y6AszazOiU62PgoL+OKh21Ei
l9aP5viCjnD4iJHkhNxjFraYcG01CY6ID/9GFU0eO8beQjTcoYrr92SfqpxiWEPl
hf+Schh6hSFijeXvvZqUJdadZ8oU6iyH21yFU6S3EyXuNwLTm9CUlVtBcKGMNMnU
rJup/g6U0Dr7KGAAi8jD7jrlqm+HZ4IW6/kl7OhfMEngTUi/CmmBcSvqVJeAegeM
I8lkoHgjfqOw9Rt65kUYUcM4z953R1K3f0713f+1cCH9lBZGp1BSajs+aWFXcYgj
u6y/vC0n7ujCRdi8pJB9D5rshb180BQLKhhOZwDmHoTiDf51d1gkTbZDE2LRyDXp
vvoW6g5wQw46GAPDyhsEnQp3WBG6CNzJshI8pN0+OgWXDacsUUT599G8/W3WPiCN
bOsZI/WJ3gfxBClX2Sj7W5nZDano0XP21KFvzKRLy7hyofSWGLHKKcVMVaKLVSJ/
iwhmrI9XbAeHgYJ2hjsuEhWSo5fg0so2KFHgcdnkCYPa8vHHaWcG1BiSOad6Zzsr
lNWG42QgeaVoGcd/lXHrnz/VP4ACLHiW/fPghdUynRTt0cdJBnmQ8tMNzj+sbFdA
b19XrFIy6fj8TIbNewDexbxYOza+0LXvPHk/TYuwGNzWNctuBpaoGUuhMjhI1GLC
aRWUDKdnIl6zDlGozz9VpwbS4Pj8duA0Gd2doQqKANG7g6KaL3JNvSE5UEapYYXi
Ko1N37RYKunXQzsVlS1yJ7crofOntscqOQCWvq3Ntms2zZG8EJlXI8cNeAA7lzXW
XdUV8PcBuMZ/olgN9rU6D0wNXnqfuzKzuHQhTZDJQVPCsnBV4bqA8MW6HJ+F+2zi
a0oArgAHTbY9VhAXVJ/AF+dpr431nkpkP16wNo4WODIrxXPVDYa4KbUUgTDD+EOg
UxJQDBQxI9f0LfQkgXhPx83QRd0yPG1sx0vipG+YxHzzQdtLiH3Z7xSwOnTMUARV
hnjc29jNuMcbEVUufUUUbQ08dGhHdGqK8q2L1aBF7r8cynInJFg/FLLjZRhIRdZG
We0LA2tydlVLrhU71rgjHovM7t2+KNzoTENFJB3m956RcFej4IKE8ZEfxg+u665W
YnwNMIJTSUDoi3nHALj5NwM35JVSomBoEvn2HdsMT6h8NmW24ZO54we2V21VYG8B
F0JBxfGAe7pOgHGJmoxCMknClAD4SEIdHmj9c5L+NV4WWxGd3N4NvivqwTFsUA4A
SW1Bp2tPAtPNIV+un0STa5jlArvUx8iqqdP6Mw8U2BT0hl3IJOTb71e3a91iXCya
fE1wzEa6n4E9itIWfznp/sJ4GQYjc+50USdCyWC4FbdaBQaIKN5C8qSyWt3LLAxC
WfHcRc0BA/iyKHjv7LvsHuWYNh9riX7Esq+f8uSIlSuA7TR/zItvsOfbZT7k4Rx+
YXcN2JZOVjcsbqvaMvIVDGvEsNoZ7EYapfKezENpXQUkYXKgCaXSchv3/vw60fbn
iW1PbbE0obmQQfPgyNvBBcRsuj4eWvZlxDVtfXzzSeHWRH7PAQw8LGzSHK/kXP3s
7o8m4ARGJIxhA9yOfJFRKaeY+F/koktwH8zThw3cxDNW3qxvVWQ2leu2FlU+bZlE
R0hF0/FmYh00Qn3rjCx8Pko2diFbI6d2kyopDkskv6odhje313p95zPeoe7vHTaL
PPi0XB9sMzFaaELflL7VsXcLhUPxiD70Mu7q4Vad7F+zQKRCJxGxfdWKjPxbay6u
IM3DgOnHMXa4XXqxlerW+XXglbM4bVk/oVM+ll3QUF0mBXJ/qY4PHBat5Vb3/dO1
w+EkXi0wiObeD0p9m8rNq9kpdaNcQkPEu5I6JE5NNOkhtiPaTmBbco26YEIkoyR7
kW7SEwoZBUl5Rm4YAftU0dKt1oeTWfOK1kxEqcF9k4jAZA9xs+wfygqHjLViEnlB
hHYTAfaPF74fHGZujwQacgOqO9vGQEfaiVPt3galGygpyAFqjgaGsQqtbA9wJ+nt
XhOLNr532aZFKLqK0qiRaCUvLuvFEZV1HqU25GOGKZ7Pzgx2vjo7GJVMn1mIs4z1
CogdSrhsbSPm93Hqg6llAAUYRS8HzPtbcPEQX+aUUozQ9BZt6TxOPiBSbF+EVFgH
UUCc5Pmt8UR+gMXwoQZAKLLpUSJnKf/6UqAVcScmE0okkJ47tYr7lAvAwtcJzuFh
+Cqh7NJLFLRvVGwwYzxA9RyCM9S8uimT332nB/PmyqM0HcAyWQ+i4pitATEK4mUY
QfIaKsnVEi+my4qUajRMdLH0IIA2bLMdsLAr2MmT4NiXAJkmcPwFZ6QZ0Yv6Awaq
ZZVBGWeFFdVjUJdaAoU6oSPKK4flvsfNwSoSxWmWqmM4EYT2Vs8lfHrbo+wOiBZz
cQAO1LIyC38smsO53f82HMn2L1AheCFLSIwq4U+SGpAYzz2p3cw7qty6OmM2CrT+
Qgh8zj+1a1v/sUFgvF5LDJ527hT/WpH4xVYh/peD71aE8+hYlaljtskQwCqCDqF7
ynkuGM8kMw3eNm2FIVv6/K/6Z7dzKcgGMiWmAu/dWXM0F1ZDhz6/HeVhFYgQhsZU
0LQi+nebE4vGx3g1s30pGVpPjLPIFfVuKf/WKCLkaY7lvhJzJLS4ONTROTNze1Xj
cl1cA/J3Bz3utseS0xr9dtO4OP2iebHL+pEaKAE4KJaqvJ4fjC4kivbx1kK72X3/
Dmd+baBbXas7lRmSLIxacKs1Y9garNKrxm3ETjKINPkiEkPyEUo71La8cofne45N
R3l/M6TS9DROcSnBYjnFiBtJXjJP9ewO3FWc5Thr42KAA+uIz4yVISAoBgaTxXK9
tnjavzIRi6cMii8F7s9K7e04iQ9LY1CemCStgMpPEVY3bRgCqpEfvRacqhle/OzC
dvMdwQHpaOiTYw19ArAQRVR0pCivW97G+MN1o9dBlFQ9zFTbUe5+4hKJqevNB4eq
t83MCo1Q53ErC7JU11tXRRrv/Heh+/Tt26Aw/JDLZr+hvJezzZLb32oWsL1py2D2
Smm5EVmEOq7Z/pNHrvlI4QGfhKrXe6MLHEt+Wnj+KOy0nSCbArzexe2g+1d94H54
X4aMmlkfUEoNBpB5Pe8zThRka4GSaf7eYTv8ZJWZoDGbxtcSYztoSroupERsdsIN
39UwPiwHsATY7yl33xfiPiNJ+QxRErgZvFsvTfTa0uVNODGzeVM8ZWXFwRwKstw3
QvXp3OYSFUQhSsZLcJKKuRnzYj6oiHwiEdaECBeycA4cwjlRfm7mAcqpipML7rAt
btT/paPmTRg/J96iB60krEj2dGAD+MpGlOcU1d0PSRpofUI8VdS+i/U7oRhJfxnK
3zhHQREpvJ1HT6nJ9DVSYT8H5I887rIwPIDfhihP2SUXc4el/QbK4ofS2/28RHs5
lf3NhNftRjtDyGb8Ggkb525zJumBm4eu/8xHyQmsrcNzvHrFEX7N6njUwooO04yT
eizsrUjz0lxBrV+D+/n+vItrHSV3O/lLF35DqVTrAZ+w57TScq5kocLGNSvOwsNS
FDMyShvYI7mMPErLmi/PGNY9r5TJmqsyWm8G+3+fSxbi1RgHqM34ViOO3sQFXzEp
AIzWrQbpkRtrHzigIUrh7eWIiLJyusEKG1pns9tGLEvi3+c8kKhzme+/XxpoVjwN
VuGjAfAxXH66h4StoeKYQq5JLH8vgIjP1XAm4xAPh8XuZtFgzCrV526YWwyKjBXX
SLnM0dKfIlg3QdK07tdagvx8FSzDKJGmMM3lzBJxaVzPoklTGCciFYdDpY03pygd
2mv+d7ONK9i1ONDq9htYI30EhPW9O6pQiM4pGr2AYmoV969rDd69ljjAdle5LXO5
DKl0l3hZQKO+YKzsGMUMWFEYKg7qXJVuqkPWiDSdoNGSCP/d6qZeooa8uQMiLfR+
RH1b/PFfzB0m+IbUHXN7PseYl8Y8tWLmqkNpIyTr/rdMJnWQoPZtx3y9/9bqJgpN
Vzn7/G5xHyDd77ASNyHK0Drh4nAF9eqgEBTF6Eu6U9yXJsjgUHxPM3BoPvMR7GTW
Uw3m/EmGnggQc3J4FgfC7rJ4EuYjRTWnhjPq9Iybxuj0VbstvGli9/SPd6DYSMLg
PBF8xlOGf3KwTKjV+Cpyb4iK23EicUlJpC9Orurs817KoVz97VLyCCBjLKnlOsIA
Ziijprz3ozxSNE5/iqluD/JOvwtMVcCCMOv2Viugbu1vuqkqUELhY24QiwnLhDOk
Z8TThyG6J8sUtG5SxhS8YYiPr2VVjdv7PxgmB3afwkuXnlpSR+dFcOhJ2JrGxrSp
qxBkTMCzJGqFhQ1FL/+AoxNLa8ISyroDkvCa9qd4NlZ1ba2oe2VB1j2JPMWyUhN7
LvDnpP8xP4jMWDbYpftgy3o7JTnnehBVBlXFlsAeE16dBMHFE6uR9vzKZlNkvOfM
FSw2I5YWgHu81wII80NlSg5aTxrG2pYfb0k09VRglRMELf6J2WcW3zNUYWYxHoKA
uOwzrYwh3NjS6bHBemPhte1kevK7uToMzjLNc8dKONTRamfQ90+ZqBvCrcJi5jTj
WkcJm9KFOCfb1ImKBbhKT2DYWMlNqaEBWG67nJIF3ZzaFIznv14iu08LNN7mnN7O
Wnn8Fai7z8brxxWS//nC08kZChDoisGkcnjPowehE+7ZIkpahMaerIIJ2UyWDrM5
SAi+ByxyBMBCbCgkP8AtBfRNUGixOvHjo8MC5ITP0TnoNtLH1pOrLpTSbEYHKMNP
UHC1Y0gju0hEZ608WNcvxc4TNujU4dJVlvUwqIxxKZ8JYF9Kiu4ERPIdVx4uikab
wGgkwUjwCUwn8RtbM+w3/8F8FcbYrSIbzTb7d41LRJ8pl3WspxRYoUffGflvbucc
5YVS1iUcunqFhQCescABl+iXJsGWMNZ5ikM2k4/Z34p9eFUN/KX5z42oKvizp/2C
WFhLhoJzXgVnY2lgJwgE0GlzQx9jfT4iajqGo0k8b9euwRuDfhLB0qYndSs/kJDM
Ytg8D2UVeszTOo6VjBtP3dbI1aS0O4TsqJca8imEuro4NFNVJjVsJyercfWO7j4p
sOPiYV75H3zEzQyVMEfvZ76L18XXB2b6p6lcozTyjtK22GL7234MI4MYcQCCASF5
o9Coa7JwSAT2trmU3PyvUKKvFmMjc8NaG6K0Q5gUNHxevlMOLkrQiGX30fdcf+NB
ObXJxn+gHWFi4O5Uh2zIa4oDLQxryPyVDV/jiuLX6nQmB8n4YnCjA5EGhaNz2CqW
Tti0I0PHGm8StouEFYe+Ao5nDncEkCG/bMM3ljn/4P+7MfwmyWkegO9p9aMPlV2s
8fCU0i83QrXBkdtSo5wH034LomwVT6Gumk4QH87WmClpMYO4kTMKsPoPVXwE++7u
SwXu+TSeeg+vHjyUEvvg3lg0DRLAVHpVaOlRVjg0721KeisaGRPc6/wmIxTOiRcy
MSuwhSUofiCDKEuUj5ZWyEogFKPQhsoRB9sYXtCwssVBo09dpQyzngAPYttxmp+w
O2i9Uu3FsFVEs7p9wHqC0uNZ5jR+1TWpXxecrRg5pLIDMH530v7l08SPE+sW2Jpo
suKWf+71Y1ephhGFJwXXEXxiarvA6xOVhZZHqZtR4D4ws4/kxHIzploeMMKxFM1Q
UseqYWgS21zPPluaFpnI6VHPsluc0mLZxTVxr2jgzvFUEHes9mX4bLs1RJR9CpRB
KNd4iKa3t98BTaemHGrt98vaAhYVbuHVpWH6Pdt7wN/b32foJ1YkTZVFiQAu+7vK
zVdbRlLk7k3DcqYRDGtHsYXCWfL9LGLy9+HRp+5B7qjybiWCHhGhiX9HewRL4S74
fWWij5Bc6w5t/D6IpUZmpQ1Rc99ZVnAwouT6UN7wbwd+SlsGH3TB2C6ySmMRttSu
+thdeze7SJ9ZnYU0eTo3wJT8WZ4CU21K0aippnxOmPEkoaNux4/zrdsImoJiQH7y
0Y1T1XZK7W+VDMQYTpy2tjxv3EWhwe2nlJ36Lm2Ge814qHWi21NVtpx8O+EjwlMQ
qwn6OtLVGLV8ntAMM9h5g+7td3QOjQmw4LOFlbbofUnaM3fytxqBYtdIp5aKKrPC
rAIaQuzOTNbAO/tBt19DBocq7odEccbJ00bWVn32jI1YUoXfDQRnXXU7ablP2ISI
XUwaMyheD4dIwKJeVUr/tHrXcsf65oTjRSkt5bSPew8+FK7D6EJd1irw/q8IFE+2
fhm4Vd9ZFvbaDphjuKJfGxndMAVDeWeloNaE2HR8jEJlnSxS1Zv2yVqXEi6wNhq+
hZVmGM9Vew4seVHwsofzNRU3b6m8BwT2Cxuw1StAnkMBwy+asrI2FZ3gw4V6z6ET
qWcfAuB6IZyqMoLyZUXLVAhwAZws5VMJcPIjmlc14m8InHaVwkJBuybxNkDbRhcq
u31H+iWgH+iJK07SPrdiM9dx64j6c7liXP+4aVo1NncVp1XA3WKjktMJCggUJokk
yMH9nNC632TH7OrQnXB3O97OtluM5s7vNtUlfQxIwk+MgY0phAYX2BWVq34CGoo7
SgcIjhzNsLKxRXLHF1japnhh8q1XuVkruO9cJfnM95ODVnmZ50DpFd8i3pz4cPsr
EoGaZFi6fACGcvoFdG7bxtn/ZQEybgInzXIRI6zSNETFB8xQjpgubfM0FNYFakRt
+HOefLinFBIdr8XF2NoclYKWBAqhP3ZGt5i0D9gGwrH0tfLZgD+ed0e6bEWvQOeK
ZxeJLp5r5KasPqRCdXQOSoG//o3vtiWK4THaAgmreYAjqsXgOLuAN7Gota6HidBQ
PbA1A9q0W/xCk3AyzW5o+0WQ0LcPeyjtle4d9Ya1cwBfAaCIfYjIaF+yCCMPAkk9
WwV8wDJutXQo//Yjx4sfRoDaHrTwskXcWktOIrqjYjZjW8mojma8OCUzomRMdlB/
q1fuZ6IxrZ0sDuw6Qn/JkAihYiovM3ep8BtvnmwB9GWgnj7/494mEsHo5Ca/UQrn
7PzMPt/6wyJK+j/3Dj+tk5BiX0Nm8rXOkQg02ljk+P3sM66KtBrpMpswbWO2tI7+
0rJy0AQK1efGdjPCEsnIe/Y/won5lCBA7QoO7MKTJvq37uevk8SzsocrwuFX6fdO
+90/K8HOYNq0PUdKp9szYCumAqESSMg6OvuFp5zC6t0QuyxtQl6AegU0T+9ctsyf
i2MqqEfe3UinVyKUo4Gx1wK4NuTd3/B+L3XBHwtpN2EvcF5lOv2zXuCetzq/I2Pm
sqxV/+ypVopaKYml7JtwtMVIK1XE2+yRfZtkMvFXUudPbv+I007op2I56EjrzMjB
Mpxbm4EDQ2c8KmAKdCNYbsAbIEkDn0sldWifa3x2spdJ8oXs1elhGBbd901UHuMP
17WdIlbrcweGagrDqnZAA9H/rzD0W7FtIRILlJlJfRNfK+B0MDhRP4EXlkykFC3d
jwxUsblX7qAdjf6TrvAV4KE0ZkxREsPiFkh4aCVVcqdn3LCMvXnFfdocuO2xt9tR
1cclxLfe3F1e4w230EYQTgLsaAKgpqTJlyvpLebKwTu76D62UKtdbCMyRymHDJkf
r5g6ThCoCDTJEzrPgb3Yu6HsO7MRL1oTnYpAIzb/s6ZORWMd0hKHm2jCGyJ9X8a4
hVUz8Wqe5/Dgkvachu5AWJkKx+StaNm7Zf+XIfEdvO+x87UyeA64ksRTjTQofuH3
4SYNWA1ZQL+Wqfh26Y4f/zBBdgyg9hyIt7b2bv+wmD82MA81Q/QKieoIoJrhpwPd
HRNYab260A3H9zOkPMU79RzjrUI/CPs/KGN1NopNuwhDfB5fg84b/Rc8aKoMD+T4
KL9Cz7KEjVmFvVfVNisAljrnXnxsWS1RL+J5HTWY1Y1Lvcxt/0HXbwyPRfJM6Hau
dUuGj1jKdLU7prhMlk93icJlZv1DpnjJARcj6kXtD2RSU4m25eeBKgVtC4YeVdM2
nQakNbrOuetJyTPNNUX4gby2i/ZjgyFjfKveynpo0PlMScwlAB6LzaNrbtfDf5rf
grM7BZjMGoVGJ0FywzOkihjS8h9I3p8b6gZhuloM4TddEcKRvtiI/pu5AA8AsMQb
l4KNzgTmcx36qrPSSo32qs4wxQBzjkMTJsEn1qA2HWJuEWkbyAqHaSc9js+yMPfx
xwYKwH2RoX7N5RhYHzEZsiP3d46DStne3yamJo7/C81PUf1e2aw2kzKGGqWUM++5
44LsloOLhwS79lCsNkEVs5IfMaiJdi0597epulCjXkRIXDgCA0KBNC3Bw0CFBXYB
v6Cc/omskExCF1WzCFMMnRzkjqzKrvih+EmokPKtuiTYe86wMbyR9/ZUIKrsNcWG
tHZ4RmzZ4vbzyq5dTR89uY7F8J6JMz88u7mDHIM6YCzEFGIaCfXPvR1zLnlZyyc+
K1gwsyBnNYrXdU6HKejs6LIOhc2bpIRDoi1m5NYfLYYOhKIsSi1z/LRWRcZi0lII
4ARM2J80BllcprFAj3xbSZfgghy2/+TeBw3cYAzqaA26+mXLTlOC7r4ZmVur51H+
BWRxMBwG3KJTdz04L/DCP2jY4QSzs2DG7nKOQjiP+rVXx4/PcK2jfevy7xf4NjiW
HbFs4Mf7RQKJjk6L3APxcnGMiLpWqG24Or58brArebVb6s300OuwBywLHpIbfnI6
XVeQpIT3mWmoU0wx9kwNI63rjE4zVUekBiDfV1hsjeMPV9E/YE1G0V/0P/kfJnfi
Bg4LHPv1R2gsbyG4q0zSm7TWV7+syVU2k+fP/A/liavXUwsgTsS+7BsfGXq3qm5U
chjB6XRS7LOJxSm5Esz3XXDukYyujP9mqSQdHiJmpbyvrp4im1bIlYPYoeg2ecVA
GFpSA/xiauobJw4hZ7+fL/kWr4srKQWQR+q6gf0Dg7ZFxdnGZjbvZ2l7+li+DEZf
IB7BX5CrHFpzW54gl2TOZxYfBiW+3iPDHdg8eKQ06J1XMQCz2kMovtsRymoQV7/K
YJSKf1VuuxK3qoQJfnWUzfgGx8MfdKG+tNwx0eRZvfW06zZsaRFnp5nziCMao8LH
GdRuGomXhnCT4uuZJYRHip8DjIkPfFPpbs1KYxZDPBPWH20Fi70I4TudlViEa6ek
nhcZbPxdiM0OlrhPORBJfS/+89Jz3A2nhaZd27c4niuTCjcfWjShlUqjXGjHncuz
Rwl/YkL/v3mzzASTWS03Zpa9ezF3jbirQzYWJA2fKXlzQaiyByCMg3+IvwSFtxZP
dK4ILAiK/jpDedBzqkQ/qWkjTmW66gmzIATBEaeWCP4yu4PaxiWxB65jO5CADk/6
4CKeiaz/Go2I386M0mz1FSsueMml6Kg1KY2iiLTtSD+IgcqOXNe2Ho40al5dttZP
/8Z/PU/NkK4wY1ceVpCZXnSBUYP81tV8+amtS2DQ42CX1l7i0qliQwwvaJ/G3MWJ
Z4pC3oaOSwwLU3dWg+lnVii+gGr4vU33icR7Jsg4qJQEznPPA9tVUNEdgzJmTWR1
bNP+MsBLZPvcTb+UkqwGYW2GLR06f0OgoDcNdPiGHV7B96tJrNhVfXq3ucQsGFYq
9KMrDwzqqu9MnRb0RSYTTw2YYkuFj2IKNrhxae8va34129UXYWNY4lnJEB4oxQno
ZtrNsj1gE6YsrRmiMrslShW8xeTAo9ErkEEuSon9W9CJP0ER21eFQL+HGnjMKdmQ
q+18BqNrGFwBUtfHtcJGKrdsLlGXE3YhUIvvQPwREbrYq+A53Cn/qktqQM8nOyOQ
`protect END_PROTECTED
