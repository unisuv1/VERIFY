`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yRnbxagyFOr5QI+cIj0BVBTcsq2M8HK9D/6tlFbnB11SN+xaNMDaoB/cC06str9F
Fya/tJZcYvkzJT96MyNB5H4ffhVJgCXYaNdeVKMHn1C3HaddErh4sDnZlVhdlP1w
LjT8n2clF6fJxzNcXtFy1Z6lu/zmorpKAxhQBMJ6qy7wktArYLjiurrnX46TWXHf
MGe64LKprW3lv4D/xRicTqOZwHfxILE0ZnY3IBR4R7NTEqdVI4ae2nkH5t4f8kMt
YY81oMUne3HhgRU+KlsiaNnLXilqhp7Fdq1yh1FG228dK0JxdV//ldudRiSso4om
IBdqbhgXb8+p7kYV375RnSXOXiFaPa7alN4w8EsgI2PmqEyNQnOgUYM3CTnZlrxL
QAM0ARROs9ZZCE+EORgC+XTVPFkBfkJT0Y9m9yW5f0rSgsMUXqAXEjnGX9VksywY
zb2xrYSMMCwm6YE+Q9hHz/Lrnwq3APgqyrjO12IH3x0B+eeb3lojukusazZ+AEia
Uu/AwL9wFzupr57yLLNlllc7+7yJEDwZrlF5Q7Nuu2YbT70AVkhbRzxE0QjRLfEQ
w3tXsksRSH9QrhHjIN6Pb+lXotmKwlHa/G9+8f3nPVxoKf+l5KuGVtGnSPmI7OB9
COLSsOy6JG10RrMF4BnRx0MJbldXN+MeTBzgKr1/PLqVIM52ZK6yc6msp4r7YQND
ktnBhfbMfZ9Ijv2dJTnvALDShGvlmFtFMLk9IFKKwm2UhWBW1/440KXgM/7uGfAw
TRG67PyCJfyLMFXxof5JfHvt/ObniYXrwJAvrgPZGhYfM9xh45+l7wpchj6dK+i8
+zJDEDjsdNdRv2H5js3PR/v/KkMZSYpQmxUGopbpyPnOxZ5BFGK5uba3bBuEkYDu
b0mY1/JZX/hMBtiTc4HaUE8frLgpGlasd+KoaNs7w6q4LQN2BUzqo8xNzynljya+
SR28JR/1lAcDnYnsNJMR6Xuc5+Rw1PoZkbj+iccHi6WYRUTDUieY/01gT24X59tQ
jkf6ujp0TACiuMKq9xYgRwXNvmLVS1iTxP/C0SZnEV7a1v70VXgfnpBRQURWK06X
1WN+EdEncE+dzp4iBHpvW70tGGQQJwbf2v84xhA0GxBY8YE7LiKuy+MleZIg0liw
Mer3FBPr6XCh73dj3NkUH0GQj7MT6sw3/i8l//ZzSn1CPD+5dPPkcFBpDWqdLg0/
J8bmR8ngn5j7MWA4i1EvnOMkIkuzqV5lT6/UidLErk99ZPyzECe4NLeILp4YNXDv
78TX0BHs7+ADEW4Ge00gq1pEgIi73S0Wb85BPS+SN0OlxQmkLWakWJp0sx3KCKDP
7EXz/RlU2h6TC3sUFbI8f1avMkLO/sHCUkhx+H/GpydtnD5d4yCtL9GPOyMF5ruI
X1CT/WjRS374Vs96WfJin5u3PNG2y4R594sLLkJXEc0cfdFzlPMl3ugi7cHqaN/u
+8kVJ3NbR7qjZ2puSl4NLm6qv7ea4Coxgu5H1B6rMZPouG3HXlhyKmkJLJx9TUy7
iFkgehJjO/snNJ5VIOb9WwegMI74pK0RFarCT9p2SIW7A4OMZyPQ32lde4Mm2tr0
g4U/VJKBQrX7ejmkYogRZuzNisWuk19p2zSyoO+R3xZpUzBqckjDwpBqYakZzoo6
EHp16mqZYFHnP2e5CmAqjrUMa+4FYS0yT8ntUqRhdAguSIrcbn63C/mk+cfhdiE3
YMdspgQ+NL3ggIyojy0HbQ5ktHJ/cQqyrVsO1hemcanC18OgIul7Q7FuS6vYHqia
szXhpsr8ujzkrQYqlK4yO6Dea0rOiu6lKJX9lUIObc6h48niqHqre2R4epUhThCt
PLH+9AT6+lNLm3uF1m2lU/tVJnl2k4QXl3rnGqYB/BQej36q4jzlj1nWsutN2tRi
FC77MfmE46eGFHoVajAMcW5bW/4NYnbSNi7xWA0+sGDfGSNp1xeV4bi1dKBDkytu
7oNSqn2WPsGY/qqsyPkt8l6MY2kJccEwHSRwW7XmSbI5QbtPOW+CxwosRNJqlwM2
ayh3CPIeS1Hl36bpFz2XmlzMoI6k2s9ZrIRR5STvgIq5E4ktJaDFIwRWWP13E/dh
QiyTsHT/78OhwyCNAPnE3JjbGWa6ZRK2d4IfKLF1HcFAXTAxNhTT/p8bYTC+NSZH
kqN6aoTRUrLEef5FyMY4NQGgeOR/MwhQHwbxEqXTZY8p+SRYBHBPkp/op3VDyQVm
ajpPJNm66/Tjll+RlDmsg7N5RHjXMiXUvWS0k7roFATTaD1rp0Y+CuTL8DByVIpN
3F7VQzjWYXMejfA5CXNN/2uL93O20yXaxqWS36hFYaz4RCRqCiF3U1QMwMK98A1H
9BKfkc5/K9yvkoqJiB0cpHFjc75M7yGzllBefr10IJ3HBJTh4yDjD9zRbdh4vsMX
iBF0Q1LzSeW2YMkPC5ZMJ2ps2eFRS/skNcj6SEexNlEmJ33plN3kdY2PLvVRlIHZ
Slgur4Ua2AS8xOjXd77flH5emAT91dX1sdeN+7JHl4y0G1BhUM3b7yMi1+Hlm4Kl
FQc3hYpql1/NhrDpG4F5W+7ioVlSWLSwQGwRKfUkwjInM6Wxwt3RnMsxPAnmh627
29wIrQeYAS5LhzLm6zgSGT7e7S2FW87uAmxjvrkJmrb4OmjWpigsjgHBEjyT8YBN
qGlGRaEk7k/THZnj8jLBKtYJOc98TzQ2hVmXIkYQpFadrMgqthdI0U7lgykcoZ0A
V3R2lSGArOuZ21tN1rXAIrIWm3zIvvy/nIvPuP3sNP6MwyurjXszuNc7nWOeEk0W
sekbJ5b9T930rDATzSL425mTsLzKVtBaz3MWTd4kpxaSb/jksM1s1u01ge7SVPtX
rgD9giHKHsbLkikSZA1nDXYBhQVaxtbn/27PSo5sGz0njr4QfnsiU6/Q+ybGwq7o
jz9yS3PZ/vtoIfTMzJpf4KS2tpLU+2KZ1vDC4ABNGrShwAIcy2JtDtw2aZvM8kr7
PWGS9F0xopi8cM7R7Qt+7mFXKDjYjlmSZPyq9p2GPPPdfRDjVnaOu7SYPmKIFOF7
BiQA5cv717CtTfZgMH11quyGrw0NuF3qZrpli3nepOzmE/F4VmEyLH3xVT8lRF4/
UzqTogDr5XuPuYdWYbffpYP3G9FWQT9n/CMnR1mYBqkc7FweXrlYSxWn7GyYv40P
viTLecLEtkn61np5UAN/VVz7l6njs1cypjdpbcS01mXd92PUjvxXDOAEpNmax3sb
NzU16nznKZl+XhKMlFwXSvQ9ZWLFyXLcKdLAZk7egHyrCzxUqDD82qTn2IbfEU+o
XmnLMH2qtg/RYQCHyBzp+7Qw4L1LL2Ujr8Fo7qJtCVv4+Uh4hJPmD3VnasAd+tby
HVLYGfSE//b0sYFGnYRtEfZlw49QBzeAlc/GID/u1XaeqFMFXDM+NVrXmvPkpVIP
RMXdU5fMsnwRpI6a1DWB/2JenNzkypa356H3UZ3Gq7tRAzoFw3h6ls95s5IF+aMl
IRHq0K7jp4V5mY1JlfsGbv0gy7jHBEVpQOa+mWT04PCYU2HELYiS9IvSTUU+FH8R
TwY+L4Sg/kY1U3ObOu5tnGpTVXmHWqfEeyu3pCu5BE7Ooh+nyAKj4iKxFgVV+Mqf
UjjxCvafZzxwCPQAo9O4c3Ex5IlcD37UhZL/YDmfEtp9Yg6cX2BorTmLoYvMeFaC
3ShB5a2nSdfolCJ9XZHE5TYkSYR7UkHnTTp27fcTzVNDrUbXwJVh2JRBKoA5C5de
nugnLUgL9xk1gUTIPPxnHc1suvjqtAOjzgJF4PutqqOdII1GdlMSUT/xrS1FvFvN
03uN9Inc0ch4yDc0p3QNeizslS1TQ+MR+mTwDtRhjMyJO7CqwytMb2T++oguUAGT
BM8aPOtuXrfylJbTxGScqDmkFB0t+ESwH8TndUnYvdOCWlY+fDF0/jOuWtS215mR
9P8hWy58QPIdWn1IQXkas9WvBo2EmQyvtytIxBH9zSsrdZYpChMztm7LKXvybTFI
nhQ3uLkPk0TCsWbP2gU6r2pnDf7mawFxeF6fKw6z07LORbURbmQSKyNHw/6aEyNq
mgI/nfzz3XRyKl8neSZ3b/4Q1Md22+jqFr0Gct0UES5PCMXiizF3JxYXbMikheDt
ZGWFnBz94pyU2iR8+XOmVGNwqJQhmzJFaqfznZ29vITOmOloyWlzkMFQwMD8XE9J
qjPRQ1BTDcmS/fLs1lmwIDaHw0FJNYgand+gcolwo1CzovP+Cn9w94Hpvkvz6Gpy
ltKH19RGHO9pvznwtsj1LQ/2orotr2pfkMZMgTKn8yaQhqIEgO/GCpg4rohy+E5X
jSUfj+ya5IWfHN3p2nAvX64kewjCflqmxsOWAM2k4vZCVVG2NBRhQaejx7SPR5XM
QJIa9P7ueHRFUr+ugvSCGtvchvA9NVuAB6ei5/TzlHuThFMzyiM0aFEZf897mIIz
XjQ+3+vzFieCmQ/6afxQdy8udcAtPJjioGqP83HsP/kEJd/i/p4hE4Lf0i5ZF2EN
uEr+PIUiPIwduKXI1+zxjhhWLFrlFX5pOs0ccDt1vsq/us8QDsWaOPQHorMgmuhd
Qad2N4BUaOLolrV4XQyhkvP1aEfu48cfWAtLSTcPio5eKW5ZeP1IThLNahzVOzgk
+l2r+lZRC3jd+5jEymBsjqh0VAtoz0xPqzv8K4cNvP8EvihGBcPXcjp2Zllh5esD
sMpAEHenpR+G0z9997DOBGtXf/YT1ywCzCWH9cUXHEt00Wfzo/P5qXf0JO6en/W3
FveOp9DBoHnIloF33GyeuQePtjPIn/4sGpiAfIpE1R9gnVbEqhpTSVD217C7arXL
790c/gLuFtYzD36lSBGYekg9qYyrJi4NGObXo6RiiOzVM6AhBSVpCInGYayIfGBR
c0vtkrPRmM3n37x0kbuXBvJRml6KGKgwNhkak/3wqXsQa0Iyf4uh6yZYULdyJ9XC
tjSMuIjgKIFV9n8HFc3lvpLA5PqECsM7gxX/fEULASQyAMMXzpb6D73NalDFcQmo
oLtq4QZyob4f1URISGflGQHJYMjuJRyMAvduMG0JdoVle/tRohDUpNfrihRaB4qh
tEHnbsmkqhcXzOWQ5LikzwML1FJ2+N0UlR4PqQhIvY7PnvrwMTEKcaAwp0Y++vcV
kLeu1K4ArSfgovquNyCBrsEIu8PwsFsgV0Jj3VdASzTa/tLdJlxIgC0137ySY3An
HAWYyJljy/7Wo4R9oamkt+hiIt0/OuTPO/tymZT9+S6m7LBkcj2iHxEjhWezxQ8c
V78hZkQ/OCWGS3zpKJg843cbO3niKiMMjmxVv1Nn+uU5l44Li6roYSc3d7bVv70f
uv4L97OCfdpvWMKgX/ZogCXo13ExrQumKhBV3rX8LfxpoluVE77qy5EPe9xcsQ+7
h3jyZ0tE3+yH+uiMM9JTNHlh4JKfA8XB/0GC+BIV07y51BMvKuGpa9HE6zQv5Q4F
JOP2Rf+FanYHoMs3jKbSDLckTPEiS0BeXh01ixY2TFPbC1FgyclWgak5hOJwBYn6
yxLKpBLE3KhEhngd8g4HtRUn9dZ55j8MhlYkZCmVrpG1q9oeHI8QFwiNY1fodkX+
2/Pbg3vPKExQWomXRelHBwm+De2sgJKUoRGSL6K5+97KVP8+flWLcTNX6wQPz1F+
kAF6nh/duddEWc8F3WqIf4PnkAnK4tQFT2woNGOMxCqNjRL6Cym1vlSQDLHvJ+FP
ntZ0BvLhr1R6qXsMUPPBhOzS5+MnlGiJDQvLOpfgTBufYXwqPGiIduSicivFxOwr
iq2cesu3pxF+sW0u+xbv5Ef7Vev3CdMZ9brr+3bUGj0XGkeBN2MavaqnMYKMs+Yw
0YMI8RRiRMcSTa3tuCFrx8XU45ByQ8uoknTVWkYC2ND1rX6D45H6o1LA9nHpj6kq
lQI8jq9lIo5imx8S8CH6YrgXoYzlQEe80GHs9VIxRdhPLOwBPmkN61cWfWVubvst
CvqCm8NDST18lOqUv45ZgOclVCZtBRAmoqEljgxZ12uGJpWAYms98V19+JZDxSzE
fy9dGhisnv+UJHgBdNS6DfV6m4mNTqBd0JPNUoTo5gCpRoOpeE/A34aznbg/xo1M
9l3vRY0DI57Jxa17zdFTKIpjqSEE+wdxaFZ5VS9UP8wFMWDqkknoMPU7dJzk95O0
1EIOia0VlL6S70JdZCoGffsdxB9DxeT2/JKF6z9zFxJ/ojAj93L9MsyawQ4hKa8t
uRYD1KkIULUKu8CTLoJXbL8+0jgqQTsaDiyOcUF/ki4rmxqbPAIHSY+F6kxlIg6/
YM7BzUrNZZF9Wbz37k1hZ6Ek9NaUyO1Xk+43Ybt/vy5sRc6B4DPq5s/SsEC48nSs
3AjC6+Do4Are34WQUE/4uXwAfmK+dOox3NS1UPvxTYIZwziAXrZiX2cnyF2JizzL
BcAD6211VO4hDR8R+xqU80fuQvyehbGgIl0ZYrSjBtP3O6v0kYVTl5L9l15/p0AR
GyCxlsa7OJXcGLzzfGA08MTSJYV7EF4N4kaQIy4QjHVbMWq3hRBiVJNN/Ygp8AUH
/2ogEgwlJqqzF2+18N3bzlO7qJpY4XtcXIR5dA88qj3dMubh7VT2+n6BUBQrwVI2
WOo75bXEuEUo5CnlkRQF4wrSA85dxfYexuIVzHZ8POR0N1TPWTgCGn7ysqYULzjU
icBR2JxvnudZo7ubYQExg13Aw4i11jClE5YoX18v/i4x07/EQh3MFE5dpfgnEK3B
mcReJrH/OiOyMOE7FhDuH8XJHcWeV9B7jAM07/dqFTKczmxM9Afh9hsu7EoN929I
yCKZvkq8b4naQAvoo6mMKlq3jH2jqjFSjUMmuHGmQPYJ5vHePKs68gU1JvtD57/N
K1F8HMNjDFeKu7QHTgDf1j1bSJcjChLBGcvYl6vrxJQwPst0wSYHKkNNUqUj8oWc
rrsZ/4NYmcE1xGnuO1PpNaL0/2d79rp8SrRKGoDDmFFSJi3sJDltwjy4nvz1V44e
WJAJU6SC/eSyLn92gqfrjFS2aMvmslcx+agDNkcDQZ2cwwg9ccdmYTZtdUBaj58T
DGGAgYTra6vEZ48d2ItrQ6iMVC4B4U9Viip+vm+Zc7i5TySc40TNjV+DoPmTIu+Y
w8axsBXFkn01TZPENynH0xRF5FEH33yEqRgQB3oXbc0hRfOyKeTUmU2mwKlVDgyA
KIh+ETE1/uK05MO2VilExHT3iiRU4OazI7G+TOvbWjsNZcPJexuRMhr1BHiblJbN
+gLbKDtc9OJncyGL/ewIWvyds5lRYxmfxkHWUjqCS+Mdic8EonQnVlzFQDFEQZh/
mf4uG9XMUxcixkFZJNaRW9qC+YxekxsokkpXyyzbIN4vGz0zuukeDd5gQVSsk1En
zFDOGd0IMNCR9L8V43U7ejP+pzV3nMJITdQZmQ2rMyHn/NA1OBVPkeMv5qIFnpL0
oYbjTcrMwee99IXVQ3Jxw3IvpIf45bE9lP168dPjQ9NQUZPWqEM+UCK10PT5HezE
fVkC7/8hAqqZtG6/6kPr1nJ+TcHbvvVuHhfNmVEw8M14Wq5GLCWMg30BDLjdtMoB
3rmKRuBJD+Xf+EBt5Cx1F7n4hxE4ZlEAnrK7qDlTM+laAMV35wYECGOz3L1trtwb
01GuzIoiBl4uYIpvhLtVACR0fH4UEbxr3DAlKMJsW+PJPCCbPCfiR4/jY0wQNRE3
YAQO14sCh3tWmA7EBOA48xm4fJOheEnoEXNWiI9QOwc0IKqoaxxId9YEf3bJtxCP
/3ie6A4UPHQVudScW8maYAWWhIO1Wsr+oXX3EUVVEd1fk/f+XqMz7nivxqD5jrwR
6+0E76ZNHuFig37wXr6RUCiuA4I9H4gL0g6GiUSZG+1BkSNNY1FcaGwFVjY9dluS
NBAEs0dQyq7DIhozkOYu3iMMcAQQLZmS8gOur188gdleM62R061wVpLg0O5P0MWg
yAwOrtK/t9FxNDREgCq2aEXBWQ1f+DtDdfo1X/6yV5OIMHt2PbaUQ/2tXRK5cUlg
Gj2Ec+pHxCL3sb3KoB6KfvbFyswaC6bgfhmYzdQL5xKO/4u9VXV9iPSXateuJfNZ
RoPYfQ4EWC6JxQnCCBC9t3nxgMBpcfhQ/1l7uV7HUkmvg0tPHZJYTUOqUqeHJDRy
LmVx1+ZLkLP/DAsmQE0awMy0rH7bOoikBeg0G4H5N+2kYcLOBSg9BHaOj4rDnxaJ
kR/cmkU8ISwqwFCA1WkYh4mw9WqhoIyjuhw4p0AmTWHKqa3Jrg+R8fvwSwxGVSV9
6c2cRSMdtLiYXApQtvM/KKOc6bOMWGtHCDmtKcAdqxEIJxw27honr0WJuybmn1JO
j/xMSt9x4ikzG/ewiY+PP786172Fp/R6RvQy3Bul+/+2YQti4rrJP9wn3zJ6dH7B
eFDs0KPBYuO31sApSIbqBOdmEyqfwL2hhhSxVz9LPjT7N5nWHZCMvRpSH+IOUU1G
kbg1RQqGfjUYBvf4r1uAv6yghdVLK8HLA7DrHmQJqOeSTdgkp5187+8zxxF3PYov
nsap1yJLufSS0j/M6xuIFTd+/fLXuwc7aGFu28+zrs8axfcEWxFuleD+JIMhv17/
Zfe1A2xwDBTzoQd8HnwJ6enW0gGha82VxdGi0+ii5a2RRQOxa2ZvMKDlsz5KibiX
IeDPe9t9ziELftHiEogKEFFnsJIMcVGCnKGBxMAqwAaqFiuVVmGK7qbREneJ/lLQ
T/CvsyNNtnyHruJZrpNJNfnBHJaevsJy0cGk0tJk0aMJ7VcAiiv5iMnr4R/CYJzt
kQSyKN7MLK9Amd64mBaISgokQ0BJdIacZwVmkU61aYK25wA6IEgOttTbel5m+Zrb
6/NgkoIdO9duoMVryxhCk31rdAGQ1dy4TlBDA8KQrZEUWaYvcIfNWKvTuZ/MPb/h
pMPX3qmoAzbqjO6Uv6JYdi7LkpQKq7orsLYLR5GcPQY7l+bUSgdcyufN72K4a3nq
7heKAbBGie4IfwxFAZwIBXlc2LuS4WQJnD5S0yfECD1jbi/kwO2Thn6hKknVC+AG
tzOoqchRKYdVyeMgG7kF5ExZxvqxZDupgNH9ME+EaXAvrkqthn7bSThSXTTYHl4D
0VEg1oXkNYLVIKdyVysl5wUsLNEYbjL6IueHOIjERJ70COIjwvPIZloTNv4gWrXV
yhhBQ05DjnJgHNe/mzJhdhFbQcgqCXZOxsQvxKhsELRxhjK8SVnnMtzGhdzxGNLj
eT5cjYh5YB3mpr6t2K/CoaUzp+PmHDCSXNfbXxJ4OuCjdrnwPc4av/5gp5S1aFCg
kIjdJlu+HevwVSbw5P5b9xxAYMmzEcn3Jc1DQz7tywxXMfNVqu98YP90mJqODO7Y
5VHxMKHAaAN0O2/9J5pdGSuCotwkc+xHHvua0Ycjp9ZBBZh6Vsw0KKTa2ay8ZfOp
sfyqKGXy7oEn0eTEmplUl78ja2VA6kVU+pwmbirIhxHEzNgawEYI8ecIJqk+gIRH
vOuOWpSMOBD7SYQAL8PUxqptjvZPYkaWKgvv3Ej2avRrdxTr8dJH1TSeKGS7G9ji
tdWIHTW0Blaj+gykQCwO5A5zIzLTCxH8Jhtxdl/oFYlW1/PxNWCEOSNPBF+NFsS5
/fhbr0i0b/zYQWF14eF2orvt+r2M3dzY1Y1ZUnW35HxRQmOs/FJWQeML0hxYgbp8
34gi2mvF/piVEJTywjMOtHYYwjXPu7AxlZ4D3/2SiiMK2FmU2k98qbrckAXUhRdb
Px1KuttIci8qUKdsmuEJmA/0OAwISSEs6bKGaZnIKLBV8ffaIRkOY9F9DsZkZOh8
oR6RaFPD88y7NZ13MNMjvD4AtbHVVu4ypO/ZYaMK3dMPA4eES447N7tD1pH9vODC
DKK8/TAAD61uJupePSaySiWx+MuItsNANPuRtjo3Uuy/Gr2dG7n6UC0d1jorup3D
tctC9JL33GZ9qRRrxUvL25t+y68eREwM64BzPMtWTWlhUQUIo0tZnDXSHeCrMprz
5JFoyc63aXHFtABnE6NsDwh+iuzTF9BzPSUv6G/u9+fmlt5hVNLSxgFLrmSTmuIU
hJdMXLcMiA0sIB5FdYHgZsP2h59ZTyv+8a41Z/HCRQFTQk6uhUmPgfCcywJH94gT
sq/lUdKR0WUyiO3KnD0QHa5SN6J+hmbNvbXDl7O0nvf9W5HzkqwGvUGkZVgzSYB/
A12GxJGJb5NYf9qS6Sm8w+e99fD2xqD0YIoiXGmAFAW9ky/TGzcGNXPJ1b5YJMMW
MKmZt+ktpMI7pP8Oju5L+tSOpBG30n8zowmqCNCOjDNoKIMLJPySMYPLxJLIlDC5
PZV7/2z4IitfeaNfKn6kej51DctG99M4tw7qyezkOrgnruOr4BX4598p42+lh2ow
7T61q3u8N/KzYL/32HP1M2xXOr4xIRJGZvYR2+8d8tf+/ZMfWAZEHdp3gLbIBBD4
WNrLEqkV4pGztipCm6IPt1LyLAwWNZeGixDYd6915+b2mEMMsYmsKKa5GtNRbgL7
zTYH39QntvMqsXinOQiQnCyOT/ToUwOmUTVsD60pk2ZvieCdUfILMAyc6cq8uNAG
616XNQqcs6jzMDgYk7byn/p750Gy8P7wythYA8NGLVp5HIngPXm88PSKBIMPlAtH
K3dCgrsnFmUMHIlLvAqHR3iX4bI7cKna34u0DEtO7g5tZux/yB0vpWPFshc+/2OB
56fv4STNi1e5cWUuqFNDJoOfEFHGa4zyGU/pE401IvSURL/CerAvWuvSOdE8dL90
TNJb9BSNBmexWRvW5UrgFAU1/YQzqE1ELEwR1xjkKpsQ9O4hh3CruIXeop3i+WL5
LIsT0fSI39jQhEwXDm3BEXCGYxKgT08wfzwuEH/otlaW0Oe822wceURrIQ8ElRWD
yIqf+jH00n5WEbbt8MhyQ/6uxTWPbIsHRP+28sODEy/Wp4QHQUn57jJSUvUsm9Tm
t0v3zr4iiU6YXkwADDduTyTqTYutlZtfeXSw+iDCjCPBynmOHn4SVHvC+AGzAYr7
6/4zRZ5jjemMzRsVM4kWxuJcL2hSBpa00j5qXKB9Iq4avxyElGCykSrWOuOYHani
sfTAMvIDS1np0Ale91ESVc5M35uEqqB8+m8KtK+WaNbDWOPJh1dsXeAZ7RzU6SOM
DCpqWvXiCt+FcUDRMNCx3Q/vu4bxQ3uEj06M4RTYCVj+py6vkbC4Qf3qUS5eBoXz
dA0cScx7khU9gfxnUCI6qqGdUMQQgJ4loVTjmZg9IVkfDgP5VobsLaQP4f0x6q29
gqvj9S3yRWsT9qys/6InjJbrUZwZ8GeWoAKwas4u+XjLDETQAW5/FXtRyoO/MRzC
6AewJ6u0asfI0VsUoNSawgY+6yMofgrevCisrEeMXPH8LihFGIWJGtuAcs19DTR2
1fVWBCZTajaZOk5ZSMam+7PGIQV3a2gnDZbf6nUR6M0tgJc0dRXyCKWGe812zHo1
w/oSwirODZrpermti2N/LTH4a5NVKG5P3NOy8wE+U9iTWw5x9Ou+9qNOf3e3NlrE
0sT80+XzLvFO6ZSEcO0Cqw+3gVyr4JbGV99pFgbF+J4OmjtGG74PbxeIy4A+vGHm
inNUnQMToMD9owedwXZwDfxg8A/zX+8Z4JzDqXUOs/cbinx2AKhoD+X+AR951oxF
vuZ66Kf/aMR+gSrFkMI+zq+glY1CufiahcwmExliKbSqcKh84z7w3FJZ8modCyK2
hHcWnsX7oiFSXLDB7SZxw2E9O9KNFZYVXufTr/moAV/9tm2vTttsCsNH/WbObm9U
j1gtXw4ddeu5eBwTDiZd83IzB+dtRtsjSowgGCfjqF6scrNOdXnlev4rttyPKVRD
/ljJwOFwmG9z1ED1L7f0MOlwxXR/EEK0WR2ECkeZVmtS+v5QSrQ2evLSbA0pRNqV
pO6nbYL5pe2On5p6G3zxvfDKxbqJTC7sbm64aqJ4pwKARiWPeXPI0L8G1kxmoo1/
ooxd7e4fXD12gMTIRnKGCHzXK11JnVu36NZG8dw+INRQ6o6Ne35pS0EGD9LGYmn0
y7BYsCUq1Y6tQ7ULjjz71DJ9hTC1ZKYWSbwdGofQCJfphL2IYDBxqLIJFSz7jTeh
AUVWt2biv/SyILyWenzpEUo8mBaEKjv1eXP6S4p5ay39gq6+SuM/GecK8DRgpkUk
YUt0i9XnYSvJPvmusrfBZwU+gjSpDN51sVhr2GlQaZ+atljYafbc8pA43YCKd0MD
FeqhhHZGsGxWIo81j5dfwmDfhuMqNv2I0qpF7qgPR1iXWpTYak/oC7UbZxICeCk1
quyY7x4mN7eZb1ettDEsJKXmh/sR26fkwABM8y/zkpuZmEPawbzLRzorAgl6rWty
3jW4Eds5nN/Ankom3bSpFHSqSaGrKIxOz4xfREW2zqIawVhwA0/rpQj8WfGrPNig
+AFrN+96CialSs27hYTrtwYxCQYqWgalG7Drz/leDC622lJi4Dpv2IQogJbon78R
6azxPtJoTe1aVfoUZM5uG57lD19LFfbK00RYAkdU2+KRwTzZwmv68hX03Gk70t38
3IbovbApqnSOf0fm9POrsxta5mMULriR11Rx0pS8w1A8WofBxrfRLoLyRFyOCug9
L8MoldkohsWJ5NuvVZJE3Ld/o6kvlarQ+2b3P5IKFHWi/BTA9G+hDSCKpaJ1WwpL
1Kf7+vSqDM16gBa5qWfgFDoZmWHbrWVIq0Uta3RO/pQJ2UAwfc7fDDTUL2Z06e7l
tcKqv3Zlxs2wnm6t1cT7kJ3uMWdw1/DSh8i8dAU5BPhOzofVexbwtTgVIRF0tXZs
LHx0kYCavLwXys/FVS9iPr5E/Ue2Vr8WLHQ4YUXfmSjLtD7gRKIUuRBTbdY2wczR
Rv4JWE5mPv2GdkKSFg9WyBM8spel15UhwTBzDhBdc0e867twpEd/oVizUyQAU9/t
HZPPXUtYySPIean/w50Ekg+bJaQ82EWgAmeQcTElyQIqBPthqI/37emiOJ2iLNvi
rpY750S5qu9SvRpaEYhBVCxxRo/VcL4iwO8RwXOvXhTqP/xoVad1MRUltkH9lK58
gy43pFp28QMDj/PhSOXah9gx1mlOdR0t4OFtBXxkdSlMUCEjwU/WUotGda+K3ZKq
+FoLAkUBn3hD4upqwsBhYXERTjBVZwZo4E+RRxXSKmpUgTJNpcS74TUX9ZZgffaQ
5b5J5YAz4gGKt2TyIuc2riEySABAirbBXnAm3mrr7ak9e7U7DL+Kx796MVq/FkbW
ycmyBK32IxSyZF9NkBBd9nU4QuWZZax9fxVJncadzCMXZSXqgd0dG0JlZRezVwIw
XO23y6TY2B4YPvEMablJdthMVLC1ovq6u8XyzTkDcuAv9qg73lyR6RbFXQjleQ30
R9fu1fkKJic4EMgDd/iZcKzy6Gxoq11lAs8QFPKsjCp3iHfAQz+gwrzujmVsgH05
QviQmJ24uyDTWxtgsPr277v7KrEHDwN44seZ92g+XC7vSI+eiGQXaRozeUIBGcSl
8aZCDEp8j3TYW2av1VJOjLsguWrJBvJeAjE3UYXtq6FFv0RcAVsZU8tBKqlcNFqj
Xas6ikDCElnVnEzwyxOhUIMoswYLyFm//V4xbENFbl28wcrIvOrbaFHLu0TSYoXp
RuK+vz5ya4sCU7PzQ1O/ACH3SaaKHBURQTJLSfO8GTE7dim9DKiVE8Io5M2qAGEI
Nwn4p/xcKxqGuAnWo7mGvSUN0h0sKXNpKatjE9niIPEnB+uBmUrGWunkPGBRrbyZ
FX4ua3nyYzM+cYF44bjNbDEfAX/mqVtNPUf9vhcJOTS82paH7WQ5j+byO1UJMIlF
I+JaB3VP2ND7gOqLFQ4+su/nZLMH0TOQ106OR4gFBP2kqAfrrKl0RZ8sX5WD9B3u
VTcXm4rJ4t2IVEXHztzvdjvEq9YaXpe2/eyyIIW4bx2AKfPB9KN4oeILTug7jZDH
STOORyYz5YjMT6/C73n204Ftgj0YF1yozZxK7nZFBBBpb2uMXHt/reizaUJy+MCz
hp5ysEf7+3+P2gCj2Rw10bp6gMZx9NIiAIVwuJ6MFlbEe7wP+48cY+xvExC7X8ss
hRdD3C0Mq5rQvMPWvRi6Td3uNsGKehhj1NrMijjmAKLcTBVw9S9UGba4TaQ2gtFw
XOHBX1NgM8YTsxEFLvTCHMYZkD1YuQjPc7sPP3ScOFM1MYDWyq7jOj6PCcsVEG6t
lMqvTrwDFM3QQWJDNORV6llHZKhAAoRSJV+H4X6VKg02mBZi4U9tWGDoWZnrruZy
6EgxrA8fsOOUt6Hg36oIxy+GYimpiZ3BIFX8FO1HP7rvtUL3WA9zpt79h+7Y/L3u
zzb81JlC/UbQS+44Df7A4KmLiIc27FBiBSITjDPvFvxtXBJlnrCMuLzQ9Mas8CK8
6IOIJZtG5Yra8685TM8BBZCyVl9mELC3IIH5yCundhtmdnUciiyRwk9txMIyDnap
aUQJpAo5R60kj0Xq+9rvGV+NeVmsU8tljontR5GSSayQrfon/E1QBUy7nHXY7A14
z51FAL99yDZ+hBMNUZNo+0CKpHK9n127IO4YzRR1YU0cXqibrkuAo7QRNuXgiLdE
e0LQg/fDsYeJ2O4jMPrUseD7XrLM9JwWbYm2KmigaWpJFTQHRhdB/Uorp+3vSpkK
ustUPC8AsZyMd1G5CDzuPoPoAjkAl5LVAf6ZZsGaRCzi6nc/PNKx2PJ7AWKeXawf
OjJvLgaZDwkF/GJHvzr3mlqRokK2Yml7cnIOoCIozX6HgJhQTi1FsJBaUZe74z73
3MuYlw3m/R1hn21kXrqfUCUmPjsEL/kIYVLcIVmkdXMWlsFItCp6FG0kERBhiuNZ
XF3b7O/44/y9YRqF98VoQASqeP3FtMjRm6H3iHwO1qc+E5kd2M2CunPJMl//amCC
jpHE4ZSKyYU80TQ5MECY5egHIWMUO7akAMGQH5GCmlakCWrdKrDPDA/QzU3zuIet
tNqZIH7Hi/+7sfc2MH4UCnOU7EMAArB53W1nk6QRXrq+71gqAIGV3eDnLcMMT0EU
TVkLZw84CifapYJoXZMwyhTceA7wRVy4deI0S0bNOEqDMe9/ttJdDw4EeMtzs8xq
UsKD9xEKq2RM1MaaleKvsQr6u3Ytmlca4SNXpL0RuvMBElYTaT4i4q4aWRDLNeTz
BoNcOTBvF168X5/4cgCNWuHWbXTXHuIafZXu8Xr0W0rvXgk88PrAU9xAupmssAMG
PaxfPz/sqtWFSKAlVFBvNKUIIMmSnb16pPQ54iLb/IOqTtrQXxmWD52ZdfADl+th
wNAEYahpy/PL7KC9PQlF9pS5nAQ7NMfzewWTZkpir+PFMyUBX03uBgM1h5Aflzdu
+kz4betJQXbsxx+Pjdr3MRN8gzAfJ1QONN85m+8nfI8KvszOHfGdFPffzfYWDlkj
5MvDfPyUDryh2++YRY60ZLKjH/RaicEO/7Yi8Y7uAEAdZEvLSFKfJ8Rmkx1Cg+gT
PNVjVdV+Tt0Ma4uQyYx+riX4GVgUGKguixikD5YWMbWU1S84s7hPiLWNX4QcP8dk
6ZU6WLggCjPZkt+5f9T8RTqzY75o1od/ozmD+ob/hODnqJw/vjhI5UMRSGOcyiAR
hUCEat6ukSznfZfYGM101qAxYXZVF39eZ1w06oEJD6qSOHIJ+RMDM84B6diDXfXB
JdNDhcMG82byMddLsZoZbhcfDXhN0BCrRfdZM4A0XJPZ4Rtp+oiyhQ6TolKM+C/l
q3mFYim2GePejjrxB5J+V2Sfmxk38gKd6uhk/l2SbjyY6MdaDo20FaF71viYLaZB
hrIA5uTrcTAyDJPa0J3LzPAGM1KNOoyJmUrBBY5sUfB4AeSfdqEoqtE+eQkjLbTp
zWMvLVYL+a2rKQs/0yJltNwcjM5MVK1GJzn5Lzo8eUjZIb2p0qRmYsWUmP/HxEfk
HsVbc3m9mLk5sdPDozukTQHqKa+Jh+5nQAXnVFrnorFBIgPd2X4cBqgDOMRd+qwo
O7dGb3bMMUKAC4ZWg/ZAjiIYqgjLNap78nYtnwWDbc/wLp7ip95rbvkSYW0TnKOy
UShabdOsSFWDp+DOiNZ26CfKCXiMBerdDfg2UPdbUu4u7FvxELuPL6JeivhoMqpd
EWvBuIrpGyCJC8z0rL12TFNg7Md3epitiUR6jB4bzvXTnYGRIDeuqeONiUtEksZP
8GxFESjXRij4U+srCg5TNEDm8fZMXQYCzIELFbSXK2fwielNfHB7l/ldaTITV/5M
qFbDmMLLZ3nDs7CSAO2OsLPKb3zYzGZrCPZc9OF0olOTEdty893m7UIrrN43mT8A
9wr7Fe4F5hMgLyNTpNSUSOEJ1G2qrohVWAPyDaKYnxfHeWbU9COaB19uFgeyfqt1
sR9BBtlcz/XiCslVGoIkFUxEGmcei6kGbc2d0jSafxbXmKfD3eXLsG0E+isFPn+Z
CSk2L8wr0CSGUFt1xR2GkX8Gy3or1WQL3nJhw5BOs1A0rVK1O7R/g60ffSBQFM4S
QzJ8mayiaFtxyHhANfR71jbDdzzugb3y6XLzMDnaF9tIGdkqdZdQUtwaSQcB397w
t+vt2sBWRpXL+pe539joO/Xdct1rM6aIpeL8cEUMlJ3nC3XHA9VaQzJPyl364U73
nP5XWeIKuKJeENb1CgvbMeZyfM4Iqfqrw+f5U4c67+lhZ4A3retjtsrXuHb7o4Dr
q1UJMUYzr5g/glpuzY+IFrcqHWL0DtGbE+LJf+BMn05GEV26VsDee/0aDdxgn34O
ygMVaB00+YTyhpFXNWEfKguu4sk76zH38oRAHc3mJNySKw0+wAb0jxNnNqS3VA5/
npz+EcF7GQx9RHowEO6TnboUXxFpn5/H1VVV0W3NKhFWdSmCJCnJoHjUgxwSs8V4
3Eb/h2XKxEfrmm9cwdNFf2EIRD7zvSUVhYyn1oIt66jHobL8dJj6CJYOagUQZkKf
53QFi5OlR46wxI0akDZOgVF7evpddGhNGDDqCzBwNIxOowYa/LqWeFp5t1jpLftm
IQRYdvYf/XXpWFhIEEeQdeFeeDoqUIOF1in4sq3pAh2ky8/4RphpJNCZNx0p0QLE
avB2bUAkXR5fzAtw3vwa0yQ/qrY+d/4HTXTQ/zk+PcG08t/HqOtlSeiLtPAlB4kx
cc/FAM1DP3teaCTCkuJ4o6rkddxQGKs8esJ6FoBBo3Oex0RUoJCxpnxgrMg/9T4W
b7jaLqOifn8oiB4ZAE6OAi/KSwJtmH6O6ytputH8y2U/ehJMZinZD4T6VTqNolKe
upxWEf+5XaNLNuSc+Ai3l43BqL1OQd1R47yKRRw1MPfITK/JRJFeV/EarxlCWJ5w
7VpeBd/J543gHoNkiw4hL37vj8zKsBUoaOhAV2uRVMY6xvZSNGCOkcZSxZWnT1MZ
Z06GccKdH4wrzL1CEX8tON4XyjulTKh6rceP7knDSnyCn/7C8j42tc+iP1CBfA+l
UACLO1RhPusIw0qV46iUVL0jYbOSsl86SnMIkc1T5W3JjQcB2mIN9UFQzBhyUpCW
gVm0QEwuBSlSCpTMTwXGyPn8RUqskJZJMwmyi6k93u8zU5kWsml/tyO3MRpDu/1l
FzXxk9JqJF5DOo1nUWWzkSmKHCfwYpzFJIM+e1/SKu9ZwH3qgJP76R541lWyiGQg
7AZKA/H84A00sGMgihUd+ybAY8QBWnyEdtYLDsb/aAR2InaYakY8GFETgIXWn1/b
8COnEvGImSZjO0BrG18IgujyyK46NwQHbBz7vDEPtWP1iDQ6n3JLvndE/O8l+qa4
yKW6DAg4QgNncHnxl998vD8A9usQ6mR3vAyuWfHV1wrzik6aaOAj+RPkjidT9Btq
S9M6Dhl2GWGrxbaEtwuqHr3eeBfbkFSTK8TlQ8FqJRFcQDxVp8cEMwJ9oyxWG4P7
NmH132mCGSDtCTtmW+m/8MB2ZkIXGfWaXxgPuVApMem5gqgsN9zvVApdhBLmsSX4
8s7gAKKox5gm5Z9hTYyQj/mPVn9xtKDONOOBTX5wZ/1EwJiqRtK3+fEMAiGH/gkw
30DJSGqSok6QX1BL4KgSn8w5P+UYnqgUVxaMysbUqDHLlq5sw9X+qqOeSwONGPG1
o8vCbqbeaEzoYnnBSjOKkWQYPfvzRpg0LmfwhmjdSOBIpmWVRwDJLEAlbEqt/hbs
A972xr+brorrLQmAFjGeIiXp+iPQSTLs5zCG+YO8fxJ2tkRzVUxqjqe3hZeK2VNE
vgce/nQIyt4ab16SgXcDuXi1R3HeTC5KwAF1/K2rHmAo62beV/CsCNPhqHAdkC5E
YO7SWtl9tNxdxCzZ2V3JafTS/6LDxOp81oBKTdiXQ6uvpRJm7nEropouK5AlBQ2X
YPlyM/EfLANPXnfxZ0nbmc4zFu6ums95AQqCqh1uRuda4MuIrNgMySmlpGoXcDEZ
1XXJ/UjHhNTqU1oFsaWxMHJclNc2Oa6SOQIC6fkAp7NNAD6fChPOl6sUI2WqLDbI
i9MgZrnGd/MgaC99uPSjC2q+r1QUdd3Hlx/bhpE8Lk7dkI1jTuBB50yc0gjS4J58
za9iUu4LfnTBxcZS2iwQRefiiV9MB68eJfwgrhp5Q2Ldk2hT41dEV/eQbYJ75rzG
N7TVZeQgtC9G2L5Ywc4e5IAv69GlrjtxBJwCSUYEHhoXUySW/qHdgW+4tdHtbNUV
PvMZkBkdIwi5i5uDGIIbfUrklA0uPg52/JA12Z93N4QipgBIWlFwSW6M+3NTr9LA
FAxlyGaPyacjcJ3tf2+LuEXR57LyA8/uaJ/ETgnksoPwI1qne1BmvVWwlq2HN6Pf
aHUXS4dAYdOUXtWnmeQXGAk+x0bdllJIgB+4Oc2IUH5jeLVGXL5AXOn532QO1SJs
RaHOhLtcZi+UqpWITv3ClMGTZAdEdG+pJK7xZSmk9wlGmixBQeNIqQ9siWcnmoVc
iKbSZMtcXRHfHfYpGlrBopQHUHdr8qhP7Bj4DJ8aknFrZvZDx4uvOfiMp1Zg9jH9
KkTzJlzyUc70mo/IJBDfjs/NGBUFKS/T2XDC0WPwh7eS4cJeOnbK9gTziTIq4Fog
1JNzxfGnQjdh01WakZipGDtAr/DmzJFeUKsvWZfgmedNhU0mAQpHpXSIG4yQCCu1
Yo57+O5rLw+8/XSz5ip9pPJYSvrVmzfpd7vKFqhMIRqDBNWKpzEoqlEg/7JFkVT4
Dnfn/cIHM1i0RGy6LfGlXj6J0t6jMqNM+gtdSUgTXg7TMR9JmPX+odEZiF5Djn3X
Jr8SaKvbx0TgOfLw0EbC+tUVATpdSp19wTTmBJEG2U4OZLFj47tc9EdVVDpVZhKb
nczEdJaABzYTGlLkl+hMPba1G9xjlvlh+Gk5axZCNOuMeHZSSYDW+L513fxey+c9
84IMIC8STGBhGIUAOoOjb7xOT6nKhOJwYKF10yj9/sT5a9Kp5aixb5pC6uqsIOBu
VOznIXbk2DCcMY+EJBaYtadLFtSvY75TTQsM2v5itsjg53DgePfqidHQ1SRFEhuo
X/Fsi/mxTg1f0PkTZl/Cx1Ft6kThVZiWlDKM4SJY4FNwtod9UmamGwikpehQbIU3
OSuEjEVFqdq+mXOGJL5vMzqfOQ7nvedN8ry8FzBpxASjaE3wPnE8lF4vkxzcBy5P
9t5Jd8A8cZTN4yFq/beVB8dw8uGSkVSIUvdJTHKSuvhu0WfY7ysIHJpBA2s653FY
nm3C7eGgGR18JfjbdOR4ypM2tuuK/gffSq01KOZWBupsxF7l5ZV65R/o/p3LRMiK
dRHSuF80X1S60xmPr+kz70kdxy8Zvu4z+1EDZb12auT3QNtlyOkaKdU68YqLBEd3
8CnbHIU/gy5fXsKvLP2YSqXmadG07uXQCFW3Sw5beQs5+TAAOhoUlk2s5e0IZhQc
GoFa0RRHzGfTxsNHt9RONojkjm1APPey9rn/p5rO5H3pvd/KOVZ91n8x3axw4/5H
MEcIGyvhOyKNmN3aV+FevNT3q9pTOLvP8SXznyTTwJ+4kSw0gUx3LdGGwS7TZCko
8JlVf0xGw2t0kBQMlkXj2GJ0MtKjftdeF8BEi6HIuIJUB8si52oKezVs64NCSZKq
7aVOQZTpM74vMa5FeVNVs2C23mD5w7XNaMkbdupA9YSX5UEgiCd0O76JZxYqCVly
Gmkg98pFvvsUlbR+vn/rgGyUjmCIvj50WkVbMwIBiXZFwIAgnDwQAQYbc4qp4UR9
jwB0VF2yguE4aZbKRjXgKy/Wg5WmqaG7siqlg1+Pwyv+5kPiMDAFmhYgGdhKdc9a
EMELL2dfretc2UChFtqY92GNyNApGrU0euB1SA/bsqrX9oWCJKZxw+e17+CTXAXX
62YeSuvsctampgXlCuI9z0x3pHG/HJ9ykFiaGDVyTeLqDUtUvbM2HpQkwayV4NB6
N/jXunc2yDVKw0G6ujoPmTwOQajNw7tzC0hefzVepXH5DxYw0eUgJA4X3UF7rUfg
Zh5mHKkEemIoBBGt/aSNlchvhCF5+f30WbWyOfgU4LTHKW/uhe4wN4M3WjCCBqxW
DtUx4rIksD8i/fhEcHV0h7vxd/mrtyF9ys9n9JhcMwBIfj/yjdLKPv1OmyR1VTXZ
/L4aWjnt5Uw+CUQ7FPbZT4H8SHmt3gyS8dZ0AbGQxkmsgBF9/uAjFuhkKfX2foZU
Mj53Rb+0pmSvvxM7Kd8f466p+erzzK6oZzxJuW1CHLda48wuBJZb8p+DyIEIHyoo
97tMh2JhHKaSuB4nQwXVq0t0PBiiB76SRNqgHtAckpLk4tJW9oQCehHduDcoxq2g
0u4XGBnx8W8YYYl/YEzhq5ZFd+mJSUVZLmKvaljx8Zocv7Ydhk2v8vVgONgXEf/I
AeoCy7lziwRpJOqRhlmSQ3OE9yBv2RL0wWe00w+/W6PKopr1qEgxDjcHgUz3NFMB
RuYNvPZ7G6QqNpzd8xOk8mdyqELeBCVSXuyoDscnnN/ON/ErFrJSXr4BRcEEGeHn
3e8aRvtZVX/RTM6emSFLvQiBwk2I/RrgTI4xdNlM8liKUOxLurQv8wMZ61ABi3SE
eDVF1hgRWEDwWbIzUvNi2Pe7MYVpa5iEUGrrD+4D0D/lnws/jre8skGbZ1wfaPIp
rQczXZzPrXmocKtsoIS7TEQvtHm7Alc1xDW+HTCkRXU9BhD1u5wRvhtnaN8+aYOd
ovAiJyAAjhtSlXRBN0gWS89zQMjEe0Dky45WlAjRmvkYvAQ11YYEq3aPvV8hMZjJ
Fu5nmM7eoIgnChCwhAaSlFS5fCPQLM1yz3YViWpGefcxBZcviL1DzczB68RjNXE9
Qfdgy8cvSgH4Fxtb9FA4fvrDH7XmJ3wiVtQFtJOJ2Esv08FImT8pY8MOv/zLd1+5
YNGEHL7xr/2yN7XZPqU174OWk7ct4Q2thSrO9HmC0l95bEiq7rnbVqLwbV0KuShW
CNU7h7PXLUzYCNwqI1Id3OefbHR133FK29KXDeasMscDr/JUhNxDJIsm99md7zdc
It081Scs2tbQ0ncwKhS8HAGvXgsOLBJmAgXCv7me8OUFLMQ91tUsf9PDzbm/HQq3
W7Yc6nPS7fowlnmyXLu7/YtkKxd/I76odKmmJvstrFunRtp4ecerJHHAllFLTJjC
uIENJkj1cTraxadEHcd3vWDc6PvTMiLNLgTMNaSjE1tVnXcFzF0vTxpLoHz357xv
kLdfKeZdd/icbEOrFyddSrOjCjZDb+3gA91HDBJA8XUdkZXLvexBxpDFrO7/wUt3
M6ttb6xs0BNuRo/UlPUtcLpLoqIDTc5laKHlMn6zl62ntl98c4QfxTthjPGtO78T
ollp01i6WL3tsod0q8Yg8aIdnDaDpaQrgUXVVpJ2OiL7DMUdY3+qPKQAl2S9y0u9
zb3gcmZlbJ3JERJZlow0DmoIHQ4KrFalDXN2tyh/3s9W17Fr0pKelC8ElD6OQ6Km
ykr/U5oQKs9KdGU3Q+i56OIfquqXk48MDXf7YMtcuELN9ujEenWWRHS02Ur3oyf2
BK6U6EskT8Su1fsj2QQXxcZpmCf9aMpaSgndwOn9kAgnxXO3hQt6g/wg6Q1gxBQf
XUajnmqXp2V4YoPtfMeZb6uhrJFX12M38//UIwPui+z73Zx6sLNv2v96zCz4hMDJ
0ND78m/I3lgOAETLWTc7MUdAeI4oGqhHGcLkzeNM6NyiSDINCadCN9DU5hjnY8qR
5iAd3/41w6CMMNixxeTVAISGXeyLpVs0/C4dR+ooiK89LIvu6/T8YhWrQ/+EJAoV
EwkD/SW4ifOvd2Z0OlWW1KJgx9l80TioxJ78M6/QT+XYOn8qX5fNXgFV6fCyCYns
oGB9+JBG50RdwwT09x5Qr4gUKdKsg5CjHS4fop925tQRivQTMNO0+VPFwaCi3FAC
Yi1jxVYTlNXhBEuadJGrcQhamqR26IiZpXLGN/kBw5qhvlTL5++49W6MYBuHGqD/
AQMs2pzzl5KJpp0F7DtWTDha8XRrXINkiNqPBfdWLLbU6W73x9ZtVeOzm1smLrVx
4DLStOf4jv7Gdcz1woTq0voh/CsqmFCqoHWKpyUioI/UYdP5zqd68DNt7WN6T6mR
IOFxt5CBMMurWL4Cc4uk3w77AS9zaH8QYUtcVl7CzvijjJnD9SdnLsV1fSbj5TZx
yt0TuIFVcnMB7M9DktLsZ4ugS/zuwXsMwEXMJ2h5RNDp8fj9O3lrfKWmuugAtqLi
EGg40s6vrarTg1TDcyFOfnspPZbvqT8SjD99NcPJc4XDV+gIxwrFhyJvOJ3LGAN6
TcF5SqkVvnzOTOPVsZQbhck60mcaVjI3nAgUFeHloqlZFVHC4hC1mXs9UV0NDIH9
Ws5YXQQCJk5RxcX8Kh+1bhMPZp1njc23f7HwNqqQrCpWhPZ3rjYifcafOJ1SoaXl
/7MIJS9KEU1v9+CHrHrtFPQeSUBUO/f185Z9dChV+rQVcEg8v7IigWnLW38XbdP/
WNVDgdaugjC0YHXjT5uQb0yicWrkPiFw/1BGVnrpiifhBnBc4E/NHCr8nulSE/YX
d88FtFazpYVhlSG1dtj3a6/LzoZ+fc00ghEN4xPN1s+PMH0CnIFjoeHtuCkO1a4k
PRzOkQ8tzN5zrNjsZcNI+FmLTlXbcKFI7sC50H9Db9pXzJLyp+9fjFov6LAu1ob+
h+26t0IIYXW9b6UqXQM1eJmZ1o/ez1NwQWnh2vcdBhsIEJ9kbxW1UnR1yxgv60/8
2HlW5h2glK1ESl9Vd4EBR/3Sk3ZSmzzpuwrY9LpjByS2+V2G6U42QcgGzdUgZges
+Iw+nu+lxNfn+x/uigl4bCTheDUwCU8DIbisUy4U1rNFD3cwKLWxDoNCnjZ3pT3v
vkzDyU3evs0dVibcFuC8seYtH/5QpjPxIUaMe1RetgR4k862u3NcP2ZVNvdmOFIx
sd05CLgEnjWGcLq595K4T7bvNkz7oslasjXm80O7wHZDKHxqSe0X+OvPu/e7Mj4B
KeO3p674iZ//yQokME0miXKmuzKF3ANaXD/ywBZ+mNyDEswkqwBPOCt0hoA0CLv0
NbH9aQlLRkiQuir+MLjKPuT2O09qsWW4pcV5V9DIBM5rgqws7wepAECGCPRQ/rE+
icBaxghLLlwEZI24s78nViZY6zklOijzThxyR+/kf5uIgY+WXhhUkobrLTa74SfL
cTY6Vt6OghlcFCEwE83yPsy8/3FulcLfnuMC0hktTsfkRLhtVp5Xy69xCIUpnenP
9DXyccXm00qpnG5/4HMGTlGMyIjwOOBg8UOOJTXy09i/Hd1j+lNKBx+/45kkE8MG
vHmuTrf/T6HuwXtPC1qH3Uuj1iqG65RsaHLFG3j1YIDJqMRMpkjwta8IoyxOODid
YpBtvtdQLh68i2vNK38RZG0kPxgataOB8s5MLobfapWK51QhZALcUdqfJAc5nQ1z
KSdSJYjHkANIEJU6oPGjjWPXKcglE8OjF/k8f6+S1oc5K9LJk5xo/kMYuEFCDMsm
UAXtnQap01p5RwVC87auH97jVx4KMUkUzjAQbzvXu5GkENlZLF+3syagaJFUP58w
Uz2+VUg2LwrA22hteyN72oo3HyE2l5OVJZHXGKK/I4SZrwr7s0UU0HSkWsZWbGkK
ZnecGk5ka4dcqKN3vHW0EfWuWzBkSdo4lLYULRWO97CTU34ouvnSG375kD9RMW11
9bIhzvlErdd+X2urltTRog16LIwKXGI6Pp5AgdTG0TpWQWabINWospMfCEgWNcp+
uXann+ZRtu/2ZWts3UPJKFxHwut/3ePPb3s8oKBYVa6wdQaE5cGIAILxd49MCOOi
WO8Hdc/L1sYbGv3viGGNHG/IeQln4GGrEaAyuF7NDWLGaiy9ypV0PiGId5n3NlQW
U1lylkjH53zXNQyOOz9DTpGS5XqVS+psXY3uWWu7HpPMHHPAGdj120zBVJfBICNH
bQlODE58JzStQynjRgmNsU0rqH2RvHmnPl4GWK77eHuj4sj0hByJ6FfrEHrkoYNd
EQGThCfEsaLReAkUm7A3Or2uCkkJzNBss41shm0VCjQWO6Y8QWeS1RvNBwJc7vXO
zniMI3pFEUWxKLiElPoT+D0ewZdYnFREkj5Ufe/oXf3Mwa8Y87jDX+oTNMKuz14s
hn0G7z3FmUtGtpnRzozYH7bCND6e2Z9BGHSKwbJZUZVjJuPxorq63kxzMiy/LNI3
OUN021qgjRLVX9R5hBQAlJmHZM2ywZSQusVubywuduP2YE8e+KhmDhhthoGxbr7F
WEqg32ZKXsl6kOvb2MUiUJ5mnwrtWfVybinp+ZxS5RpL3w5BKsSFDQDVELecTiv9
pNFUxYJnGIP6QHYFfitDzKfL0Jd50eCPNmiTU2w9/XZvioQbldECmCWV+XXy2oi5
YMr7fAYgFzDYaKTZZH8njs+exow3Jw7RjJIlW8rZwb7WkzQ/MWO/ir0RfhBxY79X
fmG0Og4s/ovpPq8GNgB9uitqsFqVTjJHPpd/paSmCV4ilFhoakHXmTy9GILDMqa2
abcXYw4/Vd5MNaJb7/4D9s1InITzRM7KHdwqA03K5nYQu3GvbELl6DKKLtR9/OvE
Pm7abdx+7lWa11YnO+8goFwJ5Xxn97Ts2ST42Blz1Wg53bT0NHOFmQTH8jA2mnYB
fW0jPMU7HOy8/I65Pd8aaMQF4DuhQthmY+LEDNrpmahVbqKIDQCid3W7d2Xhd8Zh
n2Sw7ak5gLaLcdAJokTUIVXWhFLx1v/9tfh23KD53Mj+hn3lBe96OZfEdprrBJuO
q5Hl4CFfXOGqCOdGB+oRwQZtYI6862lO7i9XoSafw7mO8S3nf/jKoqRgASDEMHge
gyT1FEzCVS/51u8I7vmZPjjlCGmq42Rjn5E1HJ0El/fndjLYlzyXB1PTKR6AFK/O
IYegjACxsFM2/Hh1FHn3nCcq6Yios64pvAYo71m8SZB2SPN0sUyvdVkCayykgCIp
nMRcJ7he8qt06MRC7EiRwDt5RXXK+0HQAlscB7QcpOAnRC7lQVfuwM4SiaKt4Joj
x7PlrX3boNiTDSG9PSivlNGNUMWdJ7adZVOVaydsFmILcbWuFsvWnfWutXrPpjza
VHP5BjUQreu4Vcn1nuAm95s4EJWSWlaAqHi3dIGyFZVLQ7Q7qRkYk4vHMoEfJEUp
AJLFzDDvIXH48iNinEVBN4NupKvd/R/xLP0QFWU2gcccG72O6hnGtRdh786XiGcq
nZyF0VbrQTtTqv1qiVms49MIMr2Yc6j14mtz+kG8FFE8EsZAOf8r//fODut+F1JK
dJIxXfA54kv+TaxDUMsCpYjCkurJlIx0x3J4yKNkxAhKJvRnpwpbYw8Hvnbs9j+l
TvPekpd9nS1ha1hf55jvuhHdZ3UUd57muMioow2M7rbx/MQwRPdBMiQ1fPT3y3Yp
Ojgjkvu+ggMbXYFEWasUXbakCnNnKUXD2pJ3YpjJIW9Z8qf8w7kXfrz1JfOdHnQx
BNZ/TAixrgnJfm8B0Hy6/giw2Dh8Ch1S7xzJsYy9oefjG6c6/AuB2GfyOOPdIuqM
4fmCfet4oJB2/ZhH2mevlKq0w2vR0IcirpG9KEOTJskXs/0dTLp3heW6cXwrpWU8
Sv6Wp62m913EzQ0AoyOxK7GdkTXM6UzO1KuWu8E1sJR2BGMntq00Qd+Im3+xzkT3
HwNL5KiYhD8Me5UEMBigVZ9EzBcrARwt8qTti8GTHVgARjbqtsAqTJo/FfhKl+VS
V0gxAhs2xkkb313W/Fc7wubqLC9KPK5witopwthYFPwOhl3h+43WMtf7AYRWMOPY
rpCcY3GpihDl2skI9Cokz28+i8mwM+q8cfrzi97w13E9POioT4O36Mpz9l3R9KS3
liMogcGgqTjWXNhaY74Rzh+Cg50TmZ/hITcyhZeW4zppUcw717qjiqpmC3QCRG2m
YxFqah1puVJwyB/i7fIpyrtIch/cx2iLdXnO+xxLffJ2rNz2AO7NVx+6mZyxfvu5
iJpea3hXn77+fioVSo6j0fKu7B2gbJtRGd2Fy/kvJYtu3g3cKXSVMDMCRzdwuqwn
uORXTRk1WKzAz1R46SLjZuc4POi33YaM4up5LfN+7x1yOkSCWudVRkZd/IuUuLZx
hVlwtsCbm09MaqMv30iANb8sLhx8x7ugqR+ydr38OZvj3gaUjR7h2Jxjs1xJgEYx
FzLCsil8vsE2w5iP0fn0vW2oxjUnt+R98xTNRhDsXd7X8LFImvb27M/3NW/pKqtg
cS3C0uG6CIgiRTud7ayDEZMRuAPzQ0oPysE664hbcFfLrYh11nexhVq4BmOjTU5Z
hueIdnGYTyrFgunTPoRnEwA5B45vlaxp2nn7THvWsbPt3qpWDFukbYtJy0/f0tHM
0ftlOLoWwA6Uet6ynam4Y51nw4TA6HumLGW/s7fYc7Ac3iP0sGTQX7OwTTKmVtjM
0TMZkPCri/mOf9vEle9c+fADBKPnOSp2cTu7rEz9nK3F7yVzcZIzZUd8JxmweIDj
nA6w36XKmriuj0Ll4fh3UgOrOBC1WpMKYy0Eeimxip2LU/PNMY76j0Uegt912i99
o00+r9t3xbDAvdsNMhYd9dLoRW3VR9fNxZ3/XKI6WU1TCpc6RBagLc76Z4dyz0iD
C5f3Wl+M3Et48qbaCvj1613lZ4QKEedqAK1JPd+l3G2vnsjiKnFdtlZpyaKEohT+
V65D7qIutHT3tjlSD3WWJ0Fwdv9VKvO1CnmqzUvZa/Q0Z4jJqoaVBqDXbDgMXITZ
1rq0q8KYwBwEMLOGWctT0QSgKbKnSNHolyXnTrrLlAo36iW1JEz53IemFLihhIwG
s9Z3WEcG+bUSEz5rxw/43RBDDN294JQGyEnFtvlFTx7UY9TZEXFZIB7nFyWztg1o
MdLtfV4QaDD04V997u/RV9kkKwU6/umTmTQFhJ3TpjuB3qwMri4GHdAkXN4JAEEy
gE2Tv83Lzu4O2VT+8jPFfRu3ve+z0wDKfhUTq10de/7Pyje3Q5vfjP5bJNwo0bIL
WUeZVm8OdgkxEC5nwDto1kilWZQ7r1t6oKLVzdKaocobU/hv+ws7EhPzLxqQU0eu
KuffNsEzYkK3nWOIP1OuGxxRZE89Us01FFXr6IKy5JGMs+bO7g/+hvWhFPXNJO5s
owYNbkbLKk5hJfdh6HCphduS5xcvauzZMdTDv5gh13gjlVC3p4fAWEXKsw3G8zJk
Z4WQBF4qKQzeYyVTucZIGnmRUGnUYzcyHAVvu8rBWosAwe/jTcNFBW+CubSbH10S
wag4G/6M5hT4rPN2gajn7IRlTvKm+v/SVdrKR6NKTNsBB7iijDKOnZSKCXLRLTP9
zPLz4mO054rA6F3OO6tIIEsii/VVJ59dKqGHxYH6NdxL0/yneGVaIX1JpaAg36mN
FOcGdVX3RW+TArqMDfjUW1LcUDv6Z9SfKbe95Kj21vqWyfB7uInvvX9gTFpBO4D5
nYQhdBIwlYa0mB8iUohi9rDKWoYDMfwNSbROvf0IndCYyyqxs5ZITDw49Ph5s/JU
9pmQ1XvNZPVPLDMY1OyNtGvPHEdS86PmNhn298D9LzkwgURBAcoC6xlmgE78P4fm
vih5SSb93S+gW1T2Ssv8fUykKc38yZlzAQ2dHCfAdkvFsDTaeo6qFIpQXBdTSNK1
Pi982WHuNc1e+ec61dLBA5Yk+li0jxXIEly82JRrz8J59zuNzHm+N7+b6dOHgMZd
FMCRGdSrQPhV4KfZlge3iivnV9KGtci/sBpw7tL45aH0t8JlhrfMYZtSFIE2IvSW
V0vecw4hLaKKM0xT3VzdH4pVYQ8VuXp9SA5pBSHa/5bzsmPDoh0vHPpVCI8mcWSI
J3PaXd70WEDba4qLiZN6gdo7q83d+HmP12n4DbkD20E93Tsgk9thwF/QGIFbnPxD
/nWmleNC6bPqjKNfPieyzhZFadlH0DvG7KJEnHAC4z927n1HHWPnxTXvG+OHL/ef
4+hXJt147npB0Ml+Mc12zG4CSdYrLn06pgl2M3Y8pUrWAM2sGGdoLz7YrfINiFpn
7+TcLRiNkv9XF/CGby5ZQwNW62sjxVs3H4twuSqrum4r15wMqq2dK7ET+w7yAm3F
OhXVseQtAFRyWNXYrly48mZn3tpJaNTiU8jLpofIcOpzYAyOMlqcXxghnULHd7Iu
CwLoJr3mL8/CAwVzE0QLICgTP/9ftlUhjxyJA4hWggHJFpWPjTOab6HfiwfDpGAe
IGMkpZoQktdaZbqFFUOVKQGOEsis00haq2zfD2/F65SktsFz0fNC6+h+RiaZS8tJ
OPg3UWdy2XrS9t2f+zplsmJeGut4dIxouZ+PxzMoFGPCbi192rdPrkPN8nxG/E4X
Qn/F8MmhxxFKJHLnRczvx07qUjq67rmsg8s0zVwgPuJucWZVmfGhvRd2XyidQQRh
7N49xaQifEV1oOsB9v7/csUzHBBKHahltJ0cCDNi99MGXHDxnIDm3J1sL5QOQUkm
sl/0Wd4FxxqtxpaPYOq0OQGqR15AKdW63bjO2vxdsbFKZQCqKVAUCeTUQvSMgAhq
KugXF7BbtIf4i//JzaZoTInzkdbbojR72oXDMgq+Lc/vb0ALfmDj5ZW/yyKJFpmP
DMMontJJJZ6xtKX8VtdZFOvZ8RhgcOs6GlibhXpI+RId7mdVlB4dAYbO9HT4jDfS
sDFc8v9WDa01dRdk3LZqVp97CP8drh2ErMvcVRsBzrs2naD+ACwplF020lR1pgr5
2y4Oz04H59e89hcKtL3TA9mNaL6yTSXWuq9iGKK0G4uofAsGJqttpOEow5ucVbmp
ezyD9vRU8ErNxJqFLZqiS0fEzy1FYZOfjpHlakAeadrjD7avlqL2fa+eX58NfrA3
qgpJ0KEu5HzO56XAdxhB6qGhVNvciHAleP7XU1p8rH3f1knuEHqKBnp4SmWpjbxn
Se+EvefxSxNROHXleJ30kjlGSTH/+HkXLWl/9U7NytNSTKdDH62hLKOOytKNhjuw
xbQJdieXnm0XkZspqjBDYIJvImzpQh6VfvJ/caX+Xv6AXJs3ntNyyJpKAZe+SqPR
3IodhhKSo2AEk6zFvdT0EyeT0TOMVsDMc1YVynmkZIvzUGg0AD1/ApuLvbw4AD/I
NjaE3pPvdWJNHZSCiyQAC2AlAKvQHJg7D7kHL6g+xwTJPCgAx0W3PrKeHNEVm1Pt
tKcyGPTnJHurgbb92L5ED9ZuqCXNBZESG0xx6Z74CatnAzhHZm0MGGrOkbbCi/rr
Yz2xP0r4SVd5yhioh3kUZ3P4QT3Dq6bQX/XIpJCBMyc0/JkkvxVa2Z2xhtuu8ZUe
oLJsUyvoHnCv0sLb1fCzXi8lja/Im7H3gT44sC0lIN6CS+Wclibh53sFb4ybxb1i
kTArRX2JDtpyFFSPbE3on0Qqfk4wJpVMI26eKjFkqYMqra+IAbEQddgux2/SE3kZ
n49NhoZNJZdVteFzN7NfzJVqyz9gEIYFbSXiE8VUuNTMeIcLSRgDaxQDAnte2jDt
p9OW2THv76kvXE+HxRlHdwCVQndLbG6tgNHTW9tIsCgzthYCm5NJAV9aChiPysf/
68NSeja/Sqwqrtr5y97TczzLHm+pBAdgE0rEYqs4llPZiuh93o8ZnA8e1iaMGCCx
NFjtZPAzGDaQFx0ru0+N3upBf95a0OsQh6SyUn14KEKwqlSnDLqa3kRuUhIKEZhV
1aVP9XJNM9oWQAkNdweyjjH64SpU8u8Xohq7RuDyVI4SrDSNedC755LQ8nc9JOE+
3qPbSteMWrTMiLaS9jmogGJzE/twMhggoQua7xWQmIZCR5Y2ySokz/0+svg2lba9
qayDigmL1/MO0ZqO+wvsSNqBPXzx3+YExSYmqyKqmrMRpsMC09lmRRQciXXZLC6Z
py3+SVNDURoh1zv41mZt5BhdcHTsYOMK9RR3/1JnjIh1wlcBOIt992bYU6Uwh26k
IqwIpEoilaxr7gJDz4B7flSrhbmh529Kc5hWzTvj8EjznLopryftgMeICFhwUVMG
1FB4RdAC4TGNk31ugbR9J+7H7Y+hQX1Wua11WsLZ0QvHmy3s0amj8LsJGss5bJAY
dfvxNON7fXn00DgrUpezrbFi6pCGkREV2mrle4aveZweLm0Kcw04MXXlzNpcK8Fn
BudEBdte4lAO2AEWGV8OinS0Fk8RhJXg4fHJaj92s4XZ+UW456GeNLcy9+XbeJlb
jEDmp/6qr44PvfXrVcSbWtI8DNCO4+ptORS6P3T/nDPFbrnrL4XOvjcLNbeqkWm1
V7Dt9pv9ojSGfGFf77/MVCKmk+Tr6MJloyHaCqDivWr+Nvdvd5FVCXYLid/96Vyn
nJtPWmEzLAF6caieJEDFCMVOnsWHm8aMg+R1bNpr8pfXe0x6u0ZoS4eXmjOdRiog
jXhY1fnKwAu+anbDiLfOHbqLqg4jvH0uDYkcydiqD44H272HkH6PrrYAxzwB+AtS
HjG+UlF3L520nf26ba9wnwb+coraRPZb16hvZXSyTvOVhwShN4V2sz9q1jXbtkgj
pCPTezLNIoceBBpKoiU3e+fiTTfpmzC1Yk1y8vn1ZtpXHeLYUr8ZE9/j37UVL5/y
n/k5/ndAbZoRtIum/I6g9B/lKkv5AHJ6TIBfO+xcp3l08eUy3AjOOWR6J7FqsDGH
nxTmQMFxBjRTP/g2FsR7ANKe3IXrxpKLSdTqrQF0F06wwbyVKMTkpVOg3BxqTIiN
9R/ihSMDOtCGkdiVoDmOiSaBSAj3DHwHE5s/1kd6F4xFQikUjL7VpJCIhJllGqmZ
J6AX2juMO31QMZkL7ufd/RHkQvPqhQ4B1HhFWu3PiQ8+HGmwx4snWkYjivBAjQYL
nna61/wLFZPkN3qH/gLmJ8lZwvXY4dIIWCVCq1irdHfsfQXLVbvvtjuN7ruBSPFL
4QOcfFUyqdbevvsTGLDgqBRg4JN/WcT9y115IGL2ue6U78EtghylCxGicGTBIs7P
CcIuiZ455aGJl4/SsKXMII3tNhvdWAkWFiWAoYaR6fyOJSCe0CxOS/8BFKIMANcX
uQx2RiIfy/ndiP1hlTUASQoMzJ9v8ZjkTRKK1rcDEfq66vszAfGSmuI6qTNFu+d/
HruWQJRfWO4XZRyDmvSF4VnkIFXCEgDJBJEG3r3ZZ905jS0aaNsir+yYAy/6eIel
SSoM/GyHbRe28EzlFna8aKKV2JKMLPtJxXFMQNTeq3LjXx30CoXXVolbqBIwkYJ6
to8V0ItKx/DF/f1/VcB0KDS4pnIVHldWM1ZhoJ1nMjxrsEy4mTz4AG0k8DUhAbVf
x9iq0dv6vWNo1c8bYAm927o5wHKO8rELWJh/wIjQBLHQEYbKnXui1Kuv19XrgREk
ZQQOsW8RNg0ArrEjOsSwZ5QpbyROXDvY197guPALvNe5oFy8rgdWBfBGkLQNKCBE
gcjaek6eFK9jhON1wWxVU1lzTXjcUExOYf5t6YjVu5Jwj4BSSKvDph3FpzHIiQi2
qgQkZmlF52YjbN+U4ZEhFNNtM7t1qXowNLuMqiPFmoLUgjL9tWqKvj9knK90qw0e
HP2ARqhDnJM+vr9EWN03j2RC8e850bCKsjh9JlhTBF5fJiseiNdpKYXt9Rksd6r3
giYYxCf2sJrSXvZyMt/uQoRTi0hLvm1X7SubwnAyZUu2/Kfpd3ZBht7KCfWXE/Kx
qrfW7spSxSYS14XzlrNYFevGZ2UBon/wSz/tj1qoJSlDhIlOrwWiGtfMNM0c5ZdF
IKAEC+7JqL66LCYCbKGOQ22rst+s+yV8ZdtL3Ljy8m6fXhCYgTuRG8Mv2QEC0+45
5e1c/hPZScpXrwecLsw8iYoO1kIZA3moYJJJ6PhUGpuQ0jPCFZ91sE20cm28BSza
zQUowoIjP0FY7dN9kyA0aOHdilfQCWzZj+9vm871KVwgslsLfIKlzenY6rG27Yrf
0vKyvQ4S2pFOJFaViQiQoZ74tIQh8LerOuHPk3T0VdxUOXepJNiYZ+Kz0mF6FXW8
PXIx0u1++FSV79OFBI6Yk/JKy5cVkzRV9Sfirbkd5gvcydSYdT0UqlhI6ppmEZiS
gyf3zDpPWwBm3AIp6H8tY90NGSy0TiVO6z/MTwhNQf2RCCYRVyyNZlFnD9MVqthc
zUaDdvogYl3gJwl4LGJ5K15R3/GMeclJlpyXZ/GlhJiTvUlKvqZ2WferOc3Kpqvs
1BVWV+UCKHGgSR8pG/uGVYmDjTPeCLc1kRCeW2lAZWG9oUpFxjHKNqrPuz+vSrBG
2zzuwFestqH2t0VMdCeaZdM9o/+HDdYP1nYqMWR3QP72iyvhd8lE1jevhswkT2x3
w7vYHvp32bK6kzB9e8a9NR5HAEY8eFBi/y4tohJjP4+AxXZnwbR5q4oWPM3dwhR6
FGw5nizDTAu/r4MU3xn8DXgIl+YExc04ZmAK6ExbFn+DSIjTtIHeDjFifEyRX8jq
5UKYLTUFBv/9kIzSUgDzEyyC+agzSQdiRCl4pD5Go1/N9r12u47uGaxOLpJzcAbZ
0qo6waFvjHoggrWJD8WaVz/ycSKNUnJrPSSzvYQkwXKhWAnhPKBDG/1f0j/+4vPl
XWG3roEGe0npVb2nIFIpORUWdTjP6Fz1aCKzTEaGJRcVKIFDkABwgTBPeRmsW70J
P+CffqpYONrWLN+Ntoq+vZWP0s6PnSkpxYT0TRiUE17VLIPzUFMzwSZWxtfauwoB
udTi7wAZpbZq2rc9utQ9v10m842DurvBuBa61rjBaNTB3dFth0XvWSM2gbp6NfMJ
X+cDqoGmoNaPJ+/5EngFqaDwBuZ0EgS/30nQvb1k2HivvGrNwf9/DnA+X4Z1QxTG
LAcM4NZh+AwOv+yS2CNMAdOFnKl1unA0H/f8es0nkUeDcrs1Q2Ebv0ngtl6mh6jT
9Su4pnYevjuwctox1HCperwyGUbKss3dSbxvbF/suDMDdfxsO/gWrd+Nzb8NOm4g
ILB3MDY7NBJsjoVirwZAQd5oJ7/p2657LaPdUhT072YYXIGDPWvb4Ik/9dNirVVy
t2rBlS5hDyoL0uwF7vtFIbYcvvRFlV9vR5DMDjHOLpIz/IWMvesnd4vvOdiNFA9K
Wj9rIsrX2RKUdwEy9MkXSwCPdWlKbx3D0NRo1S9IQuB/OrNrI3qmZVbkYdsCiT9V
/iQGP1j97wmT0kgtEss+TDpwlZlE5oIJsuWUIuaEOQYOgL5qZWrHsJq1rWlrIzMV
xlIjCXu/UAKvdMJ6SUO8Z83otTUpkmiIvdsQWoxBZ7LQFRI7hqSsppgktSlBmoQf
C7lccp9JzkT09aVVIZYwSjxRr9d0b9sH4Bgv7xYiwGn709KcbC+5A95a+Ev5gDHI
M2z7vjBbXaNJ9ThMD8Kai8J0oB5xApsEdU0n9zHhmxqIh23ZnWh9GHiA8EfVLZZc
VoZP8+d/rNW1thj0XZmiFPT5ZI4Gx3VN2TG4s/pqg+7IhA7pPQeNp/2Ovdi5df69
qyLFyS5dvNZ3yPY4ZQphOvEH8AKMOFzippSMWrLGaawO9czDeuJnIp2NOYYhtyoD
p/TY4NaPxG+QlYGIbw26SKZ7Q3AcT2e1Go7fLzqnv0kp0Ee/2042tecoLrLWUmnq
Sh57bcnkRrGhl2Z5DoMNjKMhfvsS6BM7qICpocz1pNkVTb2GJT55K8cCTu0dAVJB
NdSS3p/GjViB/o2TAEI6nAclGVyfojy0T0T664LeDcaIDca5Q+qvwsSxqRgNBHJ6
SkOb/Cnzfvrfj5PjpiNxJxJJDd/yqvCAWnTkcHOFH3dkzDpYnf2f+L8RjWjYPYTI
6h69bFZwHFbNaklcUcJ1NFYN8rMOjoOfe58Ziawmo6HECxhE05q8rJM7LJIhL/en
vykwpatr+fcltS3BHnOvwq8wRV4aKXlDAlyipi48/H1/I6wRBF4KDsj7EPiS/IIM
hBGwdl3tveHGE5e/oEFLckK5AT1DJgRixPxSqT3vV+SaFUdKa+WLxhQFiAbhEXna
HwiabizvlSlv+cHu5JjhK9+KaCO1PkIWZDmhNft2bsThbV7DknCTvA2v3Y6I0IU9
AAteu2J6gxVfTDs+pazfRevI+YNoHa1Q+j+21483TxIxS8eccdrxgFkRa6YdNy+B
DA7h3in9wq53Lj+g8wkYcvbiU98+FytDgFK2mBGedeNXvjZtlvkTzvmHNwG+tOhK
SIXwaKzUO5n7KRPmiyiqf6CSX2O6t6/Uua5i6NvxTYv3yVQr7OHPB+fRolGzaVn9
tTChnADwY36OUA56bZ2AjLLbv5o+Dj566rkRX1lLLN5G0dmoHEEVPAmbNgwleVmg
HZvCk5TKsuwM03gqWWYC4xcIhSPXoYND9rEN23VxNNahjBbtWRvaH4mQ/zzrqhPa
BmJVV4+68sdqsltffUEcNe1lmyNkwUqPTuBqzgvN8Jw3UKg0BAoWX/cW3mhm/9+4
ZcniGhOKaI0I87vQYkHBfTalGeCSz1R4mEaxZLwM4Dii8jUjAapxYd81WJCeW2Vf
1og5RB7a4NS0y7WyUKFGU9INPQrOsrApHK9b0S8JqFQXMUBjgPaYfMYtHcIPKlia
WYlgyWUOp/PlkEYB1ZH+EeCNSZgiV/N91ga/I2HvH4NT457SWWmpc1bPG+ei0ytw
kjA0IyUyaW3ogI6oU7tngufXHC4fZmuWataZf9doxf9z+MLWg1DA72rMBxMyWQs0
ra+NoLpK2uhczWmaC4JMJC8/wKzhogLUziT60q/kJv131NNMgdM2Jb3AE27ojeOv
k0rtvvO2SZTqRAxFITjvAIfaYQ5PQpSlQwbmviH+/zBhk5Ux7ShTEee4it9rB72Y
7nyvtM6Ce4OpmvE4OYcsMvxaSOaOueSj1e1GxNGmPeLY74xW900wVykdS40+TUZm
jOCxR04HvYzoR56qbh6jP/TO3fEtMEbA/cQjOUqBNZEjeybLHRfAFZbqI7K7hy7Q
+F6T7sz/dDpXt+nA3xMn6vkHHg5HCDoOQQz7G8jGNmAXS+hZHrKdKRXfJZQugHJI
pBgRcEN3fHnKMru0nYKt/QcrLvUZgpEWsLpkjI6CWpkiU29x+zUCfHeTn5/L+KQ6
84Arf7q3Q30XyMXCWHrtU8TvwEo5xnmDq1O0tAcgfadoiG+4XHepZYiml48sXorU
+l32SkmUlucVhO/VUy04HR+tcJWTh/ikOxu1VzOP4x0Q89etu3gefsGncySGlnKn
4hlVPD0ESjbTM6MVI7ku8Xe3SAsWrky4SV61SkxlWPLsnoTyBLpECBOPg/i6p+lK
RgRaVrbtSV4EurwTZtoPJjixy/sMnKUDlb2p4lt9+kBf2osCR5gR6QfRo2HnBq84
KPSGcpLKdKPrvbhpUqxek70V4RsfEQDgWD/JKJaJWCYTvefZuXdID+WV+7Esw91/
wyLApgyHU4wA5qQ89qlt2sMmQwC0qiNTaZJ9w4mLTo8WLRY2ZmHTpz9Du8qNptKr
8avvF1/sjylEOybh8+W3dxKkFwyYin5aY4X99SimhqJ3anU8Wpou1zdSyUc1qMPQ
pA6I3G54q0H103GBCPtCg9QAAQKsAlcSyGf149b36+nO5D8+3e+oL+3qK29V+6R7
31VPg0H4CXpIbWHqPI3HmUM1WohdsDRE29cEc+JV9cy1k1BfTlIiqdoK9/kargCj
jO0QLK6RCSpHz6/lL2OMRFje3tT578aT5jaXM0+DChmwLw6ylkLX9z4tzEDSFLqW
u8AQXO1THrfHxAf1O/OUiAK2S8UAoh0m56MSxAwZHNPbpcZ8NHBCtq5+TzA43RSA
RKeAGMOjHOqGZQgZoxU9fx18KEiB3SUz7X03NzEsXic6R/CDkPJihmZmeNueZcvo
W9YOi75c5FfopPaJcYhdNSNsnm+Ts8WTAkx8EkEsy6LKwjOAbf9AymnKPH52qWS4
WxFdKquBhtx2hr3ewo7I7OktJIbDNE/dzhdtFjpnZpVu0mnE+rPsiWlTIYUyEonq
jTCXLbPyd2XiD9cMIxENZTrbJWqpCDWB7RK/TJKS67nwVns8L8LQLu+okZfP2G+k
H1TvWLAZhYgPJbR9C9KITzXmArUhHCnNVz5AJg7o5IpK7nb1fwrCnv09/JOclUV4
wEAvSN0dAdHYMm/dM8/M7X2kf9Zn1K+Ba3e/ONXovqoxE2cEkMqx8VR+WzPC2nTp
6K2NhYAa+w4Hth/2GlEtWFs6AQ4QkYtSqRI/MwYFYWbmpoLnuH30biGuTakEt9lS
5fmyMUqSDuigj3cIImwpUGjDXdvuKWqBohhhpvsvHTypMoc9SSkab987/pCiAzi1
6baJSMrEtmeE7KP2oeTs8lbMz4miQ2mCuUKIO6ISJQ5P8h5pthODS7gald+WrMvv
iv+fIJSU6WJlXv8nwwofZEL/shwwGIyOVTBZmFw1IUaGXHmrmO1pB2E24E80IzXt
6GFexQ1lXXs8em2BoOiTXOqGU5ER1CJHl7ounXrM/1jSN9x3ZdH1bQBYehFjv1AS
WeZZH1A7vokposXCdrtjIVW2gNKJFqzpQCUm1eltNzp4dOPQwcTEaSeUhgepZqMS
Gk228fn393oTUVH4jU6KmTwMgOALmClwOoq9N0fpWGp2605b5XJg3pk2mOceTqjh
Y8w5xpL/1+k8cZOR6R5/NHoxqLt6/6G6/9DAVakBhv13XhTAKOPTAC3wiw2r2BLB
nRSPmZPAz5DNMp8XbxnH8axdnbdwIbJ8eCwgv39ETMY2ShQBy7mf0U8DtVFxhf7g
tDeYyeWiRL9scy47bYpeR3WTishm+wfx8TfcQMpr8eHmRLy4NZZsw0cNUCrC6IyD
7zUmGiZULBjon8NZIGYjid4pMrx/L6IakHfYLvMDNLaVoG8jBR1Z9fCl4x2YNxca
y0TT+3PGe4dzyAdtHp7ghd7LODjMpXprIMZTD99CbyJUpz6oVW6nYga+RJ1umu3O
meeidWjxUXb1kE+ye2w31WRvatoKCxoVT0lYDSVChadmVHjGYMJzW9IkEK59g9Bw
HUuLTPUIemRwy+/5MImX89k50EChGiFyd8OL5PmcRnFMOijr4x/N94dV95c14T7r
hko1WgLA/zhsHC2hCZPfIjKiopBOdhd/ceOBh9UENi7VqiazAcq3AkEwZSTz4qV0
M3GvOjrYc1XnNfiybCT33PnT56IcJzefHZluUFp+AfwkfTbdo+wJ0v7hzP8kSJPh
igSF5nrb37k2fFUva5AOMhyvfkkWjJIcnuWT2rC4bxtltWPHEDzLFGdHpEqYhjjv
pD1rkfMEF/cAckbm4air7Sgx6xvwmwpxspClJXgbmJchddNqTBDVbrY/rKXEWvh/
tBFJI7EzO5DnfZpS4bYKfee5DIeU7KBAArJ9Y14zvEzmrZtwR2TTd7K33OnIGEBp
rTtEU4fKUyPc0SfUtRNW8Yi+HuXzf/beBB7c38AZL3XfHq2LBQsGfI4rD8nCEkSb
s2J5x1NK+yonAE5xG7Ov0EYJM0WEDWbjsG8+SJgvDGbQFwkmwb9DmyCKQ8lKu1gl
upvNqIO+c0gNdnIhP5nV2GPdIAzS41cS+m1TVLhPK1dxQH8rvwsbHhnQPz3kSFTH
iHrHWsWiSedJNxizkQG+Cm/AyMimwfdr7pv/wDInrpsg9vccqFUPUCQl1GOK5BAK
ZoBz+0I4+EFNYEPhG8VSsC1Z+7QVOsHy9vvZcC2fWaGHFb0ShuU7rkR4ZGM9FMkT
FVz3voSooYJhKL0dKn6IoKQHGFfMAKdSXdshOkAGjNgg6MEI6dKBQGBDeMQHXKKi
AQ6Ac/3Iw4J1/I6mXwaveVSGJ2YVQBlK2MLBUFTMwjChzGUlsKfPBmyZuEzanSmy
IxC5W2A2nUI8PpetDQV8BuOwzl0C039CBSaZgeXo1tZEuYfKwuHV3xGk69jINy5Z
3FRZPVox/dst7YpSbuoBWYXNup56ETsAM+q2CBJPNRLQRRMd4ZBAYg66Sxq6BiuF
d9MRdbWC2tfgSrRCCBnULhNGV9mc+TE6IOZiFyiH5AsBoxBvKwKDUh9W+LZVgBMs
/fZdfXAN1pmYeGsIeeNwRno7FVxR+TaSJ20pKexydqWRMrf9SLY1jAs/7bYF4UrB
49tp8XJVflOQNkQlWvs8x1xrHEhY5H2MNC4b3gV1zzDNcvx6GlpFF8f158h5jqhh
Uk/jr+U5FCJLlBnhRycSl7m2y5MGY3O1oiSI2wHQD7w5hN6pYVIvMPW53I7PaYnX
AfE+ykdxwlh7/aIl4pM9Twn8PLpmRGgdiJiG88omy3ee6N3G+5dinNyMEhemwq2r
8AcPnwaMPjRwpNAwrNEBStaM+T4oOsZYGqyHnoIxwFdLmHD6AFcYv+5QhF+x1yWs
XE8wxj4nyLembLaB2vJ+x3NF12NfQDIJQFh4yjMCCbwVoCbDDRnrAJq8/D18J3Hx
z4KJY91C5hZAQDbDuhm0eCFwvcyMCQPbtYEVweIYtMtuF8ELUxpxGpntKPWxbSbJ
D0vhOAwmgYv+ePF9Nczgbd9s92pdQMoFVuigbKfJ0GzM41pP3SAVZwB5oLiFu9n6
tJNIrRui/tO8Zkp01+yZg2Fk5NVOmtj9XhlyO82EXJ54bGEhVMAOtLqfm+eDc+xx
JrcANITdTNA4RD2Cm4Nnt9+ojBEL/BEGluNi2H3ZpeUdkhcfjnDcTYNHQ6ot3f2a
T9BOs9ajlBySiMoq0V/RGqogxrMZbmNnkgQh3IuWw/Ux9C4KsBmLFdTsy9zSqgNO
gvkLM2pJuGSWOpG0pgdr2gHOix8g3CHtJAOr9zevEFcwi4n70E8d6ZBUxRNORpcn
ctTP239livFokpFZaG4b7nhVx+Bj2xATmKGELYhSuxU0ZDPy1CfDtFLlnCuvkZCV
HM+OQSG2U60L8Rq/CfOH3cw3pJG8xe1TrKQodCNzaAmTx/noKfHKKAYg5Cick0aE
XV+MX2eH+ZHx03uS/SiBU29/ZHhrGMrsRIn1RI9RtgWUTE+dc33yR9iSfzMK5epP
oObFvMopFjdhNKv/ogwYE/G+JF+vZQTSgB5ggQxtgxA7h3omQqBQ6m1M9Mi0lr0G
fEXiGfAQEXrnop0InS9wz6y5lS/gPsxMMnjZNhoKGrl+cQwYub3/FhokZsjjopPI
hnY3DKXFM2Y06zibAl7bz7ibXyCB4xJz0NX9CMoH2j0dhx+owYejfbWOjFFQHeBY
ylSeJ5JqgMiG91l35ENppQgg+AY3E8bUiziVNDFPdNnB55C0OR+p+2ZKupXQNcGV
ZQRMee/2RnLUEaP43wwUbgSw4dtgUUzfIj//4sJgq8tVNsT3oUeQ+XLg87J6pvju
7NRSCDXGVMifN8fzevtOuvm/fUWBDYCGtjhR8a2R90eDZzgJYHGldDWksJtvzx9s
jnYvx4DMMeyE3s+Ixzfl1FzFoxQZue0HleCdCDWG1W5S9Fe722YuYWYloKcp+V5D
QSH7tDmQrmQH+bq3qfc3rCbGoLSnuPbsnD7CBEIKTleipQHNqLACEBTBL72bI++C
tAaXtHfdrPSyzh6fRhSDvwjPqJm7m333mSnAPsY0WbaNd4ocEl4ght4C/4QHln9z
+baZkIOtqBWIatyZM5XUHxmAIwUXQxqHqxJ1Vz7Mu4cFCpkZmcRZcuRkJAZR9RDV
1jt889/n+FeKyjOmP5kDqUe5bLlNdRb/JvUU4moU0TO5JMZ0gAv4eMY6jARemDAI
SFQRWvUVA0GZ+fp+E7iZOs/cyluu0530wgUeNHkVZ3TKHZibA2ndwIAi7DX5nZqe
96UbZHxmIe5RaTnApratjbfGHx5bNaezxPvBfNSZ4KWmJ6hIDtw9NhlvHtO4Onhn
yQknPnTycmGXA3xv693Mr1Ix8CKs0K8EIu+TP2RW0WbwtfBtYh4Z/2DuVlDmevPh
F4NfENzINiBWBczTT2E+x/Ajboib/AYhkPuKSshulux/BAigKRf7dWmnykAg40+R
JTJ2ghs3Ikrc233r3lkJn824oIAuksz2tUKzvQ8dGGcAWBpElwa39Zj4DdD63XwN
OKCsFWPr+f3fnc4OAtlfzAVETTYwYxsAJOjhfnf6gUVxIkZYjU6h24Jq9MSKtvGS
XqV6rGT0fKUx0/uw15xHPISF8H9VzsbxuoYCUUFxzpnXXUft+Z+1tsgViCMkDVp1
8bu6NOQmqf01k28jvNEzxgCha4C95Mstg0MPxlvw40U1QJ4/YfZ7gXMnLAN/BWT3
1OnBAS/4EXDIkGLPjWzALW1ERIpbjnIY+OvSKWpG2oblIX4ZRfLV95KBRTvIKEGh
W992P/9K0Q4EbQCSCZjEoX0zene5mkM9TEQOvRTW6EIRrqSphpGWhk4IeIXGKCQR
8jw8JmnNyWrGSrraOySCtsrdOlPQaz9s0ZqlC73hoVgwZNbekWzS1RfpaSaw49Ij
/kXDFS1YbDbTQsTUcNuzV2BhkX7UBL+ECxBklQJYIyQFN07VaQu44wsgniLKIoS/
LR1J86FWKp0yImErQySBgtOUGFpk7kN4jKJmaknlihm2hv0QK9dmeeoRsgguWGgi
QfSA6wS/cHTI7CpbYjEl5F680gy4bxIII4P6u6gN5Jl4jue4dftMzy1cDx+KD3ep
a0esomFmfjDKbnFbSNkAM7awRvA7ai/6Vcurq4hpVymgmSlW/37lC6W6MRois7tU
g5WAbXv/t3+OCKql0vv00/8yss4KNWqtAN3BfWmApINR9CSsNH3Ct+cxtJ3Ymc7/
t+cc062Q0Isr7uDBHlbM6s5ghj1zXjp6lpOtYRprGr2pxz/S3iyTf4YGyOAJinuf
goEpDNdCfV7kfmzINR4jesUjwGk2GCB3jG9+AtiOMxiWnJsIrNxjsjAxro48eOY0
w78tS/Oahx+OsNJMFF9R2+OUjym+ly7+6sdkarI/v6e5xorRoB6VwUwqcoqh9tCS
8rQMOZrGXGyygi8tmyk71tHpEmJvqUMYkRRYVaajKr3zv5U///yp58u+0GN32WnN
54YzAaFFuq5JD2jtZuhsh8kuLu73dxnVnEZtSDLqO+wISffw8NNsZG7pb9WN1Zcw
MsDIsoDNaORPOurEky/v+EkIPsyDtkI1S/Pv0D+/PsTLTRWh9JhxutVczMqSy/Hz
+jA4YRsODJ7mKL7pY7mdzKTfHECsFmuNimDkVwFmZau2I7q1ItiGmiKPgtTohdaF
vcmOZ3tGxz/4G+fhi5FE00qafTrWWtMilJziE7/E5u+6f0KMXfXC6us7poN9QaNh
Yu0izoAH6Klrcd8zSyYJVq5a3LW1P5htPSZLdWmfWcV/HKF9oEBMshqIZozw3zd9
zTX4yC9AZZIE/dpHeliMDjdNa4JEd3PFwHyGCLTzuzat7KSbry02o/ipBX1SSE+s
Y00O1fe4YLZCTerXEg1gMs8s96ACumThIbX+e/3F3hStg5Qwp3YVOEGjcFXhjx5g
o4UQQvG6ook3d5IDPBysjBLMD3AUIiS0z2WaldmaGF08BRy9xFnJ6Dc892ybpgmv
60vI2U5HLoDJkQHh+Y1qhFG4yMmjc9JaPASfwI2rVMRwdmn0QyobXaKZqbd+Jic3
bMw+so3k0gWwtZFOYpQ1OyKu9mZdvkuRkG+/QaY633rC7y8WBn99mpaV9n7uHw4b
5TC2i39Dn9G2Bbh7hzDSsUuNKEUfUf2EDzf0WioO0c5bRyOjsSxypHCs7zxloyFg
vG+/7SS38m0uqhOf6Dpx4yAEsfgId/sKOZa9IoXEdWGl88qiXjt+y+Lng4JyRROM
xAsWq5hf3fMdhx/EM0dJvf2r7jwymT3VMukV8VwmqyP3UL6r6SibHHozNTFBCsPo
RPE0VTtV33XhmGKeAkKqpu2Ryu1goCPISKzWXSd9WGZKgbrCP2YNU8JBa1Y2x8Ts
Ddvv2VmJYA/8r5jfGFJGj6VgWDGmaYKbi6HWODiNkpKZ2T0MX6lJRSBkoYkuDKU4
iMhFyppLOCbr4DKSb3lJU/dE6E7XUwKQmbm3wLlIhXSSpOmGnsOxv4llRk1khOyy
mPrbs4ape1B4I+Nmyy+tLZea6QTRxMU+gio0dWTkNLSSM+ANbbyHEI8Eox2MwOOT
YtB6Ac49/YfpyRkhyBAZbo1LnexZwclNd/gqR7U4BAUIz9L5c9odRdbKVx+HOz/J
QxGEf8Fyezyu5mnRUP6r1gbtl8XDrEey0YBuO1RvlXt8aP/nTppnHW2Yp5VqUTZV
wU5sxBjkVdEHIiMVYlcXH5G+A9ReRxAnjSfoKP77OCvlC9srAgFyMRz0No1ogjCj
6zupTf6PFBzLCsfVfWHOR1DqyXzURpBhUooo4JkdWzNIG/QSHCl8kgLnKVnQvuQ6
WbnGGOkSi5SL8gKoazQJkGUOIAWpzsnWOPtRFotysw/ym1ymhKAILxJY2tHd2wUX
tAw1yWTjI8E7OwxqGsDuwsRK40IntB7CMxdGvvGYoVGTtzWgK92FT4wIrflTj7ly
faVofYc8+F/r9/vkGaqMNjaGS2fiBligg+3DhzL4kGuXn7TulbwgkLHB+Z5r4Ql2
vyal8nbTtUiyzrAEitCntE8pjlYw1r2E+QULQkCyIbtPVWA3/SxNmMBFcPTlcwEG
KpfaJBLe1TkrATTU0r+wK7ixv2TJBjcbWk1RshGNtPGV0J1RyKGbWJ0KtdBjcx3S
GGaIsz3KUu800mSzRaogruMM2V4ggbPS63dYJ+thXhYtBO/6BxnCeoFI/8vJkz+U
rihSuLsQYEXc8I79Ycieeh4EPEd6DRXjgzmmiVUaASqgTo51wQEZGlDPgelrbtrl
r+csPFEd7NA1iaAv2qz9ANMfZFL5P30tGMXJQ5oxRneCEcBLTF2B4HJsrnuSXx+3
3Fwi6es9a7j8QxvTfO1fbhPJBxOoRHX/egCBDYLbGJbBABrRB92OXXXz6f87f55b
cG48ikDuLPQzrCowj6AJF9ni1IDYzRFpggda7lyu/cCLax2GRcL1Neg9vfU7p6dF
tHPQ5Wo27nOLklOn2975ZhNlOatbJ35nTBevyi2lnlrI2G0VDtSQByq+LeXCkz8p
+Lyksx9ubJRpWI3o/+S1Ej0nl3Nt4yX32lyGwNr4UZWYpMLnTYDMkqDlNmpeepLx
DiBPntIWnLgunv6Qtx4DpW0FiXx0oBn2NxwOXk9FSRJQ+vs2FjSRlGbo+7ghX+cd
Ahw2kz+B/ZVgZhRijxFmIuIbXKwNpHpU/u726ja+s+8h1CmG0M1md4UVRYWkaCbS
6Z2PQS85EIqeLrDDm8A5nK1E1CJJ12iTD3GzYqVsw25M/h4C30bnmhDbeUCS7egP
fj48whZ0CfCA7xW9VZDtlERsvbIXMddfkKveZeJeyVwtpr2/VQ1DRaayAEjlEJ+U
WnUbAHhocMtSBCF8mnTgwjGvBveAYvTP27PenN5xDdi7gDkY7Cd4L2vIxnZ+FtVZ
yHtrbNVowzIIGkNyV0XGL6MpewOjfnOiToOiz78IsN6rx+1CXkfp/tQ5AbmFY6Dc
A8ML0O0lr6B87qnS2dWLzvIBjP4pqWMJfpaQXyzDfPQ/zFzu34ep05t+0LAQMNcG
RzHZz4MWR2LjTx5yAyGHKWyCn2TWCemR6YJu9hca0NrlMYBsXx5VNJAFMCgRKhoS
UuIomTrnZyo0/a5n+zI7d7+4YbjrlmZN5imjtjyGpnGy9gf17JxZJl0is56Qmp51
A4flK9HsUs08DUKNpUOMFyxk+Lb0m2YqsJICs9pRaxmgIkbR1BlKnNc2S87e6G27
1okn8idflgCT0Auj4K1BB9oQoXC2KUk2HMZ9wsUHXIZ4a4hnUd3evgISPnQfRWkL
5KX5KnXzUpauZF9fDPKh179/47CRF5r9MvgvgSOAEqv+LrRYQZSymD+a+p4r+zKI
xJUyfFEDNMhEAGAklDrwnaw5PXB0FMMaLH1UUtrYZYvgAS7P79/wgX0OYlgyxt3f
d5YYOxfMBeLlkYujsTUuG4TJ/PWWL+LCnElz7tWslQ2J2ISxFtwv+CrmGCOg2afJ
4A4/sjzlckXOUnYWHYIrYBq0jSbT+n7uTc2a0mjGNNjn8DChHKZ7vQpnxEOj8N5j
V8ICfgGyvjc2DPt4/uMM48I/E+sI70r+RlmzP2k0/elwR6uLQ9Lm34Qiu+5OBZTV
NLCAcuLzhYFzUC/w2PudSJNBADumKLwtPUX5j5Qcch7Cdr9HN12wFD7cOFWAOMxP
d6s0ornWW4DkNAJxJSqFyu8bfCn2FrnGmIGnzXv3BMb/rK5FBsERlpzrKCo+kpPr
1ATTPSvqxBh/MS6T9o3vBTOmlv2cZ2wUKnlDwIIEAuXNwxfqNHWpLIMn4fJFXpZq
2lAhXPkNnbPi7yODkaOb4u60up+8YdUazuLigGSkG1+ky16qAhag68etQq7138Bu
+r3d2iXKc/M0g55UOxzDRzs/MnATPW+kDxC+LBC0Y4uiViWy8yDPqtqNv0j/b9Gv
x8DJQ2uCrEzUSLRLbx8WEEJ5EpXJBkcl+TQNa0ODW2ySkU52Sw0L77F6RRgK9Z9R
eSTgMmOU25WqlaeTdFztyjY+usvFbt+0aC+E7c9gi6k81bnIQOQtFFkQY1Dj/is9
1rt8HEFtfEMkwzNcxabrFPUxNJK+eRMYctRwTRquVLkVzQKRQsB+aVN7uAEzwphZ
EP8Ofh0iVgLgNymUn6i9On8laJFf1e3xx1seSqqWzfFzREscfC4l7lfCCaz5gqr0
aUvpu7GUWFzDzZtohrMUkv6BqY3qDkNM0MntpytKWkv2ozXhFvGTc6zR0+gUjRKC
N1t5piwNvGUDuwZioi/xIUBm5N1AzCPv/EpqNgLl5/tFPGD28ohzJLrf8B15hOpC
yVd0apSv0vJmMLvPV3j2OZO9XPDdA/fnmF2RPnwABVBin3o+TJwoN3WZjCkFa11n
Kr/s2ueIcAZx/c8LkXvsW7+QnqSFON7saJOhjWpTcmgz39ZUj1LNtLjfQNHpwf+S
QrbuwotPcBrs1dgZ2inVW8XH+kafgqt62u8k9Zcwlt5ZBK9gZNP/dadQWoKfnnmH
+KEeaKpP8SOf2SAVgyj+qElFvfDDUeWa9b6KSd/7aBnaAe4h12ulaP5Zl9p5Kzfb
O/mrbJ8TcRQxUeqUnWJNc9j0pMKDerJhiJEmANCTWmj+PLYCIQ4B0/LDEHkeKTgD
15DZ/yFidlqbFzrwZUn4aDZn0PzcZwGYRmitKAdNU8DDIbgvGOoUMBEWmlJCfykA
QFJq0+HayiZNUmuKi0YmhbYwjiWG1qVm+vh//bLILQHBFh9+EIXvQHHc34Tky6AY
wWM4L7En4dpU7QxZv3NYgKevWeXnKIdY53uJ/L1/4/KOoNRIpU2NphwtI0lqjkDO
hsfWYz+7oAAIdttC2ew+BoFzz7RGFd6l0mTGTDWgcNLao59ZgkdE9ELaWPTX1iRT
FlJ9X6gNZuQMOymq68jdmoO0B6bFgdBpU7c3qj5e9Z7gNLjkY0G+4PWB27SEU3yq
IWdueoNNGQuoveArmgEIq86DHJj4Ia40yPej/R79ztoPoi29lYpp0/5EnNNV1Ita
TgRy0b2mry/l8HymKqNEdVpOswo0xPf4pehtFyqbhIIcOgTvTeFRVBAxhHAjOOp3
34x7UujCO66Im3Mrqu5875+N5vFz+v+GejrPVm3lBd2ogFejmiAuIKd4csGolPHA
GQCwAU8VNuqmAx02JBfaLrHSJDNllMdEVx+HamCuFRefiFUU6SWdo6LnBUu9TeV6
2ifkZuOBejRwCx0EN8WeLto0sADrxSqoa8n6ylh0APg05GA/uRIz4U7XcTl80z7n
LjuO8GyjSeomnVMVWp4BDr/bZGw9h7Wy9juPThqxKcbeYQ5WLKmQJW45E+c8QLIz
nYuQFNCkcTW4oRAEn+MWZxr8rT11r5ge3s2JwkxUMty9VcRaOECADSwvVREl3zp1
33Ab4iRjcsmzYkqCfO+50ZxEGS40hbY8qOGcVMIt0+aPNE43NYdVqNJRTg9th/kX
jvhMRPB6nwro/gr8bnTtufawidkFtM8KxL8rI3Vx8yEsyL/3VELYer1Zn1H8rRV3
2umkJCxrdwduWRs2Z/tEST6F4tPSK6qCgY3XGVocnMoaLFH6t5RKDHKr+Z6x7bee
N9xul2Yr1asVLn1dZZLMquL+6EX0AqKXJZmzagSKwH+YrhqVRYpZRmHa1LsgDWBa
E6iL+E/Hyo6vTLEnnL75YWwHSkzSPlvBYeGOh9M4CwXlVxHX80prsk+geaA/kgya
GK0skgT4eeVQQSliCf4frogPrqRETCiF/3C3kHnZqX4j9kLWeVuIPB7QncfqmabA
yTPOTKb+Tn7cS1etaTPhQs6k3pQuPEFfKmCrS708heWX8jqfiR5FAuy2gl6LaazJ
fA5iksOZQmD/UmP9fZcUwhgncE3EUkUS4/EadwBEub9M+rWPHbx9WLdOWSQHGDFp
IrhMiNH600p8Ftwb+StF8Pnlk/Mp+xywXZU2jibfooEXoTY245Dkn8ODxyoJuv07
QwZHuUCpt5LcXw3M+hNRWd0EATJB564u7Wf/22r8LZWswVLeNS2LDqlAhlqldmcP
svHr4h6V7yhf/OlWdeosSKGnFQ/XrfLX0ptrbGU9aauH2bSnwP+t0qQwMHgpJIme
JkFp49xQYyYYd2FsvFfKGcko3+CUifeZJHlG0I+48LZXPadEe0B6JPDYubc2c+43
/+Z2XO/Wd+GXqj+AC4nxzjwbUWUQbzb7WA8YwRJY5IYpDb8aTnpaSCA6qn04gLtT
ECKdfiOe2l5aWsZQjbYVjacdaHWhYEQLlZKTDWzErZNmwPgybMzAX14Tnl++tO2k
Ja3DqYMEhaJc3lmWb1IHm+AkyKGnvaBWEqbXrj5WdpHxhW2I3oR16skYNlwmpv/F
vWoQTMCGFE3bXs24ruWBpPxnDIWM30W28twlLy+978JhubuNC6yNvp+ZrI03Ev0l
GHr3HTATHHVH87gcE2g415rHoaRmpu6BBiXVzaHCbS/Xz7YCxxXhJw6SqTOsnwc5
qtQocBdtqpP9UvYRmCvgnwCNyG8Mgkf4KYomMP4YdsMMc0652Y9Upi1ympS7e9bG
3MfhBtOd+vQoODntFuV9npAkSwt6noJCAItlnzgKcIvWY/7D8vW91e6pHt4WdfRv
UfHtSE4SrJHqOJmWghLsbLcwyaGnkF+jPPNr8yt8qQfnufiCakFVdxQRki1PMNbA
d2s0vfj0PztvUbavKVDSQggxY7SAS3wD2y8fm51iK0Tr9LpdDc4y5rV5K7hRuQAW
3qYkJEtz+5buVYvVb/USmhTOKlvhmtcLYXW0cdRaMUNscYsruZyIhvrQ5zOqsMIl
+qLTy3fWdeHu9/MkTAQ+iDFs15NK6iFrixvP2sepbxT4z6X+6iT6e56Q+L1dZSUD
YGPqyPnyx/3xArBQA5kp7w3bj2T2G+GGu/orKwKht6+oBsO44AE0DiYbWDBO8L2W
S2PLhTAXVuVdWBHkLZ6ibuavbSFJN5Y8sy6MCBJfbMsv/S9J5BUCz3uG+ewq8LKf
Wff8rtx0jGloG5/wnHa2+p9xjAI0HKG7Kl+9SvNJ9/eKjTToOJCAWER3ABKXvNuB
6qtSpM69Td/PKSyy+w27iePBG/e0dta8x0OTgAWgu8bWYvkKJ71BLOoAVCUNWGEk
m24k77LzufNgpFxUAlHk6HeSGgQOIB/CvkoZeK/OxYfOtWtJ8p5YXH47cu3p8Zdz
hwYEsOLTKDUu1ilcz2wstXJovG7LfG7YBOmcN9k3e+esd+BKzGEwWC5Y+TJEBYyy
Dwd9wxchjSMHBGWM+AepnDrdd+OoK1WeFYShjw4KegPC8t0uF01a3tsCwT7qZvHB
k4AoCsNUXpp6BvlSVXSQMQPHF4rCzcBtRhR0QooPrHc2/dQU68CgSczHZfvtl1rx
TxG8PSrpVGjPAf9fkXN7o5cB12n5B9xA7tYfpIIvIegzMIPOPBj2tZuiJ3+mk8B7
gCZySd3IqW6KxJ+3YiVpGgPq40NdRWPWR0nH2moFLpr4q8V/nbFG/1RAdC9b7YC6
d3ApnshkoC0whW3BDg72TEbeiCZHdDtJ/JPoudy7lEU21nsTbd5aoTrUTPLQSEXz
K3VUyAN9MZYn7ZyoOdi06tTuh4Es8oszBZvTCD0gAiN3fi6lMeKlsiPOhsP36bFz
Ii6PaJZUShqXMHPczA3LWNs5WKnRs871ycX/Uafh6VS/0AKhIJf9tjybacGz7mXl
1MCVhiaQ7LMGzMMp/Ft2j3HlllkSR6HjuIEffm/VSc3HYVRz+xTnGrn0wKamAJAB
jx4m6YJ8XEGahe69iTCxJo6JafJXDBRATuHvKT7ZvQ9gHivwyFatM61+RSoV3Dq1
jyMY0WTTKR0ljiKBvud+BJ+jGMZNDxCDpCZQj/Hyod6kfMiEueivaOtAoEp4UzOz
u75UpAZbJLaFfxmRSGfhC38GMszfNatm6CJO+ClWhkGYcMG+gVZkhtrhZOvubnek
ibD5U7VzT0dqHxajWPGjTiYGqDcsbnfZsbXWRhwN4zRuQblOc20aWBFScW3GOjp8
K418sidodnn/LqZ4CvFLrsaxn6rYOdRKAZFK2noS+ompWtanKKBBAzbJ+S/v3O3n
eaGDLskzbA5l4HvZ24qvpaGYLHUEOWH2qaDXGfHy5zSQX3Ka4K2oKZIAztxbU9OB
ZDDdb+4dDlcdCvA6Ln0bPdzNVGCy3UAExDB778XpmOp6OXWJ+ee6py4o4T8uAoRd
jLzwmM9QNjlL/CHn+tgYUtbrVTJ8nkbYTxNwmnsyAB0gnsgE4ijEwBPrbhRiwMvE
TmfZy/mZ68rsEnNw5dKHFMkUYWpy758WbwNKKRHAs/06dcxNCmXmJsAeMdZWtALz
GwIOO+wYONMHXZ6uoMhwUqAXRY5wieZtE9VUCzMyumO5+cnHftQ05G9/GJSbeOwu
tvbbWGboRVCEnjSx2gC7JQcixOPVi6YPfjZEXATdV9cJiU3PV050wPzRjsFLcUNK
Yijt0hROMd0V3mRTFkE8fXSt744IpM+IZq5N8S10dlVoqbOR+t/tSQBimIfesL2U
GSQnhf7rF7eJ0Z3qmJKSURe28woNdPa0+7XA7frcqTJ1Y8vOBImOkmAHEbCcLD74
VX/g/MlvlCwNhLAB2EjwhkmYwMRQMzkrdEDUQCzfFYto0W34MlGMvJv5l2E0Nnfl
DCIyfaJV2qFKmYgML3OJGcMM5T9wpWnYVr8MrhfmE+BVYuNgluzsSm0Nq4P+vlPX
WnRGo3KgAoKUFamnK+LiEOb6bSUr5JrqOi30DwuOiNdbCcx02qU/yjCvDq1Gnww/
e9jOg9bpIemCMyt8XQasQBlVGLpVoVwFOrpDVxGofYYAg/V5roGwCUl2081fhdWM
xbym15KuKMkW7nBWN/aeyctOGV37XL8IaG7fq05ei5n3vE6vtb1eatznNh/yACEZ
OtiFMgNSyOCNHw51rJY6g6dMZ1kIO5FuLT0JmN/qRsDsKj8AlEyO+0yShc9K1jxp
4HTWOvjH0MxokFnN5lGb2ez5U6GBiamtEATkVvZN1ukg2nNA91ZT3tU7I+qq8gMI
FZr4apinkqFuvNzGP4ZcLmU+2ZRuQUJOOo3k3l9Tta6REjOncYl/+qZAdlJx07fm
K1cxsFHCbnqlyUE3yLRjow/O3k/qJTQ9RU0ZVhFCkPDXjT+UDep23oJ47eFFgfNW
iPxE5MgAPbSZkLkmlxnX/NfU3IgtyXw/A9ogi0uBQuM0TrqQ1Onxv8HE3THXOZfb
teH7e0ICgfTlZHn8JiuyBIN9U+4SWudvm51925BOuoU8I+NUaWaHkqZwNc2PYJDj
JjKdtq3IfZpPwFZCd0/nZ3O0qWT+cAYLOzJqqXQWrlBP3hGmbOz8/7t/RTfUUPaI
C05+54ZpYfgIl5XtK8Gh0FPBU6vo76/wK4p5WiRqDCt5exNt+0o2WL+fnOSqGiEA
qreCYk30YGTUzSJbnIstR0OZoXQsq6EXqZJd7EnSeXUZrLCZ66JT2YjroG+BQjYa
dqSqBNUPfWcnmf+yzYuRSdKbB0FFYHjgNM2RMwN+kPYXaIEYmRhIOpL+zSNIcB3x
VDaTX/XhhExhpiWrSBkmwBZujTie7H0cVhudGIDvqbFqE6NO6nDV1EPNyWjapwa8
2pXC1vOb8B5vqEQMfVHs286DSCx+eXRtic0vWfwY41SqKSB8iKJibCvnENu9v5ge
WIS6Nu9MCCUuLqPI38FX0eh2CwnCe8nlbILnLJDa5lymTZ5cpRJDgI6VZOUVQqAa
cuUtuePV6NBzyVSNBJlxjp41FBLpF01kdRGDIyNLp4AGJ6pCK6EHNyP45b7+ZuJX
cUI5+5J9bKdRYpy0WTz4FbyvXCbxydGp87GN0IYcavfbqQZlygy6Q4iamV8alVKc
iz/EXCmWSa5kBfxsEqun8J+4rKUK4fZ65Kx2bXxIdOw/BO1bwKx1CUoJV57mv6N5
xznJ1TB3TUzpQYwT9pmW23EYhZreCQ4CbRq2jt6bIHBPPjwHiRWgjzgbzq2q4Zxm
MiCxtLKJzazSa+hv4GnZ62+9gU5M9bzQ9DPWsduMI/y/p8UPq0lR4mgJp+9Ofja8
A3vKH2Wgsd+eWdKc5BopTqyOuL94GDRWPKF2eVe81qe7rQpogAotSBQuT1Jx3nkF
MecjNJSechuLjcCwLkMJWiuhNWx8QEK2wt+UqFBQQlVv9cJD40aP+aQFV2HEMlDc
VbU3yrIsXsr4YbJfAxrVYjwZ+UEtCCgMYnoAlOY+C9Tbb3WzOk+hbgSJxr9Bjzko
HziJb1bC57/vMB2UOijSgmlQe1evhKZD+YwdDxoMTpwi34VtCWeK3rzu9AOs6vkE
b3pBF9py4d7vEXkiCzdATl+kaXypszkUEyWwFZykbZ7q8igjXVT55FUgYjMS7mdC
MwGwLqHOMh6zJfWoIJ+Wx+5XJJ9jxC7xlokZvfnyxhZWwAztWikfbYSImYGnZUuP
Zs3WzOcrwSHDa6ypMKhlEEwABeR9+A+UwetAwhGkOpisWOp0PnmBAjFnDDR/Zwc2
ZzcpHDmGmGNFyHefWWvdMorO8l1XGAkT2sYezg0k91cK8zLt2Hw0alaFcl4yHGIr
DWALUXv6G1VEYv/Re72iFQJLAs09GpyLH+43vB6ACvWopXsqSslBhEFeNb2cTKCQ
zglCzPOiE5iufC5xAHjW9jBVrBUAcRD54WTCkPg8Fw8GlppQdBaCZqQzbGXyty+L
cYM527pRoQ4cvJI/CyS0CiOL76we0fXAuhOgosc3qYBq9jzed1yiA6LDWJ0PAcf4
6xEN+3ah9Dbow2lrzfHwuKYN0cUo5MwFP27zD1hpLjNQY4cmOav8dso8sv6tEhYF
wxcUAWvCXlDIV3tQOEXUHDA7PLTLfHs8dJnTuY3CJAanZlFs3cNZGuCMIKoFAMie
vHdiBC3+5vBT+UWSpWzPSbZ++VVU8I6F51tjAshEUFpSPeZlsNwLncc5oIv6hrpt
RmT9F6ilVMQoCH+R4RdDf4UvcZAQ6w0XLejM7FhGyQ1ziPGsAe0MRNtseU2vf5dr
lyIpwKsBJRVLgKiHMkX+pAVVyMluTDxnbjqRY7fDtufnyHFNB8IReSBh2v6a7tVi
dDxH5TJWA8vblYh6LpR5ETz5zoVgBcspiqPf8kgyHb9MpP+rDnIylnvhMCDkAB1H
/g5xyCoZn/Mj9RPKBy6o9VWgHMOblsB3+M4ixX9XfMdPOI+SZfZ5skaSkcczJEoa
ADTNw9uc5U9q2ZIlxTC5akoN5Plj/K7Ec8zjRqXtx1881VeZ+iway43si/HnPhCF
OkqDd1tAkW78+1JsEir2YXB/H5rFH0mTUuln8Ij/NSbU9VUglszhGT4c0igxuJ4+
EvPSui/PBh7o2qd7H5B14h1vwakR6yOnnMtbIRKkGUtNSOzU9iH8Ub+ZfE1R/34p
6vBpo8U0WpXEIq7JIjdD7pj2+9HvqkJsfoB5t0Dg/WO0yuUdFO4VAP0l9zicbszP
3TSKQpioEKAU7uznbWTLf03a1vPRI2xqTwCKtRZeidRFMLgo6GzRH28/bDkxzfWO
1sOxPrDhX2aAUL7L2J16YBW4Drt8HPBOBj24SJC+tKm/L3GKgisA7hAp50xqxHkb
CexU9vB166roCPv7J0ml8U9BiJSlZtAOFQuNM/nGct9FClCL0BP74/8zaga9uaFZ
w22khRwlZAcJencMIpPzwUxN1lOpf8ocon9LaJkJPVM3QUcPIHgsj+xZavq9U1G1
lDAy7m2rbSGUV/1hzcSiig5jfCHyn8jq9EaFrG37xnX64GTAlwJCzTTsR+uh1o7k
RwDZNbekv5xlHLE9JTWHv1ZKqj87lIHR27yN6RcHKMSZH/A6n1SNaLohhMyYPcyA
9/ydh3vfVoUU1bs388vjvoLm9IdttLQDXoufvJ9uoTW9BIfEdTqguXxPt2UxK6PG
xWTRj2Sz1wem+LGNBbPw+f82ji31SsCK9POmEWyvCOGZfc4vp2j9CEqaoxb8UK2x
GYAd2YFCC0ApjOBFYtIWUgec8RueSAu1+ERPWbZkHuNZmQ/BRK5c9W1WXdgY0Bps
vkSsFhRRZSaEORdAGER+piz6OJ1APi8vKMY0OJ97sK7/tnc7b5oXQXZ+fU2tw1X9
7jGqo3nBrOm7ycW/C9Ni6fIx+8EP8ltaktr9POMBphEv+x17H6WLeD8xpEYZ59pR
5uWKn3WijV3rzDdiJdhAeJz8y3qf6x9eEKpW45CDLOX9jtA5d/Mx2qJzCl8+l4RX
YKLiXJa37r6EolhtGv9NZeScKMqbtvvrAxDCew2IkYIg47zSpBuND14y49VkJ/XJ
J39kd5L9ne2HeXqkPnaeBqJIbOoboCcoHEvSgiQSdceZ1IZCg9Z39COKjDPcDslg
pwdqrHRRlQ8qOD+xg3ngh5DiEkC6MDsBwdKDJFM/zd1hORt/C6N24djNwQURK6Rc
kueu8/bXAyBbkN40VOXMwiyvSXoVVnrh8ZvZLG+9teRbqWhle5sC746ozIMrEP+6
wLXt9NKQ/pXsxC4p1+PqgEjL6vceE0rCcb1W3k4+yvD86B6ejggTXRSvOzeFSPZb
KcXZs9fU/NydT4PfrATz/PprhW8p6GSe0AoammsD8bDrCmeARzp3g92iqQGz/TM2
G79vwGezSmnPcgMTvkhhOtGMErfhI2GqW0euQGO5LiF9BRffHxADZwiG+2FbiT3Z
trbD70xZMYp+5OhMtRvIj0wlFRrPatnM14YgFQoWDKkQzP5cBW0w7iBCUEualMmG
0PDOk4tRczDaO/jcHteaorOcUCtC9Sr9Y4NTev3yfnXXqRhf2iB1fQRT6AoKFxp1
Cjwkxt4r+i2Iz4NjAkk1rvmx8EWiJNwrsoXKryLp2jMWKe+vGJduKy+7sm6XUTEV
kgmLzqEmtKazBGSgfLbvJoTSuFOXMxNR2bPI1MbQlPns21z/HJrpHzCB0Akk5V56
ZLRfl4QNd4zZILzTZeZv23BDDsatzDAHnW7Hg81JZS2Uhb7mQru9TtE4Qa6f+pRm
5TYxhRFsj22u4pX3hNw7aRTvF8XY45LVK5wgeZY1vsSWKxEX0gTrDq5LqRnjIgJG
QAT6QqZkio2JGmBNTQlMV2sXVTXQc6Hep1nZ3P/TGwE7pVUcBAXx4M3KAiTrE0ta
4y3mp1AZYie3bwY6RuFArym4SxvfU6TyPyN79eRaqhCP39VjXp5dVzFGTnXpwI0m
iEhPsxdK9o+SjuKI4MzUqHtyrGRS8RLINTfLBv5mXZMUsJmWWoteSG2p9HdhVFU2
9tKRJmdoqVdLZaWWgTgDTlnU6kUd9d6VEbPRxC6K0NRr+NPFtC5IXOMM+JsgzVBA
+ejIbO7CnZlUKPxPCU340QkwcWCqpT9cRNltXvhdcrmaSdR/uVv0Avx9/kMOwohn
DU1pPd+V6CEicXuyw5xJfdFcyOf8hAcDvCosmLxhpHogAu9UqPqidZ48fSfqMAho
CFFqZw4zUzZHBdeFgfzttle/PgPmIeZvpLUKazbjvYnlFOAQi6NYiIysGk7f4OqS
iekj2NDYDfpuJuoVnJ0WT/skAU1FGlSHlH+P0xq6XWTmThPL0tPJQGOtxauw6MVd
FWax8O57Qt5IMBJOZ8w53RmdAUE4dN1gI1MqKz2gzc/YoGPxF+WD90ghySXhp7tF
g2c9MjdtmpBFcjpjZEzL3o05BUs9kCbqpYDLvNxjR22y1uI74PwIF01HH2itVA6+
IgjrjTl/nPnE0U3cpV5/Ihsam9fU7KB4q40gmYmqA9Y/4N6bfAQ9AMsJKCB+FKaN
biPrHDe72Orx0Bwst/fgACOatoUxaiCXv0JmguC+LlDOAk9/D0c3xIRkXSO1Z5XC
9Z4Z+QWolr3V9PELVD/4tcXGdmSqcQjBqZ+DPUItkyghAYkKt4+ehZCx1mt0sXkr
7YuSQYQQdn6hLx3zAYoq+U9OkPJBU769jLvhJmleEOwWFxBejDYKh9mojTtxmB0z
wGXF7YNALn/B7rxX4qVqAR+QIUAlT4rCm6Z6bP851XV22gwV+E5sc9gES5O5FDrk
0ZN4/kEpunKgdiUfO6TsUTpFNVZBoi0TQYCP3D2Rc0xKOzjUMFSF64lEsj3UvfyP
deq2TdDgRU3kCl1YSi6Fhiks+fBhjB6vYWYpfb+Y+TD40xmOoElM5ARnwm4NoNNe
QnzVaP2ebzuGJDiHcVOoims/qmmposyE7mQwv2v55MJ3jQIozeRhDx37hQ7i5TXw
Qy+hkAf57oFxKYqNyaxMWefH2LP5m1UxE9iLLvnt23myHmM3/egV7qvyFcES+CSi
2SQ7SjAWxPXZeomAFFnoB1NaaHkgnPWVGdx8RX5mtKzGWO6SwTPfALFQMnCvE6K5
0SQXhnLnqMItWzzPMK8aGysIdx28MHUgJ+PkE1m+ved6sC5y7mgMb6D7x3588/hT
T6QSYW2w+d59Esswdrl2ia1oszQE7+B0EAOzLrQ9/QGt91LQHyom8XwHtQ7A9Na/
cQ/lth2roNIRQFWzH1C2I0M9m5hNcuMMwylJivVtg/ZV+HNAFSQC1o8D+7NeRE2A
c75EEOa0F2PL2IpC6Y0MI4UrXq/Hnsw1lVo+LnpgaalI5ylqFtiHN0ccHsb95cju
tLdQmyDYEFz4gHdzc1TSDdKSz7kS9sPa7J8eYvqVg4sWd3ZAB++AOAAQZqpwkvpT
ONSg5tZZP56mVW3A9KWb0GAzaYDTc3DgIsIu+xQICmSUIFa3scCxqJdQ+RVfQmaD
Gut3/tm2yEna/ixUZ8XtF8ElP8lunWvDbYe2eSGKDy8/zMc/+ix2xp5G2cGpPukw
7DAYyYTlXSyQsq9GgISoQOFij1B0BkuCqDRh2Lr6lc462KFzR9j/AUbWy0sKw3MT
yEMeLFriXR01hsaEK9e6AJhm8Igu688DxgV34TsZxJEz5FMb+nrdIoW0EyR4Rlje
l+AfVmtcNR+p1IkyxjvcOfL5DBLzTKO7hu1joELe5IQ96YK3d3ok46d2+6d9+ahg
nXvHld2XlwJ0CN4G7nKyCeV3XfCG1M3sdhiHQYH4MzpDL6fYBgteNXhTbekU8sF3
scC7K4gAjC7/HQ+sa9NTEAr1wZEkYblQ7JnFFholWaJudSIKk92AVXp4qNT12mwp
fV/+CDB8DFpYfbmD4f4KNrA9UflQZPRus+Sfqd6ztmOlHbBB/W0eGW0wQ+BXshA3
W1ycpniN1lS3mKB2ENawWc/wybLL0BufyeaoXsWO87F7kOBovLxPSVb4AvnhhUl6
tUgAa59bHJxt7a2da2Q6cJw+WAhWQoLCwntvSCQOX8omeBY37QL2UWlNAUizlyQ+
uU1vNvFByEbuqRwsXa/roarm/23cSgKXW9eUpgSlRaOByt+zGKRXY5+Q4JouKQhS
SdlPECHs5GhLbN8v61wWM5OOxEt6gqLlT9a1PQEIvrqWuHOFC1Z0lvQh/CqhBFcI
irREK1j7zbeUJjPYQUJHHl9HsZot89lV4MUbqEN7q2D2UWY8Uup5Qmd8aVmaRErR
ZOHAdE3J/SUsdhAc7+GA6EjBrneWtcVBATUIrSzRUklw17CZYr0CReWqNyjaXD6a
QgeManwgu1gtE3CanSL2g0Wj0SzIiEMGZ1u9Qwalug0SwD7inZkl4Sx68XhxjX2q
+sSjt6dyMZgaADnmgYlM9LBcgciRZVMUvWMZ5SNO7qh+oLVYgsMP/08Y7nXb+am5
SnsF09/EpSQF2LrpwafZEF5fyc3yjNVa1yl9rK4WlSI6B0H79Qcm9jGQcVueQh+i
VwADmdEPQMkKwPg0gwmQOblMBUaswmqwOc+QvE6TpRHS9D035Lr2lOdGHTRyVv6+
EpVJPsTxysGeM7DzM8/RoUP23AQtJ79qhU7BncxDJCFRmcJm+F+a8pAglP/JpnYm
bJj/CVRx8f781IRLNoeCsV5lggcaPTC7c1U/cA1iHm8aaXn0KooKHw805mj2AwF5
Wte/DGLtVQDpERsQ5GSPoOHgw5ZrDCTNBh9QJUjt9oBEPDguvO1rPke3EpxzW1bY
jPcyCjn1LkyaNvskXd/oKu5CYveiiPQQ/odzTvtBSVGq6o493IEo4RWBe+M69WSl
6g0JSatTfzi7J+85kBuHToVT1txwXkFbCN+947m5Ag2IHDbmGdZGJ7nDfSN3cheC
/TcXZmiLqw4c3t6jaMlx0hM7B7rM6vCqh/FJ1NAuaQMvfT/gq+nF6fZi8EDUgLNN
A7ZfW5p7/cCtjVI8sxbMJ3DesgsTO241qCipnl7ARiJXcyCqc1rrigjNyywH7KBI
wrqAsnsxsapx/j1ufppzgsKpAgNTegeOHZNKS0TExc79tSu8jq7I9kgGGS4HMb4S
sTI2xLqAiqCGoZevbYjml7pA2rVsv2pRTtzvEpkGToEDDjM/YlQN69WzAhk6+uOn
EaKJ8XLDf+kXqi/YCwZEUqVH3eGwX/cexFCDGnQ5iXrGvePUFPAhiEMYCMDS/enV
UT8Kot0LmB9Wfc/UsHq6nYvVARu1x1TnZy9ZzyjDK23mG9FylAmApzTku5aIONva
is4nN2DYhJ5UINAVA4v++mW6wqI9iNVgbBqewFtWGR3wObYAb/Mh6gPEIUmIXyPC
rXXutbTnM1+1EHUcSGNbD39mFLsHYBjPm7Ktyk6AHwQrzMcgalnKaA5Ya32n73EW
7vlm+V0yw+yaT512vIfZB65TTuYuMn89q/21AlNvqiA6xrq6uTW69kfBF8BlsRhy
l/zcXCKbCyPv8/6cKG+H+c3VI8AI7ChyFbs2by77HzfRffAORCXO1i+FUeH+Svmy
k7+TaORO9lLEurD7T53KO8Kc047TalTgB8kVe2NgM5kf99bKD4++tt00q/7VTwMv
PQQxwrfZ+//Qoz08qQMFJyx0A/C4WYeYfPr8ep7rfI8VOPJwc58bTH/2VOq1r6z5
aZP+s7z+RA6nWuMvpvY3PcWgGBLqZwaI2x8i7GI2YSujgMjXMdvTD9TKPqpBF53v
QLHLH1AVWetRSofPXAqgsJwBuWPEAMZ+oIqSh4oufb8lqYXsCajjNgMXGc+YGMfK
ELJORN5sL/kSTU1IEc6og4t1fj1KwQKzQB71sLaSqtdxXrLoiVaT4Jw1zWPTR2Pw
a69pW9bqvIgbEf6C9oWBr3C8nymb5isbAm6BiN8HXUR6MGUdL/fJvrfCWfbH/EoL
bB/K1e8C+IuzXh3Bh9OV8G95LKqOamBDTjg6H5Yzci1NUPhuB5NtTSZSSHHDbBjH
+lp7WTwSOgJqnnkAkmuTZLl14G3YSJ+yfDJN7GWMbN/461Rb4pDgQKHCFTSU+C5n
KGDDN3/nF162GYwUxuWC1E1/XdJ1GTUTsDs748KGbUnBESDfetPNgUWnIXclr6MN
2gBvUBzswAIrjrubjEoSxGzijuwBOMBn4H+VGHQHNBpV3x8mAi1CE9m4r9ZcGn5p
FEUktSdXVdGCqZIW3bOM+dA3WxwyqUFvfgyCj5rpsWJePrL3ilVLjw0X/1kFAsPm
szc6dt+2gFaiB81MqN+qM5KLeDOeKXeVcUwuz1iCC86S2UIDZQLZws/HUmoDekT3
IvZsWYuXeilrcvYJgZnNSxCEbsdC5hEG/YXw7rt8GQTdlygSdRS8fKbvZ6NBfaKd
BWsvReAZiYMKdl9DRP3AULT/bz6tUHpT4lumBscl2lJu6loyHBcoL13LQCHUm2tF
29e5IHX6VYSiIAt8i7nzXrk+Ii1/D9Cui7PJdQmlJiUMzCUEIxDkdx8xuCy90+91
Q6ctsts8xGzRSrL/SnA/z+ls8CqVUBbSM8cgZWVGvEGRFfTU78B7oPjeSSKjBUQP
5MC72PgQcL59PvHRqeQCbg2pv65Q+eaA/Ik00R6x8KTzRpLnHywrU7sgETN7LIup
41bh9nqpASoSDq12QDNv8VjcmQXCntCdoRgiFSxKoOnL2dRZNWmIuLi2zSdOnZ3i
3/JQIyffygJJdoDux07EeV3X4G4bzFXis1D4K5QHVpXwOELoJquVNKLl+kZ4U+88
dc+aAFHw9KJWLf7fncAG3lxJfIJPU3yWsNFPeuBqx2twVmyrfZrU+NMKU07gtbFf
AcZYfmRcMVhEuguBUw9HCDoFq3YpsQcGUA3miEU7yxHh3aT6460QIBIa0U1YLaAu
RaB+PipekpOxJ297gXAFMvC09WBWm0sqt8Mur55myMdvTjaKAXnBhd0jrR5bsH+0
A/40CWf61EP/tI+4QCdxl/bKjQhmYnznMkNh5QuWEXFf/e3zjmhEO38zfEx809ww
ZcGdA6WRcA4RS9aGADXU37IYv+phWFf6K6LTKdP3ir7kObLJ4/bk0AF6E9PrwbN9
OeYlHtmlNhlbj2cwOvn0JEC6pIKgOcfAbVX09xpFqQkGsLgiQcOolzA5jTWRT4vK
Q3172GUwjzl92U7dCRxwZzcXXIDWXATfxrqJZF5HI8t154I3f8k2dNNLfijDQAx2
ILH7NMvbPM3BVXOYUB6K+ewnK3R7OvmoswQnwFfXGzXYKujeiQfNumWBKH8ZouwW
uRX0x706xm/ILL5qcDUUHpsCzD8ypg7adKBRnzcr1BgRxbJbHZkpcUVPp8Layd4z
Lc1LLZ2rB7JM8sSblDShIH+UvygUWuglbp+fwUR4K19tEwX5ryw0Isf7CS9B/ICE
Poq1DwGk8wm0H9eIuz0JZNmsoQ9oz8q3wZIEXQNSQuJoOJbyvTW65euaYWDul0c6
M872LwXQvyQ0/2yYEruOQHoUDdTF3q2MsEw+3ihtIdeRwl7S8RfSi/m1VNjZYKjt
zhjHM3v68hbyYcyW/XscfZn2+Dpn/iRq5K95CnZsf7xiNkQb0avb+ANKaoKni1av
N1IQqkVggtcauU6dVvygE+06Msb4soxAwWxLaaCLCLw6FhMDP/sYeXwBkj247rnU
QzJ1kT309crG1EOCOvlOQ0Mgt3N/Oclo1uXiEyvUASfpOGFx+LdYtqJwb+jjxs3f
4NKeVq3/2FLsOIAZFXE0MFgzw4IY1oAnaaptBT4B0+6qx+kVlGAaLuGEutAEeIte
2IgNc39S16zIY1uR72JZ0MaK51Dl+tg/dBDrb3pNWLLds2Cp7+b3Asf38wvCuuM+
8Mw1jiMGRaeXaHz6PHAMlrbeKY9ijDvmQye5r4HagY/RNtOVa87UMRCrVwM8nDu7
YmU4c9nuWkbz6IY5rDhQnOBSWX06coZdYCniSLs1H6tEAVgwPH9VvlioO8Pod4uq
xxMDGIwDubedThHzD28VIFCWUNkLN9+gMbTSgxAY/d+h49ZKze77W/IAvrtQhqAf
01k8GRs9C9mJTSfCMd5DLDgreys1/Ss88Zi2r6qh9fkaVOtHPkik2gsK2kVH5HuR
23Im16pPCqP0FFvIXNuNRgUxd+RIjZD2Nri93hFcCfYl4LQ3QvyfGewLev6YIwg8
l+RVEpSq5HxM3xIuAx27XPOBz+miaSapCkD+y9iYGPF7YGK+Gc98n273dBBSNPeH
kDT85OW/2DXZIGOC5fJaA9DofuU/20xhFDtT1UQKcqGXjgqcdipX2jod9Z4SU+2P
4T9Lx8zhlri10Gpf6+/nD/wvatIu5wPv/dbwghDR6GJToSl23ryfu+WNdTc5kzdM
jlYXdgNGUezFXvEUXBi0D38Ov2jGsulmIjNN6rnme6d7EfnM84AKnE4RN28mcLcG
bjYGF0iwVVR9ZE0mjUxZhYmirkSWdKwunh2SPox5N2Qir3BSfaO8ZV4xLtvVIkC2
ha3lAqnIrScUrhM7uG9DiJ6TBJO4+r5TsxmfWmKBsTyI2LiZjb8QWDHN/pQHbGx9
ldekCl9shyi/8hQQSjAXm//kv2UFQeSdF6qUdRx3nW+1JdTQulxJauu6Y80xf2BZ
AsC33Mhz8v9uERzKtis8adcTZzOKquB75uLFgA7SGxySHMMYE5HPWqLMA314l4Tq
d2wYFZ/MP+LnC/51VaKdw9t/yy2GehQiH4zJYAwZGK6fVQXf4d5hriI8W2ra7Czm
LSwr7ppyq5twiAC2xcafQuxI9hLfjMN2XUbJc4xwjeent7UFNyiwyOerUNqohaGx
QHVZ5gH5Fo29IXVz0+RyKCR6HdNt8PjwtuDgC1OL4p7vnAMYbx81fSZmxCOIjwYq
zDA9Hox+UUDIVZNKT6lxsd1o+1AT5+LljUNKI/Kbf9KU2kgsjY9FnxXSTsteYuML
5lL8EJp79GyVSX5iD0yEmHFmj+PELkThgDZ3Lpa9mdYUXwYxX4lezbbkXQVdBZzC
+utAE1G67NUYo7d+NX6Y1u/tQkoO4DYStbtF1D6q/g2ENfSZSjF8+1v4RzinQwJ6
CPYI1M78OVEIK+YDlpei1oBAkq4E74wZVdH/cFGctbmTv3sRvEjmL1U6qe4kbVhG
jeVjjTiygwUpBnDFuhn9Sy1CK/AjVP5uIUVYeJ6kiIBnBLgUiKysYj9LmmzmJrRK
HD3rE7qypC+ok/hgQazYnL4reDwtRDhg9A6eccGJ8K5x02nOZdVulnEz9TYqIyao
vDok10vvBNmDa5dzvvALHz6gQ/sN9b+HbQKRSuRdKkQQzwqKnFbl1SSNoyjV+XPa
Z5b3+I0uHJ4o7iCB7aiBo334PKyGBU/8xe7lU9NWxIYpXl3u6MsUJkMBvMpun1Yu
0/+1mGtU28ZjHyrakYyK4YZNdCYkg01KK3Zy2Bh3v9EzRVA0ZX9QHSo1gJaat6QN
BEioGZ5oqm51/gggDpD+Z8qEagB8IQR2SAKoLkqDrqAsRYMbATWelN4X50zQU/i0
bFfKpl20BYYAlokCtPAyMktMM1rYB2Z9450BFNtg76X2QEDucC8TiuxQg9SAzhRs
elsxzelccdpPXVC40MpnFxNts0QbhX6d8uoffmdIWGFU0F88Rtk0o+S+U3qjHmoo
5rZX4vphprrFrAXbALlDndJYfXd3xh0VsN1vvbdmhDStcHs4QZKA3LS31guR9ckS
G4LoEGPJJfx95wCVQNQM5AuZyAwyp46LwvjHAVO38bdF3fvmf1gfHZjFf3ZidMCd
wQsdqYNOMOjw7+Ic2Gg70S41dIv5chB5wPCIpjyDsZUza7Vhoz18HvcrM/6btLDI
5BHABQrRr5NhVwOnmNxB+FW5wGNLAGJo8OQwqDHbdhandmvMxf9w+eN2t0BVLr0+
ZxYvVpFVJpKgewJYR2qxWsib6Xi5k9HqMZsKLnz6znHoSqJT9nl/4dYrA+N8zhPw
EYXbbnqOFgPfoRM4eey/CVWFLtnx+YhsyLnSfSnlNhMN89Q3QeKsdE2wCDvtwoGc
sscUUX5VqZtLEGBgdv9U70k9Qi54KcF09NaeCBfz0SfiS+ANTipa3XqOxZ2TmBBx
AnEcfspO5XzTfN0uwM3hjPfevUE0gEDIkEvKh31Oh08C3CimEmnYEjBbKmkyB2aI
YPmGaDNKo32yxWuOJ48xwzg5c+KSBNPZBxXDbfOJpKlBqkiI+4J+byhi8qYPpYRy
E7h1Df21y8QVuFXmBpuFbpyHn60HT7tKL2DF+x+mhgWRfObLU8oTInuuNMuIzU8n
pV66HIJeM8l/FChJ0Tmou+0iWoPzwWwU/J4XYuF8PkZpctdIvXojm9EdxYId05ZG
6t3B0ndpiXZQfZCf6f3zh3s8q+55SPUX5jPwrkDaXlKg4yqeTGi8uOSaPbD4CjzI
M//xjmuHUOiZqG6lXyBf63kxDInGsni/zDwK3Kq8to168H+/PBlkPpafZKm9mkbY
pu0vSQqQRC51886nKyTq4Z27eUNJCd2ZrT5GVvuVwTE3tiQM/DiZAMHkgQXgTdkn
hwDi0c+yf9YOuOQQcEikv3ct1BjTqIy2HYrqRlxCYAF1BIsCEIe7bA/nBiw4JRx5
LgMobYjgAcGpcHcLYOp83GDJbNLjhyyzCrUaYWbwZ2dHIgZVBL8o0hf6kCpPurbK
/QAawdKBLYMA7PuXLVhzIYInhtLcn/6eHlPkIScmiA2QLmS1QUcr13sJf8D+80jF
phlt40CWDnvdNOt6jlre6zu6bBpUCWVFF/TYWH3iTNj6EwlGKp4vzQtw9srKoP8k
5aoeAYS1OmuNUxgxDFEbHyMCXsbBMAP83GoXEHdbgMuhjvEzB4q/T88fO7QX8DJs
1oCPkVih9a4PMr18LCirZVKs/1tUycFvtBhaSIyrZ+QJtkg8OzrSsxmGy7Rgkd+K
BTKsIVkB6Ma6TEesaMuzA39zCWia4TtD82/RQpAuEJdT1Rq0myvgi9wvl6ZesJIf
EWjIM5unrQxWLqHhxJ+d15vyJ4SBXLpVgMNPKBYOGgVMWr7Bzch3GGFSjJjTU3FS
w72GquIdIT7b0VB4WMGOu78hY90phOEZ+5MY0LuOj/np10v/Zd9m9PWYAHL5Bcrp
gLUvCePK5zI11fGXvSqK7OKHKmxfPLSzHRGqION0kvrtlcrOcmt5c4OviNKFN4Vq
3MsrzTwNYTa78vmLrcwj849iWtYN6mIyWioL52QvH5ZSMkz6BPNp11+YeGAT6QQc
S9zlUFCXtPU9not8WlGilqKYyt3w0s0MDK+TXrYIXRJ1AXZxB+aT12+ftOAK1HYL
JwDxdZiet8qvmvJGXHP8x/XxQGA1RqRuDSCwfu4wMHj/iGdOWe1Xxq0kYrv23sWa
6KwOyFf0FemCvM8whAf8hkdfFUsGsMuPG5YQOkgDtlKX1/b1YujDKJj9c0ALvUee
I2ghhd5rpzUisjmEq50OjPgCsCWqqySfbiobhL7K3UFzPa8GP+fMlVrdTc0gghw7
hwGYGZgDcgmRsxPhJ04/HnErBMNW583dcleG7BcCNUaj4JADBCVHBUYZ9S9zX1tY
+e53rh0hWocGR8dUtF3dyM5aBg9gt/+8Xb4z/Vwr1EZFv40BzNyltO79tELMiqkx
YQLSTu/akXfb0W1izn28vfYs38q8Nmz7/xNTg+cXRXAJ5AWFeGTF0gWdXs2qsW8H
xf37fNxtXgg9QKRCAk91uUP2cXxJPkh4a4usyE6SJ2Y44ZKJ0hRKSmr7clHxCzMA
8humBVeBhLshjWGBZbEMu9VqfuVGyGrqI/cIJ5+3SSB5pmFNe4Uec2dr5kxsg3ed
lb9LAavv920Sxcyd8Ee+UT9WHRkZnwLp1bntTs64R+o+N7bAqG5F44ht0/Gv6OyW
dYJA4y6EFze7I3CnNRM7SLMLHZp9buP3P1NLiBuAp31/9eNIFVEnwntusPpdeL/G
rM9FVBuNlnNLLsttqy8mPJHlj8YxCdTcC64gU8YWsN/NyGODJzXldt97QPOX7Si2
Xgn5AmcwIILXF+2m3AR1P/79sobXw4ijN3zwoO0UGzFjiGQK9vCaT/K1tSxbucT2
xdFN1YR/iYH/a61Xl6ms5Gmk1fLoFtGPIFgDtrr6cuWYDaJIBXqxCdKA/U67oY31
PoFA/kIlAeO9haMe06fHc5d2b6hqd5f7z/O4LWCZnfGMU7UpdkHZ3Db+v87Q/Dr4
AhwHo/Slb60/hHpUOaKcaPQLPZ22YUyag+eLdgKSTub5oXK5+1bHFsh9cWmQ1bYh
qGCWEfF3riQ6g7rWN2pTg5Iqai5VU8ihlVJAp0CeKh5yGhCFaCdMCJcPvdnWHhAi
dj/mDP/8hImJFJLA1SaCBIeki6ictSuJ2yHltaBW9cZh5lLqGeZoap3jINvk4jJb
g9RQo+YTgwBvUzdUGfYW/qrPXX2hBXQK04E+xs925hjxnSMXPFjh02H/76IZrYr9
l3hhXazkvpfG5tTix35wlyTpi1MmVIbOW65LbeoMsNxDUlr1d82abGfUbTVmyFeG
4yn75n7Fw2/WvoC+vXYmAn8OoPNGJmVpCs5JhmRlfRl1ka0Azyda2IDpm0ohmPfT
zroCHrbOeN9oKLn/boA4wxl5Ye+Z435fTtqKQFmviuVv70HLooe7hBWCbaAmf5La
YknbBLytTw51TCVElWR1kreotC0gvh/bqdHM4PUEmsIdzpXTQbq0SMTtNaYzVbjH
P0yn1JE+6n2F/sV0ajBZmphc5QWo2sdiCpca3OPzw+T/a2pp0nZP0pRRGTxfmDCQ
ai9PShWwPgun+1XeYZfqPFmnG9QGu3ugnNvDGEQLsTqSgsLcmG3iAtJYkXKEjdEE
avs0MU6jKb9YSNxLSpklSgW1UuTj9FiKWSjYba7MMkznbLkw21D63W/TrTP/9sIo
IUGnyXs8kx//stbb7D07FpB6rYtIdkNiJrAYp0+0BjEr1S8pYo+r+5ijSpXUGOkK
wP9PhB2F3LT9xHmuRaRIhZRT9pX8qR5mD+p7AT9xXpx1llrzigHfWZ7V2I+UfVYs
liKTUnmjTMnrElhenD9d4Pxeb7cvL4GlIp+lg81+TYyDAAnRqr0SwKOqRikUhsZX
2lfZKV46KOtswwZ8YmUD8y3GIACVPdC4ElIGq55weBjd/KJzedEI53gIxRakeD4g
PrCIEj36vz6w4lXKp5x7mBr0IpscUpzJwWiYZvFrmznwxMLDiR2xrT64PPSXF33H
OqGAARq/vNEfhn9iIJGn0oypFrBVY7uUfdl0bwLAM47GZCQ8MMWxNPADOyDFQwPd
A7v+CM4CUPrOtrRsoqEdxr5MKTQuDzyAWFabDeIDZdvxAlAA+pGLPJ1HKJtNIrk0
IoNiVCG7vTG+dKInBjU83zKQuJXlomCQng+JvWqr4C9/xLpGGjSPWaCbObeIZjdz
ads3nFHdk6TKkknnMwA+5iTWC91LNlrohYHAKUekWhjr5zqVR6sTV4WAU3x5o1hW
ZI2SMWwVlLIrGKOlasUap72QepM2Zg4a9Ya/nLrzZIglfikiYMzi2fvPr3LZ0vfn
1lCui2mz3GA+d5Noe2lOpWvnky/l/l0s4idGRuijxxnaRsbXSmi/9JLdR+mjJRiB
4SDd95PdmZ44Y2r/ecDcerQotYwuj6HqgZAaGBNKaygvAdh19p+4wWYhcPfZghj2
d2B/Nk4s92E6gAMUISPl0AUCkjbnjOvdWQv0mG3PQX9Xq1wGgLsy72wHGHWL1XRq
gooOmz1P1iXnGgGP9ZR8jzTIk+3TmXhE1thpXJDt4KvKTnhfA5kOW+zq0Qp0b5xg
pEw+kHHK61gs/eL3eCh+LgxUMYTY2Dz2vKbS40qG2XHWyabEdAJdeuZnhW8vViz6
9aJBXG210pgdCyDJCDU3u0z8oKwZE7BLvi8eHBwp5n3q1TxZCUQ3CnYfDiyRE3wf
iAql8ENqYJ6jn/4Dp4+iJQZYDT6ARJk/cpiRV4NXdVpsD/pruUxSgDsRKsQ2uMhQ
kPEssHYL4eI37T/3aIQtM/p3fp524EiQeuPWfwVII674/BYk9J5yQ3LD8ou+e1/G
nyT3KPnf+eRITUQ6Z6CBbQFy8aG+xzXVZxT6WstKbFpXRUBWFkuWVz0W8zRE+Q5B
nfYffX8jW3fO7osuxTShhxcy5L5xe3UiB5b2Vww8nWEM6U7OTg4CyYO8OCUXCXaJ
e4jth8vg5O4TaECDyypcq2uDQNknDRPv6ZIu26lEEa5sle5tMRk3YDpT3NYek2RH
c1ZMiOswdrdLdeQD7LGaQ8NCl8iapnS4kHMhL6IKILddq9RnzME0KWKZUNhWSTqS
XLPHLmN3a/R4SwxZGDz13oz//ois6f1cmSWQCYvhrJGfWwEqW/3hYRxXBNigGVGa
s56OrkKCcZwNn571I0AqebMmEtQmm1UfD3HojcxPERZJskJHnS7sflrP0nvZiLb/
zIzsebSSaUD9p2CSugCFzsDVabpzXbUcBXuqtD5++enUkMbDiOL24EXo5ska0uYT
jFgAM1FYIrbe7hEgth31qedaxfo2dA4Nd7j4XggR2t+QquT3U1vk6BBT55MIufhj
S1KfGmeSdrbQQL0bU63QvmcSwwm15lpSiKW+UwQBrJ2FQ656utJ9JoTmHBIgkrjr
tZjQBR9Y3ohJ0zv8qQ152jktXZ0oSqBoX0HNiebDL/fsg1KE21S4ixnS7367ZuaT
L3D8AV6i94j///s9Px8KrDi1s5gLE7ltiq1PsUSHX57uTUZw9PTX2huHrPRVfLoL
pbgE9ukXxx/YI7PVJGHd/Bj+ESc2LJGv9hK+JzLxsSsWWyEc54XRqjPORh2fV2dB
0/p2pWFfd2q9GpM9VanqKCCu5nHdNrxcxXmwHRAGhkUbbhdB6EDKvqJgTzw06PzQ
lvXPPAcwVfdI9FOmp71CLqNNs12O5fNQoOWkFUc0n/LlQAG3iP5klwQ+xy2Q2Oud
kmJeUGZ5xzihhhFmEOmSlSfJQqCEJRG1KW6gBivOZGumrFbD15oHWpnW+DvTly3f
y8hFw0f6whAWyYSRIo9as9s7YpXUOOVtSjHO9OKl3UZuS+UGevojJSlVFINAj2cr
DQGP0HkZEWB5Q4PXQDGr54so8nS/Q/RE8vZo/J9373Pd6d18w4LjtWg4+gxRwD0y
DwBbZi0kGx0tczbocDEUML/8/I3hgd2sJMARPaZxqYpMVDXS9Bklua5cgSliMphy
SDfrFuN3iZwZf10RpOeS7EmnbZ7NLZY249BEgUOre2K0vN3Lm8B2iAvhOhAmCRHW
aExa04l8tqy/BXVCh3kksFvk4ee8cqUTBNGnHaoM34+cHylI9ySAKRPf9HKhGYux
dxiM11HMPRqKSbVYeB/wFl5Xr8fOR50RKFhbtknyw7WTONgQkqz4NappzQj4w5oc
E983aX0TB/7Un+Ohk90kyAYeQ6nkNVXquXOJCT1A5Y+bBO4TnHgmGFViC7m+cqx6
2s5WCaYRlxwiYGUPLuzYnOWpfWig2qMO9gLHX3CntWGMuf1icuIaKJLp7b8i1w3T
WWRnWQqUyimM4Nl7g61ZCwh7+1WrXo/OaM3evECAkwVUIh+ppee1XqUFVZtBi064
sT23zx90RaHcK69gR/+x8rLsOEeVrF7s2C9FOP2WjChb4xE1nEBO6eUyQSC9DWOV
HBaoBp4TsUyjE2bUjBYF6yNaw1FixYVNMTpdpaI2G84LJELk1JBvc0O/3kVDPfi7
KGFNiib7uI9agF2jIVraaacsXs7HHnkRfBpme/9L/o1fl86gEFDR6pZqaavxZNPC
XxO2PB6391BR9ds/La90tcRWQyOo5zIRYES9kc5HUzCcLNFLX7jr1QqTIOe+kfB8
BVKpS/mmnKl466Urgev22fozWa2Mo8kbnZWBgZF0ZBUn27MShk33c3CqndKoE7E5
UbknUFm9pea9HMSgxJeRgEIgKhTDVqgEOp/yDhI4k4b9s/5r0TPPEVC5Pw27VF1+
yuNvA1cdw7F6vBdQqXaH2wbJjSsLTLmrNnZZCpEfRqIPSsfQnqGlgioebfluZV0z
SOoGa0uJ323P23r41dhL2zGurVggQRRu+A9MRnNDLshYL+Q8e5jRZWg7ssO88nSf
p6YRMr4UkAIfH75etfq0rC+6SlqADSKsVeFkvviPQVDosYrjSKn/GWLUwNkp9sXj
88l7KxxP0aSUAzbz3o2Smn62LM/SmQT4BiW2nch33mAaEoBZdgHFRb1yvL6aqSaN
5s0fEu71LEMx06J7clTXhp/MRUBAUAMTq1OULCxB6BgS0KSOGdrKWuIi7tZG6tVj
MxhdJ2DpsK9OUWmDFeg4hpoRwH6ROLjCDEaleEO3f2XgFhs+N4wvSMAiqGrwLxzb
/ImbtapXPvSS7byTxj3WYDLDBkpGB3EDmCbUpwIKfU55UJA25kD7au+CUUF4q2Y9
W+bhUtby+SN98s4ZPjnziHkttYGvlzSw8iHcKAbOeK/PzHJpZA9BijUwhURKdeZn
8VisWorfqfTVWDMr9Zqa0XYNaApcX2qnVhK5ZIgY0vMDD55ZoT/IXcI6wcoFH76r
HG+7kOsvdfs9iUOIcOcocNlshRwtStBvewiDjs/Bb4n4Juwoc0CFy9ebtyyiSGhp
j9Hhki2H9WAAvIVaOGe3pQxgNmkncFt3BXCoFhZZsmIR2ZsUQt06l8yKS+T+IcXA
DPpJbBvnk4I31OrdJdh07Z6VYJa6V7dRlpxhw6VAdelyqbAYExEnazkp1EJ391lO
c2aFMpnEG5RvvvWLKuXjS/CNHwF3iTj2mNPjPvIYKLM/USPJxj4x/0LfzGhRPjuM
gKCB1ZWjqv8PqpzLCUYiMlOX+4wG3oM3CkyEY/hQMOLm1AHQ+jOVVM5XqAWXBHWY
tXCsIUNiqe0k4xhaYtFq2Ok/Ozleho8P4a1qfUl8NXDkSyUIPA0jQMZKKYh+6ov0
CkWAyhcEAMUmdqVXztiavnOfxaToeA8P6KpcPsSsojReE06Qajw0KHCc9+MX0L6+
yL/jHLdQnS1DE7WlE9swecJvSMRctX8KTK2nVUz4PJA0P5l7FKX3O6YRcKU+ofrg
cKHc0ZH+OTexHh48AOfbxNnFD4rrbCyOQS5/Jc2lQ7llZ3LeLXYeXEFS35QJimqo
VeafaQU8KJMtnZcpUlbpnOEgqGadupknd3vlF51C65i/u3eMArQ72/+lX+7JmQa5
t1R9T0+0Daqk4L9YaoNqt8wOAlUiliJbv5Q8te7lPdbEddbHm81Hq4l85+v4aZA7
iQhKL/rU1pd3HtloQMb/5rFbYyuXYumxO1nfLoepIYw4AzfgC8Q6tzAYmA5ID0gB
1lKGTfBD1JbYFyvsl/OVpktxob3ax756btY8/nAVkCub0kXNQ5Kwnn96oUMaXFFT
ctHNmZA2pc9HM33K/GOmkKGnkKl4ne8AwgVWROtfaf8y5EumSH4SDsUa5OB7KLnY
hx5pEbn25LdrvZGJLxo1ZBp9c1mTvxrn9cUabmZ9N1tQ0H3YvAfhVq5MYReP8I9u
js6S79y1qvXLtTpYHS0row4LpeKS2nerK1P4uXjhdkyxyC9yUhO2gcigOlnI7TQB
iRNfRLFSiXyB/gQveT5o2M4Xme93IIIQQsGlzlh92ocpyt/dDUlW8OjiETFdmMpd
95ZM1HJ/p15yLGL2LeYZKCH5mD01Bmi98wysV/Ra5/e+0gfYNGYealOqva1geM4b
jPBB1ci/h0lS2VGP8dD07DgwQIljgSROrDf80mKi1+9UT4GPzR4w/EA+Hd1XxYMF
iKjSt9p7tcVx8LjxaTOcvjNCft7D1x/511yys4zWm1gWys5CWEy5DMNebAxANzNW
tCWlRURbo1E8UuXM33BTd2XbLvI8cs9E4hMIqxI55HbzzSKDbwVsp0CVFiqR56Q6
CtggqWyx4in9d9+QcfOMSSXncFnYx+dKXRwjm+2Ulob8UcZexFBohXJ9c5octAfX
4QqhMOCdyiFlpZtPhIrHJjh1aEthKwVWNhJV227OLkEZF1azY8ECV/zalrZX/2pN
NkiNwF8ut+d510+hud7McQyvcbHQZD0gdPxW8ke9Q+4KRKi5euPkgVq33Jvfj0Fs
FlvY8UJb9U6nOnM9HhD2MFtb+q/UxqnQztdRg93fT9iPHV4J3RwcjvSI80v8m2vs
GtZAyeHirl9rY5o2N5EVJt6YL6j6Me2mp+LtPWNZcbphNS9Ar0jHEYBBpyaVE0lb
w96tXLWfv1KlYiKLPv/l5Shz77VL3QpBb9nAE/A6I4tulR4vyLCLRN1Zd2+MOX8O
JNbtjuJqVZxolkQLLOlpwPee0T8pRzYbaZOlPqhxQg9xdzhn873BDY54+Ae1ogad
30qwKKRk4NDTaLVS9BIN2G1PDaKaET6Nees05+ZWkNGUSpfvJEcgcWBpLTnz+Xx/
NoWAG+I4dxZDLqfmPRUOcYO2IA3OrW864pZ4raTV3N6mA6hxDyG7/7GUeh9/4BI6
CwMyhsJa71tmhcTy3fnL7pDeWYtdj2UfsZvllQXfGywaRzyRsUFhgDypMyXsb4DK
UYdlszzERAbAtJmCZHaNh2iooCAbACqS3UJkY4IeOy+fGET6wF348cuBwgcrAweM
JrTsV3uEXQLvBxfJg0thXGqlO5TeJJV5ftYrZdJhoXMj9gTP79v4SKX6qocXnuRc
OkY7tmtWbOIACIh+/dUvhGfkbR8sqohItEM2WKjHf6Nf6+3t7YZgtLazwxc6H5jy
jXcYLZWZoELPjc8VBo30JM1ckrxMUQelewBvQLPcZ6tttHYwOZKI02iC/V12eyEN
tXzMjLoaQ6broT5nkhVKnFKY3wQv4wRFnz2LJf1WgmJY7l/V8AEblW0q7ydeNUkA
BtyDmPDFgbqIiXWQlovll7AFnAcb183niiuCPfGO7uZBLl9BNS9wj3qAjYPwYO72
MYSsaOHjMKItbrGrB+eh21LG9ILSuFt1AsttKUeCuEaxYuU10rR7DJhtghhTD1Pw
P7inJqHs5R8bJY8LRPRrNKaV7eCZAWbG2NlIQwmcMehy0jtvArM6Y6YJ/wTwKBE1
rj17a7N1JerlfLQTR9DKqc2P4UjGfoHom1EAaiwbowZFFlrLouR4sXbFJz1xY2hp
KYfjdG5dXhD7dmi8oSwBtIn6b629rAaMqnalFCkMBT0kkHgNqkeShWfU07J5GM9u
1c1XHx+jD3n3PNGuQgTh650cKyFIqD2Buj5WxpIKyTABq5SUp3P7zJ1p54QPNpe1
NgHBgOVZXGgVJ71yLAq4i3FoC+vhEhJULxIqvrscH/jjUtIgcwmXNvqx8PXiZmUv
yMO+1DDUyjCeuCNQPag8nzjmOASP7BXFYrO8g+XksQdS++MtLv51bD1Zz4VfPhBV
KdxR3JwUOy2xbZDRzWYTMgOB5spFOZy7oQzKhkkj0KOL8wvHdYhVZ/CLcWuZv0wn
IC4GJA9DD6tMeVbSgdbhvvmt9n7/0mFqet6WNMUlkNdxsyBJpG/xG+BjbKiajVlQ
vLcmLyciAMDQt/ZG44zxvtfIT9WwAGrGQobVKOW09KsYi6rxmjRFRU6wAbSEcxEY
IPGopaKuIOYmL/AgpDEMuGJ71cw66BPxEV64F9PWWEp+GVW9AHH7UZpcXnX8HuAW
jU8zG6Te+ulq5U7wo7VpnHuXgLol7P4GpR6ZGJIZhPZ6njy5j3t52VAHD+OKjAsH
Qb4njYBSpyYeZ756gZ6lQa+C4GH9h227Ckik/yerhLi0RKKBgdfSgP+WRrCSbIio
gDXIrGQh1rVVaMlMg4c1Z0u4gvjjGlL7R60Tbs3QcQxDWCx7pCKM6DKI6zxB9inP
q9kHPArvp5eNUxEe7wp0LHDOmrJYkN+1coMIKcNpmCvM0dBXIElOzaj1HFW9QG9X
IcbJa57GYR4WibE7cna1AOsHtozgPFWVyLstdRkchVTMGSigpxPkrxgeDGaREeuH
njRKJkrgPF00+TZ6KZ2xMf2DdPS/NE3GXCEFDeZ8FU/x+SOsi6Gvzb3jO7pN8TTT
3C5iYLTGrVtN10OCFUfxtytjzmKEFHunnVUe5VoOvfwkm8yLvGQIWIEZ0n6z9NdL
rjdaME+0aYdJddcESMqiIINatQHayyyHaS73Eibq0/A8kwPo84zkxBjuzNAdvfwc
ikTUCFzLvIfDD7TSYqNFADwWZmy5EIrVlXB6vrYJBbmggUt29LfU1tYgnQ8/vISU
qz2I/qvGvW55jnuVkmQBMVO0UKIEVIT00ku6BymIYrRst0ET3+VW2M3q0Wy7Ta2t
c09sSTRyy2L9zJE/WFZZs/f7gEQhjCaXzhUtzMqEsDulIE9ggee8OUpCtRXe8mkM
RAKM3AJ0FwRciZ98V4VKYV+mSu+t0uYFGGZ7yMws18q87HgW0fULdWvQCx9RcHW+
cDnxNHxKAVKhKxZwFAJ2KrT+MR4pNORO9FqqPFek4OYS/VQgLzAydLDYnbREEcnT
XHoKt8OcyfpiXMblzlIHJ3/MvpGSMz0YXNHjRfyyeCuhDW8mcBoUe7KFbelXsEiF
pLpv1HFxJe30xFJF2aJdStqULvtIhV6EJpfpBPWFyn7zQzVvb3ZJg83pzoTRRpaO
rlHZnZOPNCsdkn/E/ArFLluSBoQzhSFTxwXd6tq8kj7aRLL0Pum+wPTA75RnNYcm
dtav1QEoUSXE+GmoCrjaWvdgNgVK6dLQDxAc7v+6aOjHtpDzT03BASVfLxGq/jlH
RqOY3lpjqT/12ztJx9x3cWWqzS803UwpXC59+VdFALIlApC1OZU5vjs3U6Y6nyF0
03aq2F9aEirrkkYjeblGElQEjzOLRrLSpUuzsLU8pv9mvoUkMY4GzFdC28YWg+79
tkOexdtpERQIVguI1vJjw0GOnqNnNJCQ/yTEG+baHxjU+kNJJ1HrJOSgW7DOWXIK
ErJOOvfOyWPQL8eovVukemlMmJNDmEXIAbwX+3mdbmfqWkV1YAaCv99kFcExGBwB
SOdPqUgMblwxrqf8/v/Dc+pcWYxrB42lOjfbaHjn0eu/TZccIShKCBQA/MIeR2lc
FuiUwKT4fDdU3U8kp6VVcP1VCHWFljvT/QWtnlmv/URK83NR3oSAQaQMj8Ov2w9l
oC6/KWrKVSdN0Av0GuxXIQeJJwLHWb+7E5OvAtWt435ME4hRurit6rIR9/UDAhmu
WYIK/xboo10UpDcjXgnsj7fm8eKj0G4Of06pTMt51Yh/4Y79MUdcTRRpXcmzZgOU
9gid7FIOyKO5Uln4UYy92RZdgZLYNG9JSbpQZFe5lr0ttOYu2Lz40cO3XVS8W6aI
uk8SL2OIBqxsv7BsOUE5aZavr40DtuUgr78QP8fEFe958eL0UzNhkZpEO1yKFWlZ
KkyjT/k4oD5CFb+GcqVb8pQQo0gjnqw2MOY19nPU/BWMhW6IjIdkoCm4Vet0kUZM
YtVh1Ci9iZjbefxzS3NxF17zoEm63tQnBwJNxP4/dtL2edaHxE8faf54PO5WZ1Jg
Onq+O8F4++ZkdOiXi36q+MgP4WCtKUeNSh0ccfsCZxbZMsSP8RWkun6xJuFzwU/E
0Ws73fmwd+gYQFiM4ECguwdlWvrDDhyr55Io2LtC5aeHgLoFvOeC5oGDMDgGbZBI
Gb9E7IvKNUuQDfGs90aXrKd6/ayNqlcdWje5agjcHICYan8eYHWX2KojqN5GWiVe
0oRp/eBT43N9iwpcEz1TLoiCDwT3ySI/WKSpTLC88+uUvss/zGuN3vM5UGDsEf43
76I9Zdpcu8FSd/ncgL4z66iUxg5tbT8bVVNpzvhFnuGfz0wv1n+tAcULI/QaVamV
vqbCjqjHUXPTtZKNQz+VoRQwEmUrbWDwYf02AC7s/RSpDDqkSJs11gE/kibJ+s1u
8CaSOdk55mB6L49ggPvZBG0YOkLNKUO9deqkQaeJeF5F5zcKzUP4gAK3qy0L1aLv
Af24lCW08FB9N6dYwZj9gPXjy2q6e3I8fCdOho1BKzwku29T8tkDhnyZ0lQ5bhVE
lnpJaZjutrZdGeqVSwjA/e9isL52JSZiGzHfDjJKw04ozdMeN0DA/FiLkzowrDgn
QNdOr6wXbpkqoT/y1VabkwkEDtxB4bm5h0qfNbqMh7fSP1z+3u5rhxZeGX3Htwf7
soURok2CLJU3pXkjxvoeBwaKINgq3e+UY+I08b0b16t1eojkHiVvbPkoOhA4L+Pf
TjjbczB1wn3HWA1YUIA0TvPDJEumlFkYynNZIht0rEkx6xI1E1YkJrLuTV9Ttbw0
W8nvVwkMrJCEzm3w2M/NxpemFVcVBbRnVnoDmrH9AD1nJLO+csWkCIsMREjPHy0a
XtaNoq54nWNN1VXFuvqwUb54V40bVRxTwk8OaLz3osl+nN2Ov+soy3VCKn9l0ZsW
4br8rERvZDmi66dvfBknXXevlKt1rHP/ASHlV2AYzmHAeHdnQijylXOMSHdQeTIf
wjYU+8O3lGn/vmYT+JKBUgmU8mZPfbOW5uL9AQHtqUmKL72IJWEp3n7LhMwpwWn6
e/oLxbWAG1kXMcK4U0IFaAghmX7xNSLlhRsr1gAnLEnWnia63klWyY8FTT1ewMTa
U/IS9UTT3lIw4Ty3f8BVO/TYN6uPwoM9Yb5v/KKGZCW09m2U2PM3kakDbvQHSEfc
fdxkONqQPldiUPw5F8piRzLTZmleZMwXbmWAKcn/Iz5iG+Ga5XxafLmqBzHtTV8u
7CpcaOo+KpzURADE9t7V6piGmMSXbzVoU/XiagMr3o6zyNnTXqm6WcPWFT+DNpMV
WFD6f0UlSCFLcAXbT+fVXLPCm1/DAKPqbCzTwcKatQZmnDd5zYqZ+JtPWuYzS8uQ
ShDv9h/WEFJaD3ef3CoA/qdvQYmZWGuZUb9y4zzTttOWvM7P+Rryp7rb5p8QT24S
VEXAz+oroeLrdZ1ok5ckPhR49kSRTBo9EGxiVGirR7pyv0EDhEipPzPwcLuLzP48
g82m9Jo68Sm/FvatTNT2DoNEiBmaKnS0FsCQ/E9WJ6+l0L+XpuYtSedP9ZnogH+y
f2iEsYwIzTPx981lHgDptIcfndaJwbuGz4yyLzhbd5k2b1EaIYK1QERIFraGAaYd
bDKRpCsdzWbT9u+O4hAQve2G0zEKBBcgUDgPtAMZFqfan+P+IlQEvbrbBTZEPEyv
aJhvkvek75AJxmzppEJNvd5mmip3D2teGTyTsIIp6WJtDNPDmlo9tnkVmJ8VSlUx
yA7cyIZKZrms4pmIzLr7QkNqOrx0bDQtF9+CbKnhXZ3+RepdXbyl2Ze/80CMEex4
jfW2cYoTTt0H5JYW2ailGeHs28pAftYXanTz3sPsO3L2dR9fZLq+ggguBb/r4O9A
VWoTnrEC+MeeIOv6Ucn5o6NVtzo97clbTbut0eY/7yrKVUN+IFxLv+3TscQnfNzA
+PC6P04Q2pHehQUXYGX+5jkNFv7NH7ENqLlWlNbdDDWs3pzCKBuqSFmsui3sKKo4
7YI5SazkArRgx4wyFlvbiHPSHNfehxVFaxCzPxrarDyJx9utkn2cJKaUWzhZueQa
4yppmI8gaFSlIlW06x02HszsXF+15ntDchvv1ygE2K1s3fVk822ULrkF4jImW3fI
3qWzjXkrJBCmMjCvKAVE15WSLL2XO8Z4fk38SJpyaznshiB2vrAdm3Ic0RP5MjEG
7e/I5p98zFykhWi4F8Swg5tv2r4pazE7kSfZPHpkR7tCYxPY29jMsH2TtoEYzH6Z
09YKEfNexYH3Zhu+Wai/zkfTo9AcRbcHDR9ogvh9i2Fdxy63AT+wLPnLeWxfOPQM
vPIEozFSFrRJEZ52fPOsOGmXRYgn3XHjHnaXHpwLMLALth6xVRat96yRoqLKL2zB
2ZFBLIwAf+MmCpj7RBuqeZLUeH6tMMEHvWisByP8nKVqYluYnBWRf3B6tLfVj70d
2BPEwFOyAN3UA0dAi/SYOoOVBK+RmNRppZprvq/Xk70+tADZHvVjD416jWeR5zQu
uvcWN3rqbofaWgj2BjWZysU44zCpkLQGfgYXsauICk1JLz00rqdNjbPfkbTW858+
h947Nea9l5UfHmJmqBQc15IRYQhhSBDDMDMGNSXzRwnLBs3W7p5NGjUoRYQ5EhFd
Z4J6yMiEt72zYfWYtHPKNhYfBJtQe9TCMrYTaQoTNHb6yl+RR9BVjoiQUVodCByS
rqytXuU+aYkJLsQAfxzv2hV6UsfsNG0l4hmBRj1ZVYSyh3XYXUIdsWxVnRVCg7zF
2cJ+Au9dYYjR5nNbra54xE/5VJNLopVTGpy4IgdSAkbut3qEG3RLk6s/PGVbBn5r
kDysb/Km8QGZOf8Nde9izeG4ngI72KM70YW37FFpTzsqke0n3SSH+9fH8Y0QFCv2
8WM2dH4bQw4df3jbTJsdz8Jq6c01V8E7A5uRkqH1lYHdJMNkIbtkBfsOevRYILHt
q/c0y0I/5BZSOXGkf9spVP6Csfy32xfvt1Q7Wrkyk5Ly6RPyhDqSfFPAnI8dwAI9
53Pvt4A7rMV+nqKbVXQP3k2SKA2Lc3Cd67FvsWiFQc4OlYSfzdwz1tdZ/9g8IPDL
IAXXLXFIvEDNdGO/bY2BxgDhvUXgTwyOrg7WRvdfdQ7YiTYKaOrDsLdEYaABURSu
NzAYYv+FxDwg35cLmn7iE0zI7RKV+PwiseVvf6bTyis01gV2axRSLd7VZvMUvTx0
mWuhF9BmkehqaOU2/F/zRwSwsXg22zmdgixwxjWqwZHrQ0cVDUBChUvkMMzYa/o9
5J0woqO+V0oG8EznFO1gEAVPMqE7pvfiQERyrBMYQWNH1Z1L1U/jYEo3P65qGDXb
7GFpY8cMvaFFPTisAYspd0Fjrkko30TCEC/RUiGzH690B0J1JbLEUAnNCuiXc5WM
n0bqjuUshXsARVBVVlYe6CEKigKAFcIE8BgRAzPUUUM8YEyten3kJztfc5C0sRXb
r4H304pbW8B+xUWK4Hlp2m+XTWtTZNHz2T+i6hjTrQUBg0axMfbZAVFHbdJ+yMmn
9gSBiAFvjJXmNBM99JJsVeqfj+Mi2IlWMsWmA5nDd9v807ddREx5XiTqDABnvV5H
bzxCBzjHOYW+risvXIQaD0ZsJgD7FCeMwluKkujcWHGyf88BJrSA/tjdhEA6xRNy
LfzgAZQi7pZEIn1ooE7NS2Ts48Ad1rqbd0uZL89b5+mWq66je3Mtq4AFNrivh5CA
7p+4tH4pKytouLDUu8fwbpyWKZVUT277HaXAo4G7phM14ILBreJOXgLIQpouJSWO
9op6x2w6SovjZHYtmCD1K8uXNJWoNyIywYj7br+Sx+6uqNiAcGeiDk9xfrnnKkt/
WGAp1VckDZpHeNdbjPs4T/pSLdhKV18/W02Ug0sbZhxCLUyC97CYhL1LCH8ukX1O
T35AtnqUVrN6ROWpc7lAM1vr8hrmaf13AGYY4uHq7ndGIpcDj31f04QumVx9Chzn
3R5DUeY6HaQYWA/vM4riBlKkullBYC6xGW1/F2ATdSKydzU8mqBIJUl33S2cZo4a
akLWhsRl0hxhPIncT9y3a1BtEAHC7lrwYWsO2E5WcRrySHSOLnWt2IvVO+2JnJVc
3oL85XF0HToenWfLrkbPf5te6sRGT/IQkuUwsMaNItkEwxwdBgAnC9DrP5WO0POv
dDnkmSijDqu6NmWA/XEBj/KdmQspemnlcoNYavYkx485cpteOmrQQDcuzxR+Z7Kp
VAljX0MD3+Vm4tgQAKUnsNaRBAnjzxI0djs7l+fUTwgjBfFnJUzkwe0PFRk7md4o
z3oyctvIomRu+E4DJk5TdECKc+gHJnz+3xhmwLe9sf/w3ydoTCD/B1jnR0x42HNC
vkywLonG/pgugqjSqC51LS6boWeog+5AP3a8MsXwJ7YZEbu2j0+J4p37zB9p1CfD
jwG4KVzsU7QMPy+KnqEXiYfRq5cre5qt5E8kx47CDJQUxuG9NENMUt/4QGUJmfXQ
z+h/HWggDvedyaY77+ewT9JuVeSbgORXw0HqrlyfzZ0H1WPRsUe2EahAL9NJMERd
dELTp5qzaQ6AJy4yh+6yHm9ejcNrRblSYgcZtRJ1CUMyPozXEC66UxfBQu4tqowB
/tToJ0sMvslKuixTm6mFh/bENHvQutGO7d2zweHriUGfYzlvsOfoLvtYGeaytCkb
ZybnCmk0mNYt7f3WYOygA1PaBB9HT337mPY66BvprHhfWG2wMNc7k8bKOFv/Q1Z/
XTVwrUxe0izE+anssr3upmyGhgk7fYCDiDCl9zwZzcLhKs7Ew0WvJDs/o8wurFVK
xjByD5+v7kYizJErbWuKkoALvIsNhSolr6caiSSJCYJbHun0XcRXLCkM1BK0y2q9
vI81x5BYTL8/dy5kOi8HycH2Rgywm0mn4VN1H7Nrv4jHzdakVCipWI5Lsq7BpTlc
qqpvG8r13ifmf+s2zP9AHN0owyM/+pvoG71gNa+M2uRwRCiuFH4zuwDdme50uV6U
FS+JPj58U0a5LVZKaLO/VNBzcDu0uOd2cTzLrst5ehhwAhSAEchGPsFNLL/d8RXO
iIvKEwPULBnM5RxUhKfvtQFF2mqNZ4xJ3Oqrf0oZpA9PgY9SeUc5QWQ/GPdEm4Ja
jmVIopQrKM2UmtbL7WHS3w4qVoY9Ja/rkEAMc11kdiBQZlyaal016Tg8xG42iAuU
6mS49lTFLiYb1TrFiSq/1H4zpAE4OFnOaiygfp84O9KeuZBy1lw4yIRQ5Svd4YTC
dA2PcRrSeoVQEvCOheDTrYs2Vq604WvD886iNCwoLThCrL2bx0sGs1kha2NGB+As
JxGOW0pcLMKealCY1Ekb3O/MUmo6gj9LSJ84lGmd6y6m5TzkxZb5IAkRc5JWF/qK
vI+JXJmBVhkgk+te72ev3MX8Dcz3deJaZYZX6v6gtAZ5/+NdAnyx9GEruyIWnH3K
7dTrMYQ0Cc1N34clrvxafSmbq0H5A1D4vedjcJ3mSozDXDqTppuXua7YKyqBSerL
3vtn0Uax3XSxK9bTFLLEcEAraEOEGu8Lc+k8cP3Kty09hsWAwvLZDbRK7GoDvg8f
AdLtVFulhhXgy49ld6pIVNo8OtFp2zKnx2iyjuEsNUN+lZX6X4aV68PVGZjgDLoj
/ocWHG2OJFiWC/0t/b+vSPBNS4QeifL+/RjrJLSpOCfIRHQx1fZWWG2Ogajlaaay
OuOZvlruXNPcdZ0Fn2Rn7sc0ATQ1WAe+Sfk1sEYnnudTU+VMm0/fUkbZzaZrf94c
FkQx5hQp1Ssib3Es9AR9NvLXGxhLRrXS2x7F0CZEITJss+8j+vkF5vDOfLVq02pc
QcpDzZUCv92I+rfoRJJELxoG+gnDUNMnv9NevVV7dU0jxdklj5NeNj5VRrKRIO2r
HuWQ1LJ6lrbeXIbLGMb8biWrf7pEQQbrOTZ1kOnNdh8Vdx9xQJfB9wWjfrNChQHf
vGGPVO8i+PsnwXbPRKKtfTGzR07jhcTnJUfX1kzpTNnOqhs+daYWT+28gqLOHAli
ovHo7nR0e88alTIm121FNV0uCwu7s+nM6Tt2rx/9SBQsXw9n/D/8xSaVQpgCUNIh
CuMtQ/HORBaG2seXEc7+qMQTAeOPL/WSOzRj5oOgTxyDMYhdtd+2fDqTkF5lrPfQ
ilgf5Ed8uY1KhSwmpM+3zFxmgUWDzN1PdKQIWNcEzZUa3yGT4AfZMW4c77ctHQK3
TXkLfaKP226M5pKxQYsZrKZ4f4sOYw7pbTDmDNmvUcybsiwypKTW9u5RiFstER3s
TdoHHZ+IJY3YnKnnV9ejAZqgrx5mF9lyVUVS+pRZ8ZZ02FMkjbisijmGNeMVgylj
7b9YthE4S26Pte5AyKM7X7LyDAKSRucI5nOyaRsUfxvE0qPWNeiUCenpjjO1Ta3Y
LHHiqXyKIx96h/ZBzfRy4nHLk5i1wVAA78ubGOl6/YF1iFsyOUKlGyEA7fq27rES
jC2/0uCC+O3Scqa0kOz7uVmD6OsN9kTVgjenI+mCOED327OcBV75rHWKrnIfjT7b
hmQ8V4Oz5mMtchNWoVEW/HFW4mU6jmgufH6ztGkzwqt4lEb8i30GayT3T6XtTvEp
rQD5nnE8BjLYSI2DhcLt0/B0F1juEvEqsyqi9r2WoHDhnvsWyXHcvzh7u6FqbVO9
4auLGo1LmnUOA4qqOcl/pbSn1JQwrUTOp6bQ7f+ED1wurhzsJLR0iDHx1fY4Qz2g
7mAWo6DCc3Fa4kZiGkKethvobLw9R5G6V/9JCSTStl/qeyLFTLBU1rbZ4XfQwiLE
JhlCoRoVOxklrn9glGwpuAn2nLDmck7G+/JiYWzpUtYxbrLUgo7PMRqymmoL21TB
B5u9uLqPu3aVqO1Iu4RRGYgSKxx3TY7YBbwgHIcN4JG+5f5n2Kz2knyT0pLGW43E
p09f7B477o9IwAkXewNnjhRXV3DUj3UJMXEvdgkp0WyMTlru9MtJacS7U8Q9WPZH
OWmUdvTxOf4RqCc3FSzyosCvV0yrJzVZwPIQo4uptahxBaYcEyP5z3Eo2Va6flW6
LwfuMP/mHfEizoiXxEMvhehgumP2JUikakYAUArFUEfm6H2ZDsHxdjh2KLcto5FW
VDpZDwdJXYIIKxjdWDIUsWKSFSvx4zTAn/rg5Azj9od/eV7cNh4md5umAerUmofb
ePoj0h9PMz8wcgBUbC0pGu8nHQ7/YTqr7rctRgZ0QfjsPMvu2uAjFibARINxMBqW
qFv/Oc8+FaiyGOA/c+mAfqqDJa7KaRRRHHxb8VyEOy8Doc3CtRplP82iAaFTbCVk
raQSbTcDVzYLpmTJm0QePbNqV0RqcZWJTrArWAIbqsqJ+LxvaBBNRunH++HtKGWZ
6hnlC+PJVKsrsunfs45iGtVYgHzPvbNYV7GMCkC2to/vpBMMEqCu2bJ+ul2gHfm4
BiiEckoL2pUFStZx7Y47rMn4MY6q3Y1ApL6YpKMvEjgm6is7skFGjLcYzZHQ2q3q
w8b8njpS4SZcrsqpkweu/RLhb+LV2VCWRgU84uASFzZL53FwEG6Sjr1w26UslQYb
OAMkR6iIn/8HoChXqUUSxPwfPMHAV+/pTg5jtP8s+RyRrxgAttYbrJVH4s6wajrJ
RmAPd6TR3Ak/ticGwZO2/jPEG6vCxORR6sLeIuyuf4bCcxmu9xwT7wioL32GZ12p
CXDvTZz8WqNJlnAKf8JQGARvmV7dKkmeD6ykHAkBQjqBSCKI81GcPEs1S+wGo09Z
a9iO9NtHGqkSzOE3xt+ppha6wNbEy8VKbwEp8EQvfdTMOHoDg+67dd3GT7TYrvQK
VEe6oA687GnDIkxEhK7QJ4kZDBHKqbQJpyadP1NzktX2cgIJpzp8jo2gKe0QODMh
HW2wysV+OQRZ1CXK06VMDw8HVedwk0m4k7iocbTImsCm5ts8LUSZQgUXrCRhzdRX
QLeed6mkiVVsn2gouLfOmYmblU7C1xvc8FWPcIhyVcUfEdnxaHp6W9CA8GqVCZeM
r+u05d3+1OGpybAq3T7f5jbjl+idRplOWpbRSKOLXbt787NEq/I0dmqA43EX6YSX
gfCMAroCWGrkSKCGeE/JEg0sK5vFReacL0EIorTKv5y/digNstYE18CXUYuSiq2k
Qpq5/RIovAMTGVeYSA+EIkxwvFmtmGGCi4X49di3DoQk2+X2EBruTrHziR8ni4Pg
RSyw7VFhtPjDyiTBBu2DKerPeq+j5uXuSA+/inH01lldmO6Vzlkjs85amgwzldeD
uaC/tVa/FphhaRNBadyktH0vefhdruCDWpK8ZS8xm1faqHyZbUHUBA9cdOFMdhfq
3UCl18ArofSop9sCmIcGwW855opjTzb05SDHj0llfvLLt6AP2TjrAW405yO20MUA
Db7KaRaLz9XvGD4jBmZ+5V2RcIgdr0PI4sbBredwIlDmqGylC7Hhd1QYiezbMrFw
wiQ2aZOLYAwMy3F8b4uH8xL9+DL5vjBfgodyto9z54ffKeoml5U716BwjYCzB1Uh
WHHRE6pejk2/VQn46amrXww5gOSWngYt/TeN8slRyhNhKoKMEyfNslwQ+jNlRP66
ymXrc8AexyitJBWgT9qknATyerEyNR7inAOrsnMp/6zobSikO5///UPG6Wt8pB3b
ZMoqNWvdN723oYCQzpAgIsHNCNUrz2RkU0SlQGBvnYIA4I+4OVhBoauC8N+1GM3A
29+Tku76NYi3dz3xIrBNiz6vW7sMvGdJpmWM8n0roliH+C13JgLzyyJ1cF6EAaNc
4LD77dhG1SRdBKowCS0Nomq0V051SkPuB7+xbz++Fm0ktv2P1jyuVpS01ZsjdYo2
UQ5Cn2KIFXvoL/kUkNOJ1M6qxhHknEC5+vKXtCcMRlzRWYtDbSe2e1bJ7K7b5ZE/
EV+ZigPo5BuPC/ivvSNLfBRYSh9lgtH2VxnLVtKXA0feGndmKxAiNYEnneLTM2m8
1nbE1oSKHuco8i3Ft9dnps4mHvSVet5h5xscqkbNOep4lWJ/v58N1JAPD6rBqp2c
MdgjSPjVS4fVF/aSY4d6ko57RaKggMazp3y8tkTZ1dWk1F1Ne1iDsFw45TGoFGgF
M17b9j6wGHrvh266CTaursXREGmE2gkWAIjqcjjWxn9ZbFHiDFgAg7EXrJHhetJB
kgAsect9M+MpKD2Uc4o+vDNO9JaJjoZ9RYaw3mX4MsyXTHb8aBOWGwgkmf2CWD+9
0pEfzScWlFB7MFRCvWY9LBHUPNva5dWXdncmKYEBhL6J2IcF6CV1+F0zvc6Qmy4C
o25AEymnKFQ8pjcwqTDlEGCrBLLNmHlhFmk9lwLxXg22v3XMl8uiwkNEalq/TNRe
84/uN+dmWfoBSe/D2DipdwuxK1c0cLVt8OXle7DPA5TF1Zgf/4E8mmeSBW20Ko4O
Sez24wsKBjvaQPCd+8Qlh6DV2kj9pbgrSsKEyQ3ITf0FcUQzuL20dGliWTMdmTIj
YC9x5DouSCYYBK9KR6y5K9h7sXjkWREq45c9y3a+0Qsw/8LL4eqaKpaGfGJOI/sz
ERtRsS2mhl60RtheK5OBqcrX6DvelhY9UkMzHf2AhDN4oD+V7ms/lMmp+p6FhSts
7qkab+HDoq2sLIX0fnWmZoc2VtYE1JkWXnkYpiKu+vEBuTACyi/tYFj0c92R8Z9l
vCZ2Z3Z/gWf0Tx/9Km12oVvt2k6DuB8SMOhGjCIqiZjWviwiu2lO7VTD/X7aFUWS
EnZ0YUA0xQVhBhG9hb1ScHDAkhxy7CyQm6aToRkYE05BIVyja8Vxu9OHdhrgVzB/
9uUFmAAm5Db14dAD5XFTycy2gJJLxj0l+AHqZpVSKLls3I7vW5bNt1nkPWBLMVcb
3p4YUlHtapHcUoF1f4cR5SBU83tPY8krwHtQ9M9jgu7iXFTUds5W8+CIKvmqZDWP
Bg/rDD1KXwmOU6wfmjUraep+egYvZhJFxkMzto05SMOOULapEZMTUiB7Z6pDz7sv
CXJ+iso+P8Q7/HitguALS/HwS71P5fhCFDrqFV7hbDlhbEVGkY4eKh7YtR6Eb4tq
rI1SOA3Iv6oJM8Ag8YvVAovVq5ngQwvjuIi589TvyUOAvvaqT9nIRHGKwBTpAXwb
4r+hpWOYzum1CjJvZ8vpitmy4CLzuEsGtkXaZxWdBz8O/lqXAoiuI7SPGvN7YO0h
SGBLiStDFKSYPba6tZfG+EUe5GrURzM0oOlWe7t7G73lPwUtt3m46e/pEJHajd3E
1/VA5jmhTtTwx6tU3xo6UIgmAvyXHftOouPjEUawiqFDNkmputW64/fb9l6Njmw1
BRa9nqG2SoHxtaaRR+lX36XW5Zt4KS/eJMUa6p3AdGb8zVpzIgJKc7g24hklk2Jl
ccxNMYKyu/mCd9UcP2jAKQm8V09onO54tGW9AE1JYVcrakHp5K+lJkWnG4N+HmJr
5NSLkl7AMW9yim+CMkLze6KdHYuKnF23IqFdpvklV28ebw/7vh15X0jKTp/+/S3b
ie3/0TsOnY2o1EmzUatzwrJCLu4CQszZmt+4JplDqk8BD48sxeITJ4yNbZ/hglIf
YYO3jenz9s6ycAaH+QyW/0575fhLudROWFOr62GmygPsey0Uyv8lmA+egbXz7vSc
b6ecF/OthtPep3mrMgYSnq81sDZcBSXRXy7KkT/CxH0SUKCznPGcANPrkFRfachb
wILVNUPJm4elTOlsDaMXTy2+Af5Wp8XT+s6okvhozAJwHW6xnpIwq+YigqstB7cQ
Bte6fDbTlSIaMYzj9epe7d148chGBtHb3rxYcB8s1owhvBSIGPGamhfs00iYSW6P
VD8bmOjwel4gVuOszQh9VmoWrzuMok8YC9U97IRZBu64NsYlQpv36B7t05hwfhTH
drIcMlYFf8eaz3XwjRRyZRtDuBnKX0mKXOrFXdOvqlUMv3zNyE+nlQVppa8TB3rK
4rE6yOyY+UWJcaJ4k3vCOIZ6sMhcrS5hZjshWQFoJobEIaJxMbz62jMXuR19/spK
aH1C2MRdB3PYKvpLgXLCDiW7RR4YbmX6dj18DV9izh7zvsDfB0ywGpLJTztF39f+
Txt5DpL6wgB872WKwlOy/NNe3rWMWLgcOGXpUT9uztHBXMVV73GLnJ0f2O3MWvKQ
A3/gyl44cFwhw+Raz3n5N6q87bVnUqJrv7cVbFLmzUXlv4P9MjdPzCPpfNwwig3X
Vz088PPmXIq/Ox86YXlPCTIAyDEQK8TjL2CeeQb5JHKTV7PT+ECs00zeyPa5vspG
wHR1YoVMyz9vD8w5GsS8ib/a/pOE84mELlG/QX5g74HPfdUGRWT+7TqQpya3pAeO
dKQ33KGmgIxeBIGl6yOXB5VeKFolwjSuyzZ5prA7zKXRG4vuCEOoyq+s66KqSsKh
bg5bDOeE+cHPbTRrwf/KOnLD36J48srLOOl7TDU4bepWEv7QFU6hILqG4smSzvnn
+LxY/qIMf6qXx8mu0qw6PwRTNncKY1fVlciwtZFZ+hYyvAbUt6vBY2MefE6f3iG7
Rjseh7bz/kyzLxImh/12+79S1IAVqKGkyog+iOUKtBNsbor0QzmetQkui/9RZYJ0
csP60Vszxx314S9VQwXn8hWV+BT8cCC3pi5N5A3MC+Njn5iR2leV86S5B4W1jmxn
J5WeqoxHGsshQ6viu09N+eoSWBhDEKf1pREA1zuFlK4ys6sMJHwjYOOBN2HLUM59
GZKnZKcxm6wg5jXbnRKQwT/y01Fz3dIV0L0samfOVamsnxgSjIWNCnzalrKgQNoz
Hg4saBeSPUVjDj47EXnufVnaaAfn46QwksZHldS9W+RWPgjkzcYPEQZZwViJeD6O
+MYQ1KNkDh5grmQ1jJS27ijAZQsC3BZ40kTCT1Z72AvhSkYGLZ4X1fefyITxO7Gx
vAwuGLEv/THerS9SLA2FlM6FRk9sNISGZ3OM7onZiolYy9pBBmtTcYSe/mEsUzkQ
hEaK9AHwpNXbsGWs8kY/+Zo6JzxsoRVDLgqdHatcZdyA14Nipge/x+JbpEaS0Q+o
OLJbJIwKffm6BWmtpfnC0Hnjsn9+UHbuhAKSffL0T2g0tG/GPGGmOQdO7zchjyxF
fHgBhSV9veMCEESw64JxN/lSAKXFoLcO5HuFaa3JPOUsWnG4URWVgcSY6ZuS7c0J
N/bsOL9mRb6da6/mlUi1cJVGJ+UNSpZC+PJDujJ4n4izB3631JVDCkaaMzD8i9T1
E/g9IyjlhIvvNLephk0Y7xpuTDkWuwibHotmKkwtX2+MBqpFWGVarP+m6djdoDKQ
d4J5/9C+Wl527WkKqXxRwG6BYtZh8teM0je+zDBDp/kSykehjvIfQo9IGkpbMRHm
ZU7LGubaEqupX0pGDDLtFbt2KlH/TtdapOvurN1nVEuA94hH8AIBA1NhbtACU0lt
rFD8sB/Bp/FhCNhK4qKlqAOjLsvToBe1GoNnFcyVmrOwE071krv1uGg33LsRvDCz
cEKdjrld4MHADObrmIVg2XdpbIZgdsQQnYIg2Zr3fOK22cIPWtA4jFchwm1WHUhT
HbWnXtXTWetu0B1s0PQcBztMh4kr7RbJ0GinCmeb9P6wHYIMovuSU1Woxu0x/L/2
a8Mfp4W8ykIvW3TxFwzyMXMAjyMvNNzjvyOUHv86hId+J4hAJsKsNTGJTvU4hDX5
93VBL9+m0vb68PoygqodkFWiOqfjoXocRt9lVQ4RTAoXx3445AsvFNdBY6ieuo35
7KIOtEOBDjpptTgodEgW4+2yNe6ITPOi66VDRRRy/Dgy+k+i+eS9DeC3LeHOS+ch
IQT7eXaOncwD18jcEsP4rqVQPcxJv5NhKDn1VhOWuaBuVITDjn0UJS2KLzVwAzxy
/kE/NzJ3NxWBmepqhr0Y5YX5HYfBywyVcr9pKusUoWg0DSQd59Xk8TehMR+4kDUd
fzbEBZHCDf6185W9HkTiv4/CHVslXGr5OW6D4DfSPA2YOkrAYS9ek5UqPUYUVQEn
6/0axxol+YH2pSWYUGS0mBWeCn0LAN7SDFD0LT2w3chBKBipw58D9U3/9sIka+2A
F/WngaSWhS0S8kUdPUF+lvPDwkD/lxM9pVaD5dyTWNm7Pui2Z+dnPfE5QHKTnQsr
lAJc3Y+mai3MpnCUCWG2QmyIiA9sNjnPmE1KlCQbL+v8GNV+2xjNpBMt8xlieE2u
UmUpWPXfImv9mTY+/DE4a2sztPuscoBXTynUEKxup8Wixd8CI0lL4ORukIz8iyUy
aOmuItVv4SCByQkrwAi8wzDHDcUbJsdCXXFJ9q8skp5Oc2biu8auyeDcF4M56L+X
Sw+XOdV7kf/0feAQCdqzi80w6XnsSYszHb7i/Lsmic1c1r4ZzOs7M0JBcofLZneH
b/IOSB1mWxvSj9EXJ/DzWJjxOvbHgSYkiHecv1gRjkVGyrtozF2JcteOmHQF+t3Y
eGQ2rT0Kz7xof26gFDvR9Ub4hPSqoTfSwrCPlvjheN9qJL3npT2YQD3xUpIFIzLR
LASrXGUAzteOoOkK+ASRRA8wMWAXmiY7Id6a8jSPhr8CxRpGY+DemkNxJDwi34r6
m12LXbP1kI7nT+ScpGU+0ITBcYVUXiXn4+h9xWuufrPAg5aHGnf5yYgOwwiXfBzv
PFnWN2OgXZ97/okAX3D2EftMEUIscWjV+aEhSpqrr5iROGh9FUjRol9CjMS9zSGm
8DDSKKa6gVkxHafwcWkHhcxV4Pd6OfPZ6aNvNfNfUgt03jhcb0jiCz2iGp7YGUmU
ZaF3vwvK7I2/JYYbWYLG/Q3SLIzuAJnLn8EVwABCjPiRYEGSBl8G5Rr5bjAmnFw6
+Ct5YR9+dFZih+AjqjSRQuIqPNwHLYxS3Jlnl043nz1IOcbpW7cMQr5w+gmo0gAV
N+uWo3Uz8QYwajr/vUyEdtSEq6vS7hDP6w6RnJQavff6wY1UOyMl6LA+QsGZtPxG
C2II/TNwbkZ/yQwAV9S8wlC5BYu1ez22FfWUawZSN+0IXTg0tCWGE56tHfj2xyNq
AXxnWVdPMHnJ97Xhul/gcOTpantIk1AvQAs+ymroU6D6sF0EF/6wAwR1uMB4Ndtw
DoLFM7df5b61W3MHP/Fxs1JvZ383kwMaBysCW4ZrOVftwcUSXyQrnr7zYtQod9cG
t87IUSOeovx+17vZRzCM8Sz/aJQ5GMfhqj3zCIkJf0pD8bO+aF83S1eZcGwTieAC
HB5sb89oucx69b4Te4zop85qVDJ35acC8S9CqfJnBeMFBpZ5w38CFUvm7aQc8JJv
wQ3bcNQQVeEGCSzmLwYFSUw8baHDRDEABy+Fi/czNgU2CgIPuQAr+5YgrYxvRbjH
7JNH14hxFCN4WpShd4d09+sIHWpa9aVwb2EWd8081OiUnfHbdYaVxBCLzwLnHZic
cT/viX7OZ3T+wSboz5hgq1gmmtA/mLfROP+YBzKrnha9WvFadi2mM4+SNRZFccYT
vcp244kBdps3pNZ8yagHoNLyJwCu8V3985sDnALlHXE7Cu8pptCDtIk8TIz9ao5O
nr4Xm5vokJiDu3U08kBLk/UgL1o5i3v+Wm+hkbTaPDzrbJv8zgbw6h9NGVD4S59f
5Am0Qq8P85BuqGw1cvjty8PS5xOGFXrxnPjCONK2LFSdCEhfuKwog5P0adGFcq6H
dQMJD7Zp5+SjhsrPHgd5GzNZMySk3BBp5DtZFOP+bc8yKkgQMo2GkuTSQl71sdmQ
+F1wJBdweyAeYkrk54oFCDSdkOPzoL4Dl9BaqJGtz9jVnIRQbGkRz81NiS9rp8Kn
dbj+QvGzmeedvJX5B8Bkst9ZrPmTBqnCXgyN+wvuA6uTYtf4bYmyMFWHzE/0rUow
GBvcj7xPbnOzn7VwyT7XSFxwdyOO59oMHoFiqUlamWEabQZG7K++WUnfCXH4DYSI
p3TaO3jRL2LV3LnNhXIrFXRlJ2q0J6pmzITj4xzm2LNvS49xxXcxzEmnT0Ano8+7
x1qQWtWKAx2DHcRGqxxe52E9sV//b8lsFPo8VHoUFtogJpRBK1NdvGTApcog44W9
uG98JEzY84caOxUVWaUcIT4d1pv51LWb+K5rpIIUovjhuGF3S13wff8qQeslN75g
/U/MVtdZmsOyYn0AA0H53hLHgoZHUNo3Q/hZNlYFoqsAhbZVpT7WGE6MB52gocNk
6GBPdY5qbK6Ss8C6dkyKkAcAsqVnUg8O4b7TvagrnNLoW/ZMMf8JHC23ph+ejcqK
memgZfk9RdDQ5be53PSiYycH/G2ShFEcE/a6EVYahr6IUJzbQDXD8fkQlWWroQDq
S//nOMxRLSop2uCZRfBuslpTXL6jToJ+mG/MvRF2fA6OCHho7xDSfqeYyuQzaBqJ
MyyB7vbtYoqsexn0F6Z6WVun1BRzuGP3FDrTagaMNyjrLcRsIS/IAES9irOy2o5O
fSqgEt+zvDPbQLuJZEmK5zDnIvgngBQ/re2MEUHpcPaXM1d7jQPIXKR9EYYO9LXN
qjXklCxlL6AegO65mAxUiJUFAH6J7Vpaww63oLEwl6SNgvk+er5WrjcSkUmnXCKA
3XxpJ/+IW68F3Fx5U7CNV5bFEKSa0Sz67SVkLb3SxIDWI3fVUwgnXuOcIsC1lHQo
TMuwzYyZF7n2H5fc4eml9K5IZpa3xwaKts4vvuuSsK6subzG9f2i2Nokvv8/HPlL
4UoJXcNmOTPh5JdvI/oiB4ZZslhT/cACGzBJi6VXIrRlJsr4S4mR0vnJm2eZqN9V
XqXfutwBoUXpi2WBbzewfqCsxpZApJ4KnnKwHlSGMoSxTkGt4+5oRJcolhrshv4c
b1SYL3QnK7u+YQF1KslRfRdS9QlQKbSE04T5/DnurWGn0onUJaM7gKlRK1Ekb87x
BJsIf+sWneQU1CeExbB2qtPicceXDXFIR97IKeR204uRkFftqC/7TXDaFe2kUKy8
DmxQhjZs7upm8D8y6sHYQ7sTEO+rVdwF/oam27S24jYZd3w2sGRG3ZcMNrxBGEsm
sJyAHDXGJKS4YYCio3HYzsf2PzFBHoTqJX2z7TOjOZ7VGWRPm79Z54XXSjsY1JYq
Pn40rAiQkDE0iOK6YB8uLBTVERtpM25IAE1BcQbaWa/22XVHaUOwKUSIzB7iim6W
jrujURiMZ7Zzr5oDTp2QkBCXVB1Uczjts/PJGYR17k9RASV+E9iVchWMSPWAPmnA
lYCeBLoDymHoaA7kY/S3hrjjwNJpWmi+03tc1WQLBLX1xNGMFI5LJl1QmL+CI5lK
B189uiCDlxBq3Mp09Uv8VQwBzorKklCiJpOF7KcZslrrq194XHJ5lHGawt7BN7h7
Y0MMKosZz3RIJ2PbrhYTKU+zmfBU9BhOQRNSNQr9k1jxiBnvQQDGio9Gl8jqNBDc
HbdAQsTQ1CvxvcCiP5lYvY4tzd6WPN8U231+0zhqqkayUqBuTzmQ3gIhQJmuc7Tj
9J82B4/GqBoflwoFfr8G5qOKEaLvAnDA4iV69mlagKuueggVH9ka0bHIB97bhbwn
Ryo4aqMrTKnCoMQH1CSrY012EnYAUz6evgXFnt6OT+OxfIfBc7QBSW8IV91ksFmA
5JFk/zrobHpMUr3olRzjOlJDWbbEfD0ft2rJlqGRbCp8MUfsVP4B9/VPVbH/ozZa
aXDj2BV91ARlQBlMriVTckngvF8MQ1gauXtB2khbC6WssWnp/J34THJUGxq1CLfv
s7IjbctlxVTdD70yL5xXRgGRSbxRdj9A+z/hQ4B/nlPi7UpaLZn4nd8VwMUojoDV
/VqjN7S8Cga9mG0Y2/W5OUbAZl38K7TRZ9LHCFWUlF+RIXm8oAT0R6rBsAWpHhgk
AaU9PfZEo8rmxnG3znznKRrmgfWsqzo0rg7zdzwTJCvm7jjhsH5cQHU/rlUPWVNQ
71KiW9Msr8oJCzQHxOlVfnYfvjqJmReTIAYKzqrY+9345aZmuDYPkB4D+thn8Lx5
UvU9jSPt4/eRs8ihQbfxwNzAT4VbaFwjpqc4v0oOox9XO0BdJl5ro/kvsAhWdAsH
AkVt5obO5czpBLR6pK+CYeAc1GvoM4EuatMwH9FFoEBbaR89eDVCCG2cPApYFH5E
Jv+GBR+xnoW6ezCFYAPddaqx5B1mm7WvKQH4ny4egkFFWW8yupHFs1IXaNptJFVE
kw4BTkGA34BGczg2rv0yhUGscV4cfkCwBTvcf4uv1jZyJvOParCuwaIjRbfD5HlX
WBE0NU0h4RaREytRPCJwiXVHHaQGo8E2fGKMsa605IDWMZZ0DuNi0U4L+yoOlYTN
qDkvLmsrsWDTvJnDE5OLYgxzDkGYrs+gpcTuP9WOrt8+NxtZCHZNTuqqqVasAEU1
b/zS9/4AV07WndbpicRqZPf9jM0/QoEho87JlJ+resKaEeotf7be8eeyXTXx15nF
6ABayaYmYb0Kh9vCL3anzLWGYVdIbHvkcmmEEvH0q2A3Yd1as5+kh2J63A6C7BVj
BV5Oj/39cIm2RdS84aDq7Yg/b8S7eoYXrS2f9prEHFMXuEHwpU9WiuSGhliLDmYh
gMxwZhDca3er+ZcxO0yqKTY5WWiwHYGXsswrF9fqooB8JApHJGTsE1Y4Pb3lWKFe
qRpEWIFlsv6wi7uEWMtOVkqAEz/8kMAJ5NkTcaPl4xqbLbk0airVWtD8QBhZdaoR
1uIRkzrnIoJITSjF5+a95pjIcyyDc5jV1yeLAh/Rv/UKA+Lg/eMrItF5RD24Kx+K
U1doJx1KEHG35XM6+lk3frByS9E/aT8lSU8V9722Nz7wNK4S9236rztRm9Froqdh
125h3Qe+FrK6SvSHT7lAv5Q0/i6qJMD5pWfcrJrh22eEMntMI+p0bmaIZo84eMlv
5qyy19NiRMmvzhYwJ8ed/BQvxmAu1kvmvvlVrzjWnYFXorIBZwRyr19Xc4K9Bj+P
mwhATQJu79uEAFTaAcy2GxzFeOHyDNieY7Nf5iVtZzG/3Joxbq03PNbi9yiV6zhV
tohBtiIhkbCin02pfz8w8a5prHzgIOFOeuYK3zNWaPgWQiIGO52iug4d0tpdMNUV
kSTHKmmwoIc495j0f3cwxc1Jo5P+No1sd5rRMcwajAgNpnDY4S7h/cB6Slj0RHkD
U0Xt8Uyw0p+dKBsE5I8Vy9P+95I6pvb5fSy7ckoI9F8E9/+rOUWamiUSj8iMvmKN
0IR+824EPF/uz9KHjT/bZbJ8ptWqRlhVBcWWZdx8IfsS2rIRMEFQAGOissVVf+X0
mV/ZQyLm0pdmq8SBvZNQjA4RLiBDCDchU7HflpVG6ONM3uilJIsBaeiNUaVv2Cg9
dvDDXkQxTTnWk8nME+ldOmme0gWcXZ709dq2o3WWbzQ1b+DnIc1+bG4Yyl2Amc++
XBUbKEuJcVMyQB+PUzgFFGdi8t8GudsymuydEj2hPW285ZQAeFlUydfbBw4qa2H9
YhftnfmBV+7AE6MawITUJ+izALsveXoMXqzY9h+VUvpPDRFQq0HuDfQOQ0tmxu+x
MH8RVN1BtGf358La9yUNVvU4eYhyGpACFebfCFbgT09rklhepGxuliIZH5DmBtOM
shXeMXVMwvJEBtdUBVizkka7+8DIPDByOkBL3WoMZXBVep15DMhtbtjfzoiRzHIy
h/xtDyAb8X/8st99aiOhn51pc7KJABTin8400HPOEwBBLZhPfLTXnVnVlH9DnMSc
1o+HGhXX3imUa3SauCcobYTW8CjKcwSVjT1G/tjmCroow+Xu0whYmlzK2LQEzQlX
K2FqyBrhaNrF1KADrkOqUBcJ3SGhb1ej7YDVfKL0fp6U4xcKModfnQWkk+uL/obl
cbzwQbrvLmmh5qD/nwDWZVcL7xIxdsDDZdFW2sRucf274Egpit/+UC+njJ6TQM2P
Gks+2IyJf0qE0j6LcptsJrnqYL+e/pycd3SFT1F50Mrsno+U+PRlJUOOBWZHOTOU
O6TqJrufYnEMtmTbVlIUKuIk4h7vwSSNdveC9rpFqbLJ/wqR4CLvT5XnyVB2e159
GZnBGCRfSWK0dkh/VNzIbhieIpiOtce72pT2YOOggWZmo9NkNniXd2oSSFLeEPhu
xAEK2IsfrOjqYFm7/D9GveM/WFaocw0udLTb7DXhJLpZdn9bL+bEDBEFW+WDLTLe
6EIySXWxSDF1avm1Reh1EhARK64+ACklP1+AXEGKpuDzkmYCnqucoqEMV+q5qYD/
GG1dXiYoeLYag8y3PeasFUTHgX/Hp/q/TAV8KYPdHx799WaUVrNoVo+mPiD69ahj
StV09mrshVJp6pD2cE0hwBwyBocXpy9cF+nKyvX+zaAxzwlxkf3g37bcKPMhTAa0
DaExKJSuXFzok21xka5ppNySPuMzt00lD9AgXYj99La6ZAbtc++DnWOBmCZZfBqK
S0XlPIlNKz9cqA6MTD6kPs3D6hvqpR1Ed8VJ6DtCAUUblVn9yXhbVb9wFN9RHN/1
RBhgaVPNBArzSiuXJWCfPp7chE88iRnY+sed/4FjAfQ1i1EA7s7vnsnXMLvBeyGS
6OAWVbVRo7JnY80qwY/5LUSKhr9+9Wz7vGAIitAhrdts5sRPu4PlnOKJAniKHKsr
CaKJLPV+nN9IjyiKx4fgkt7y4LA2k8Un5ZQ39n3Mzdujj2N0K4UJ9ZSjJ2yaqBFh
rBdQ7coL++63Q4T2BTxKDB+RIXIAA2ardgm0LUAZaJbja8bT+X7zMgWbxGYPSJXT
55hcrIhnSObk8+kn9j3RnsBSginBASFxPoM5wJhP63L/X+l8cdWxTCT/490MOgTt
NiEZUYbJj+W+WppMMfxj6hjioEEWKmImV6cf7gruGaRRMj8p5cj80vQc89A18zdN
E5l6U3M/spzFa/R+9ld5SNdS1ET3n/XkWxkD4q5dvEDYtRMf1U5f4nIBU5gRkFgy
bI8apyCY1l7ybGaxWz2t/wCqR7K8PXXehYtXD+G2iCXepS4OwSM5mDJ2V77gNtlZ
`protect END_PROTECTED
