`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tQ60cJ1waFOjrs3asemwA0fnuVFtGkId2SodUfs3UG5niI8jAbkzw7QK2SamD4TS
pAqYxGcQbKLO8217Lwek/MA24shj9Z7nxn/mbPmo0fv0y9r/lvTf1rLLCZnIMp+y
juig2eIJzzQPwz1uICH474/DyHbqRtqP22S3t1C66Pm2M1bXv8sc30DyXlmxXc82
p1m+BhLlmhjSa50biKSFXYKmXfdD/6tbH7Il2XrNtxwrayT5CWLV3Add8Tinopq+
w3gQ1Hi7JJz6n4vwhHgZ7gH7ch1pTT1pUrurmZUUqiwsxnZTJaDwt23/hCp+nwAl
j70paCN0oy8n2J4tbwItEP2zeJ3O0HqPYkBX/EC2iNpW7eLH/ISzP2uWbMmUh3uR
WGvc91w5kJGENB3zSC23CxXLe1lNa9pePeo/lKw61fUdt73qO4P9hBbiKX6uJOHW
+Ts+2/j4LY+8kKaatxZMlbeZ8Y4Ppz1/d9R+XRBZoBI9A/FimYx0Y0s0DFN3OJKZ
8PztAn4v1XX+fVCcG2XU6957L5ch5oD0Ew6ty0Rbi5kN371elRUec3H9eGSoRwmF
/zoGxfYp8NIKYGLTCyDttlaxZRSkMmkf9mYtTtfGFL3KG+A8LVAQzLA/ZqtOB1Hu
66bQxSQJ5d8bf6eDU26EiJsg4OnruS5BHMNobYKYPULJ9Si97/aduDMwabbLSXoJ
dPz8B3nzYbF/hj8V0IjXOWzw0YDhSpWGL+CLtWa7Cgb/ioIcobL56xJldHAUDY0C
RG2PjODRho8eAlZQuOh6D9kIpHnagFW3OO8QA8kYkU0D2RrZzlZg5G/0seBL+Y9M
Dd0yft7E5BuywQ7lD1X622X5/u66OtHfKe/4HAdkVSP5TdeBlDEFrKS8jm0Cm1n6
Xv5OJb3t7Z6hrvChJbjpXztChy+pm7975AjwfGkieUdcUqlfenikRnLIFZfGKv1V
0qsyG5NmjRK0wwoagOOoWb5ugqPNp7vEtx/2wFNxdXqDSzFTy1juyOsTO/uIh5wy
1vYLKgdmdlPLsgb0wClmU7Nv6LhMuKfqTya00D57cxPlSgok/UasoCF0DDdKwFuM
vDYSqzfCFqwqz44GcOHDoOKeftdtSWwlJR/Zuq4mqamlXRPx5r+kFxm30OezDXRy
vBwLqEaqBZyJjYbvEHesn8XnROAcaNiDPerfbdGNAFsAtrcygezuqQ43tywIVi4O
rfHjv7Ve1UC6WDrLMELwTSWVebcWtkpEk4nnoQm1AnBYnJ1eDUIbSltqqQZLB6cA
pnVxY7FRxG47WoDOb+bJZhvrh/3ivdk7yOqKHCkvc13Z91fPaTuMADFfh6d4qkwU
XgqreucU3yk+1kaSTRWeO81GJWeEYup4HS9I5gSkxZtW/KFu6k6RLOxuj8sJhgHE
yx7EPyv99gQKtkfNvxhVmpMRZGV+H78iwUsCMNwSeeVTWLCBaXSJAxOtvKsZ05fc
UA8MSIRRHULx1sRhnNYi2gepyqiD6Fle1q3YY8E4ItQ/lYn8aWKsSMZAvVveww5O
X4tJfboZqjy6GsNpNfVZQHrIDhjYwiPq2a9hwVnLITbp5gHgB7mrO8sY6gkRO/qw
UQTi60G1nvpDmsh/YPifpbWY/O4PaXO2Q7/QYLfYvH+MEa2UD1Sqb83lhiNCNwIp
//pNSCDKIsLAcgfbaHjeSPLIj7bL8V8gaVZas+k/llPK5HgmvjB3AchwZZ8m8CFZ
twnSIjecZhwAHSnBEO4mRAl88hFEpKnm1fCEd2tSCqjAdRVtjdrK0ipv3EzVIv6J
+BpT8wMj5DiFJiBCb5Rte423fW4uWKb8d4Iu78vD++G+mUKY0OF2LhgUbg3TTCJY
XHQIdXkjxs83FTjz0/eGl0AAZj4ExQBeUsAk/IqI57HRlCHRx5hQHy5+/V+XjWVA
gRjbeckwXdC8DzByQd44FqEZeDpUFlAFPwcTGAE97bypTzRjEcmrendWieummJHc
Id2nikU12DgmwI3ZKYUyBHV1LHqkSSxqcfZi2/iY0nZh8zS7QLNX2D5iEgVKhA/7
KyPa3q8j0uooqCpPTYlRZxiRbX+my9/6QWO9kW+46klPgf6xF7gYE7L2OGUlE+FG
40nBNQxKuEp/4faYpDMq0qdxW5qJ9rDxWLW7vA4FsuEu7BrWLjAAnbkrqXPHroUa
vqvZe4trpuXBT/EtwIToGNt4ot3veVgnnObpyxnj9Wk4Ehh9PUY0jkqlT+5Qbg8D
389CTVRGLfo3ZsPiMogUX8kHcXQzqjzV91E97zt5skFMcZHJZzcDjaLs+uCmDXOJ
Hvt+ZaGEnGEdEwsA/GPq8zXXd14wQ/5SVOxuKFAXoQf14Lnq9AwitFPh0FZwX4AI
eDEm19/b+a4ztvNnOtntQZHVWRVY24J7yd/xblfYmvT3m9zGwUlTkUnlU2TKTykE
6fEHD8vxmbkMLYhn+eUONn4bhQ49WSut49VXpNS7Rx4fDBJxW/WB6oxo7tiFcbPj
ttDIDj7HEiJVX8YpxPJaWUR19pfJQCKZ4GBOJvK2GRv4AfvL5oycy4GsMrNJQgca
KpoO9nh+JEivmF9k7a1o7rT+joX4TKxIRmikUza6dIqfOgWeYmxFA+F5E6pJQWsZ
H5cAj0x8mGvHD+ec3FXS7pGSeURFcu7AUmdnIM42Ykm3r0podEMtDpgwm+Hg/5PF
Gt+fPJ8uxcBDNwpeqy5YJkQXfvWH9/vQLezh76cJ3d4qvlYmqhAfStyD9ZT94kwp
Nw+YsS5GMjfGyCmo36BdGnra1er9HdqStMJUOp8fKSE0Bo+OWKpDCh5khT68YzJg
kxnGTxzUFFe6ud1R7FdYfmwBdhfZu/27BneG0ZZS8cBpOESBphgl2ewkqbfHo1Q6
RHX+CIiDaJJ4XBopOckcNDgEMGx+OpkH+yPCHAe4UNh9ULGCAXHQJCHVLMIr1WT2
wGiFIhp9RLg6sLpeZLukE++fdck/Y5igEtm6BfHMRsdv1OcLWGCHfeiz7Oyv1tQE
2Rk4HJ7pPJj8o2Nt31Suv+6cz59oP9N0tHNrInAHpkAM757kmagi3NpI7MnLE3g/
076CAedTGrk/IkChASFaTTAxSHFJ9KEAvc0ZndxIw/ZgTdLkU88bsC5z4mReXjFn
lDwMp5SvNUs7m4MoMalsaFZ+2WBHHcGXTp3eMU2et/zIqugQd7XF/Z380Tje18Da
spG7aF7ILFCbn8E7jNH2TNa3aMfCGrOnl76m2T5HTNI8mXaxtbu2Wcm1na7MfPdW
XUj8g538WGMwTvQgG2aGk6yJW/4nToBUmaXJEHPjwftwtjTe5ioh3pAuKzI27P/I
3SUvkAWRLH8Q0BBNz3FQhWnElm6O3iBejgIoS7XAn/DXmXbYrHuLzGoGuN3+BNrM
t6vZ+c3ORm8fvl6GePCtkXUEThauuQmtmUBWZ3E1ZHXAGIxp9NDNUa7KJR2HgwJ3
DD3jsEN2AGAOpdVWj+Leu0emptEq46prvqXlqMxfdxGbB/BbJhePpJLanksnSJdI
+TDZ9kzUZXbyM6oiJ/9GN8qZG3u/ppJg7jMhFdUzlRz5jqxIHTe428Ojfnkw/1u8
T1pWjUmBLnsUlhpQLHNovWQeOWAEGwwKl+rUhNr/fhypVzV/fg8mMmTTf1gWOl2L
s3rtR0AedOeiFe0yi4C+cUwGoZojUGS9Hzhs2qbOGktPRd3KsIXEi5tUYk4i/6Ow
2BYgs3s04bDMQ2iu007kLyIXhVSTZUjClhSTtvj0P+NJRqsYnJCZu5Et5uomR0Z2
Evcp5SLi/yatgWBxqAkIVEkj4zb3hmqq5pKxDRSV0kh2iu6mLlOz/rq0KE4d7iWA
H46RmcMCJgBI90enid1BfXtKiHNMkyIUZ/4eFCI1acTrrLwC+3CMRQZJVENxQezJ
0zuGSQvSi00sifIdNpiM9n4M6cU1oMCRgR3Ef/3qe+Gg7+HGOeVpzouxOps0h9N2
tVcMSMp+/nIt4+boJhkQFayreiM3mDvThPUjdPiCPBIw0lG77gYTnUA6FUheD4/K
5oKUYtnYJFy+50hwXeo8hkw4fun83OaDnlGoTh5PKKobLaJrj8qjWpA60I5ofYQM
UGtyWsrsuPU7mlvikljFElHB1Ik20Yh1sCbd0eAYg6UnrXxLgZporal+LUWwlBJt
su6tWuiOz5n+vLZBwu29XePH2wkIyCO+jO4KU5z03NScDf8OvVscmxEpdemx5o9p
6i3djc8fPyekhiIRC12ty3c88F19etCxfuom2eGdPEfPZW9Qo8jU3KDMQAM9kSGt
OsqHR+cs9yOUm+4FhirMJgcYXK3Ulv73fnZ/A7lm953VzcffVNuZNpnRabYXlDiy
1TfBBq0sL4D9Qd0doOchFtpHE32qk1GJ53iaoUW4a7UQhnfnE5gOH8pj9vYIrqjd
OtMQdoYHRl5PFI0Inh+0thRrap8VmR78zacIV7hJFy+QkTf9+FvWgI+QnXsIuA/+
kijTJLUVMIM8c1A6Lqbnor+E5WpSsS5E+amAJOoxlTprNerQ+4rIiQX9f+ALTtlJ
J27ievQjVTrWERbpB1V19hZrRjVbIgteIan9Fn7wUr62FPj/aDasmmmhp9nSQ+Ww
BoAtBTRhBkrrQP+cXdohHyFT/gKVeaxsang4R0VNoN7dm2W2mqTmN0lWhilUi231
1jzZ6z0lv1zgTplD09/YmEh3HVocLN+gVIBVjha+n+K2+/GtO36KrP2MVMeon7wb
1xQkIHiTOXAbyPiVd2WDuiWgGgdAOPs2sM3kY+58SjGl9hZ5zIYz3tn0W7nxu4aX
SIeOd3B8VkkknqhEYVNjRqXHbHuO8sL0ElTC3RKor2dNd+abY2T1HraaCI8zu5LI
iM7jZoEO9/WGtUzMOsWioTvhlVMS+f6B7wmhHF6lA45Tv2tyFvA4AzgVds7D65Fa
z/BWGxjKfPe1j056h6z7fHxb5HmseD8Sy0sMoheu3HN1hcTokg9xsOhHYfEnarLh
igCdKrazQPrePR9rHpQyCi+DfRzKo4I6Sex7xKUUAHkpwYOgLIX/nsjPHc/dvStL
Ij1CRwn4zup+2R3ZtulFGzC/uyMy2nrTK9tG52WO49SS5dOdFGp6W4WX5nvsURSX
DBTGmhB7lxEb7s98Bl6Z0DRRgtnBvXCM49Uv630gMxA3CuC8PtJ8q/sphbbd9hgN
3GkYj6aad2FF2RrEiAYQHCBVYrI9fDLKrtaYHoKzecdJgY4totuzC6SUOjGBkWmw
ZCMIszPt+d2DLSiDXAib8BeJXl/UO3yogmRprp/TR3S1k9VSlM/M/jKVgqtmQTFO
g51rxyKUZmwAy4Qn83X5GISXONZ2FRbV926duX8ntzMNXqYXigWa19SD+xcB4BP0
jETWsQj1XWbifCExz5xl9jM2nNHxaMGbFH4S2ccxpqYMkJojwdryVCzw2tKE80ch
T/n9S+T4lZpN8O/Z3x5DndZCmvVifUUl8DJvj2ysslRBjm1WowLiU7IVF1+3M269
ztRVwyknFWXL5Zps1SZ4Ok4eEB81qzPnuJBzVk1so7ql9tc5qeZb9k1Ce9BBieY9
a273GQtoCZp0qVq8yP2kXHEEfnQjwVRODFldtpDJJqSPo1PdiPsC1LKH5q7aL/Yj
CKLgwPWl8C24wWHCphb48NOt2YvfurG217ElFSEqDokvj2gVcs8LBpsGHXqgnhNf
G8QmODchPVuoMMQq7EEHUJaO/u6ZcOvAkxnH/KWwdaL/BtDtS0r9juHkc8mVFaxU
htzWNgh7eefJT6FtMrNdcUh9YaBN0SQAJzEE07kfUA8j7c5rLcUcauJLKoQa0Ja5
Z7SDJE2k5DeHROpBb4FJDv9WiHheGECM/+aDmMXeXnJci1hqotmSUmCRCUsZ2Ext
Xxxyw+RRveZ2MzF0MDUPAsWd7mdHmBgzQkbJskwSBqzZt1pujBFAhlFU+qKfXXv8
x0TAAorvXlkasUVeG647uKvITAzbPNasjQE3/+pCxqSAERiejC8gW/F+aPeRJxcX
kXTJpuLpRRrQmOnHdI93uadGswRU0RWkuKss2UTVR666P8uCa9uK2Z1aSi4nqNhG
FJysReIRNvaOQhjyd+WqFVZhBjGGeuVwIj4+Y+dRNNDraUvQ77ifc3ZU5uXYISUW
feWzjcYgImk1LOrmgg0eL4xJE78YvANycxsMc+E3fUiy+8VzL3yQcQeNhboGzozD
Fv4eEljn2b9Gd+9+R8rCQlC6OQV3YzntWTBImVa5PaB/ZJmoCy5W63in0KmAvhN3
LBSaCzYZSrr0tTZiYnmujC4DkgZvTEMGdn0fhDzWP0lEF3nUpVvhEIG29hHIR38R
RlY0GqhMOtLOOfejSq/NYz/WrqatuVTqQlCElDIYAxYUGeElA2KTjJ6UBzTuk7po
ljNM6oUoyh3c7KeivQ6GjoZ3linTLvBmwJWkv3y9z8a/5yd1lD03IeKhSIb/jX7m
GMhgEw+G9Ln18GEuRF6Hu94/ZdpDzLo0lq4kLHbwk4XfKhLIEM/TY27DTfD+rh8j
bDcxy2RS7fN3h8wDBfLy2vBqFh9LEPVXpBPfpbg/f6qUqKu8pqIvtXT3fMFB5/9q
52DIbjVS7OU/03Ketz8AkX3HDIiXFtoWYhAa6rB7SuMGNrrSPu5UxxjkOtlDdeoV
S9fIObEmvPN5qQDR5kYWihEDQYpt89j49ww9mxibdN76lAj8jtJadWq4YCIFwQtS
lAj8Gh5VnmH4ONrQebSGFQC0dRiwejFCSRo8VSBWOaRBkaglDk/gxpcIhk67BpaN
R8+RtDXnra4wn1FJpVuitJ2AZ2wa7EZQJGBLclDVbUuxhfHQEtbg9pw3t/1Ait3e
EknG1c6dDCx+t/LEib88j0El+DOtk/vTvCr/msvRSD6z3v6vmyoWaZ4OXVVPKIPX
noCrq+NCUB6BhWfy+X4a5F/YSLNV1QGY8bh+K67zLKtoeJz6Lh9MmfqwFn3bHEuE
RpSxhpGV8zWMZd80XgJ2iV5DT69Fv69Hn7VJETDp8ognOvmaqbgFpORDSzD4CseC
eNI2dQ6jeO4j3m2BhEKe3pvD9I3J04wSv/IkbPhAWpYX8tdCNEr7hFGIE05+YE1c
LOTPgCgwets+KFULC+ZoRS7S3CacQ48Mf59dLQbZWUub4PC1QOzn1/qmfe8P/5PA
G4XxHdM2HQfM5c4fKwFbWHw3DsoazTX6k4XyLlV3JbiKu6ABLQFstSgILel14kIk
OTdVJyJn+kVdp3182t065nATI/CGoFF8M0SJf8/y+4Ee5i19sBEmTdu+0VNSsEyX
jfUljwvD9Vy3lJ6ebMSHkDtdziy8HoGw1T/QOCN/IueTy6hMthjDByTwKQQpXlGI
r6urwDzWniryPsi3P3S2fnQFr7tazExcUt+yRJtPF5Mqin/qJFTTrnlvx0RaD4w+
MemGzG7lhl6GNb0Tz39wTQ8+OE68m2AuIUKgyQZqiK4qwPwPBaK990ufeznmZCzJ
lAa3A3N7Yd0Onp3S0vg7jOrAWD31KQ1n8LVJ34nvogGqSE9b6VAPoCZR6dezqKD8
j+9w4E4N4W+QV3Byn44OeFw/2x+Kwj6CggciJrjmI2OeOmz+UAz47rNPUtNcTicb
xL4SeLGvmQciygU2HLDYCAlQBQrxctXc+LeDh0sl3RDKdy/IzY13s8IRLNwcJAvr
VZBTIdaWTzuoT7wHYPJ5YyV7oIWAZ/lvduhUz3md4pwTZOgW/uiCwzxOwceMldLK
qeG0UlzUM1Qoo+y4u7SMehtqJvMLohUYrQ1A1ajvpKO/+LGrN7ZuaBtKSnk5/tRB
apGik/yMema3l7y9yaHOD0Y0bpR4AX5qnHjMFUfpsfwjIj9pwgGHP29p2J5bVtnc
islYxS/wllIlphMpsszWXBeu/WFIHSbti8gm/AJMaO3/Rq5u6mmTxyXTMvpTo/vb
6VxMo3v34t7Njb17kmO4rZ3DtAG52Hh8/FPMs40jt0ZhNxFN4pkoo1xL7ZhaOhDP
wFM9ojKcdDU7JdtVredPZ8/Z76E+fQgQLuihnv+XFlW1xo+Ah86wIPj5zgBOyUKP
dmdFwP0vmJBvfSMT48MtAE3646gm63pvpDXuT9jeCynU6Pomhf65VmFH5u1GxOIW
vi3xSkzxTCDi9WkQqN74D2xc6LcsvsMV5i2oaH/yWm/a4YuExQNLNnC+b5lZYgDE
ffYqYcaJ/C/XzUrIJ6VPVDVVyLL2s2+dUb3sFZqIfrjf7lFswF+jphAAaiclv/HQ
+nbz0x9qQltOCGAgkwqGuNTP2wFPGDTwdwj7o2g7qQZzz5/N3Z7LWCzVHoKeLo9N
il0cQkxrt0h7ELRx+ocn0G3qoXW6Ge8+W0A3uMpyoeFn6YfqfwPysPBgrbIkuYQ4
LA4L6/xKgln/ltLEk/nT8dsjcBRlp7LHetiFaQ3TwAUJGa/avEqjRztnq4ILQOly
VyTQDfbR0ykAscCGpQItu0pVjQ59QQXDw7B9hvCDZVt7NjVhILoTBqqNu26bltai
fAChuBd917Y7URbmD9LFYoUwZnwb2wZP4b2tysDOxgFHA6mNsWmn2gP4F1V5i8IW
evR0lqldRNgOHLdhlcrTa1z4uL28RjT7lj4r8d2Psx6Hot/MF9VOo5Abq2GIi3FS
oFZ7zG14tuBzFl+NDDNM9Iiil9jID0uSiBNQhkzH1iefOwssEa1t6P9wfOdlJJ6z
EWRDclmwQw1BZKKrPtqPf31N42zcEmJLvuTc9nOMNKMZspu0e/Yvdq26Hn6hUOk3
1a+JMxf/rMYxsqmiaV2vO1YvZXHXHyw53uYL96x0eDssnON4IU49RyYGxhHYgOFH
EfFomd2/NDncqur4hDM1pCxcNFEV/m4cR5cts0PX1opg4t6/ZAqYjV4rIBUDUwWc
drctyY36mBevbH6DJVfkptcTCdsNlCM/gVbI6e9Et0X19tDPOJ4v4cojZVAs+52O
bZxxab6BnmdEWzrTiEkfamQn9H7Wzc8bBrkyZDWGXwthNW9dVKtWyRztPnuMOuTm
KWRGwZdOP7+dpkAF0reS7G7L2lWOeGp24oOQoniXi7ovRN6p6Icwna08Stdaz/dC
dTunX4W4walKWdAGeWHsJOZNKxJNwALBzrHNKb7znECcP1O+mtW9Tt6FSzL6tOYv
gFS4yPRAGTQ7n/vbayvi0yg8vOf7nL1aUzsnVzkibfU8fwDiPVRG75OumerMcIYr
lqGHH3FAKaR85MBY0c7aPPMvRsIS5D0fOMQpdIWM23f86YzXFIC6QuM8MKJvtYyE
tLsb5WqlCsTPQoDEmTe1P8RKjz84fc1mihOX/XsJ/guFUh9zKbv4s6CtUPl+DcTC
6NRXDl9HHGYEPK/h5utTvnRgK+U2JyOKWbr4SDlEpmef/iYKRSSiis5Epv95FN1v
NCWLnolw7ErQoZiFgKKHaE59lZmxze1CmKzaFEy6rf/Pea0SpBRGoRRiBjUk50wi
6AwuHEw8PwFuuePp7UozYFD0IA7Cow9/6hSRK44H+0cs4vnwvfOq9GACe3vO/qHJ
+I8tpvGXFCsg/3dnvH3WCzg0s85bXgZOGBqZAZ0fcV9xC4v5coAsgMZ67GRNltrT
p0UxMxhDGhGLOHda+plJFKCtmDQyqFRr7t8vMHu/WQ83c5LwI2bViN7tBdTfuixT
PYdcPLkBE/JT4FWNJoan0SIgn66Ezu9mjAU772BMtcMWLSF6THC/csPgxb/EGL7t
yD8gD54kXSM9AvtV9GXKFXLaF4553B57kSXd5QUJNDDVvKIap0gby5wQPPMbbx+7
37QhvosP9XiLoCMxNoj85ml2Pnhv9C17VFiSGPpY8MdcddL/vVKAgl5p1mniluSP
Bf2mibgwNTYcqwW03hZr4uZ6sodlcE8c0PlpCbLjbCBATGrDPs4MMA275b8HuAK1
ygv4/L02HROGEgT9p4CkALidg8UCLnOExd48HbeLu3nwJ0or6aVCBc6PaXXmi44L
E7v4MPKdFwo988jRkBxlU6gaYcoWFfNV5hEWXqjC7JJ9fp14mWrGkNiwjCvptwyY
bhhtj74AFv/f9DQFizUMpKRvmv8KaLpR82Lg0BfC7fyQipvnwSawiUWsPJhWwia2
suHCN//qSeBTdE+iqYTRwBSVCFLwFp00gLxTfbWli3P1Su29xpNpEju4NlIagnz8
xt3YuTZ8DoP1nBLbiXCvsAaRAMS+nYwbqgnwsanojIoVdKR+Z12khXuFA0wMYd0T
QIR21bgh/xL79RWdFa+RdTm6zTVPnN+IPNUnez6uxHHawLO65NTTia5/X91u8Hix
CJjOHI4rdf/0X5cE6aR+0Dmfyw3TlawlueU0Vj5fTtrzusrhxOkIm8sKWBfr1L9c
n2KOJt0XsygXfBERclUSuXjooTTjjY2KCsm68ByO7LhQ9ytVzP363cJt3/95PNFD
AdKGQ0lRTXQElTvgqBa0Ikb3x8BKP0w6pBkZAj1gFPRoOd/vwrzic5zmhY+IBWWS
PCnu2H32Ptu9EZqVs50pTQNYNjMCKIZl+uCEsU5vkcTaKtWhe3QOh2VczYxhQTdj
SNLE2H4KwnfUoqd839OB5BjcysPNRPISbKkslkIyR+M6MsZBSNBfvCDj2yyiog8p
z57LYxrfrTfduoD/T5dnMtIr/NAdSGliSt3/vvt/IVgaI5bfsj16CDQaboMeyaeD
cyDNi6yjiV9PbmhXD8PRFUygjeuLI5sUAJctfZQ5nOqx8Yofqn6JxZQ75BeAPrm0
YN872HTW8NpqtFGBpR/R4XcQX7cGvoiVk4d/Jlk2aznOkFHQxr80KimY7oAdYFJh
iwW7wfnj0fROI+BtO5kPGWEysJC10GrQgNVwinfBq2G4yw3McnKvqq5LtUQW73Mq
4ZbIjaq3Hsd/2bBzz/zwVEPpcOo8oOhXDd2FvEHuq20lCu1H6yE2ZkJS9Wmz3Jig
ZxpbhpqkvTFHrxP9W1VQiZoru9Vz2q6RXJj+nuu1+8evNu8geGBC7rfKncjso1Nf
oajgBJA9Io2mBYY3Da3nsOjgJhkEuBotv5jRftV1tzol94ckYJrfPUf+a9VC44pW
ie/PZX7rXj81+XhXt3E66xERknfjo0lSjmR9vwhUx7SeHkOTIi81x+67VwhsPJGT
`protect END_PROTECTED
