`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3BS1qAAOZjkMXS4u3LyyuCyc2DTpKbnkof7TraSuoFxhjEs6dqFAysCVPlssL2zN
zmoC3CeU6O3aUC9n1VfA+0dI3T6EQEJofDvzanvdJOBGfr5/lnApdhE6ULsxvXAa
0YqCUYv4aS0Tqnd5fkq2wDIExnIGYhx6nmWdBxUpXnaPQQ+4aR53hmfE7Y6nWBkc
RHGb4sAXXHOPkUbrwJn1bVos7UtcqLyJmcZavQKuMWYUFOw/UqyCIxRiBNvA0L2A
ruNHl5VfUYe/PPn62fCsDGgrW1N3icA0NXNNZKKdikM0kx6xFlbq/zNA/gE9Naur
2kpMOxr8O8sFDqNCByZY6+NJaq4sCmgRqnjrclHHTZmeWhGDdRRZNK4ijMCoCg4c
a8yIo534TgGMUdRBWCUjE9nt2xtpVt/SW7uu0NuJql5snv+1PXMPCxZ5LsqMD9La
sgjxAs2a8849KJS9qDdl+BrgH2/g/v3WgFRaQP6srA6L7qSpLzQzEEwaGckHeZUh
OS/nk3HbaNgf2H7ZNdhUwO96XVqykwA08OaU+SzfVGtyMssdTfvkQvFCP9aspxNz
EyNJ+LpDvM7d/hSgB9yykkTOgII8aFzWH84/cyChjR2fH6pbS3b0arj5mpN+cc8v
qdOdRtQVqmaLuDW+D5MS1D8k/+lgSbT2USQ4RMZRa/61xHNfIl5mnhk2o9DXqHk3
UivB75fy1p/2Rh3erTo9614wRXtOBeHJlsX2g58KOXdfPnvEFv/to6AEvHFmEW+c
MpiIxTbQdyALsYImwuZYO9k+HmJKBV/28WfeL3N4U9FuuQVZsoo+u67r5zf81fTT
76xukknhpIU5aVm7K7iwsoqHmYE26oOKFdxWKTzc7gm/dhMlas8LLo07OxdT2Z5D
jgTHozEPsMldjCKeN+9T7xxin0SmWbnYPM3Qa5keI4tGMWfQNXuQvNT0XKwv7qBT
Wlu4QB2RHHzjmJsuGjBirxQ0/pBiRPzbY2Dl99pXP0zcbmBc4K2AqMdrC5ttt8+a
Zm2eXFpb0E9xtQHeYB/Bi5tzvNrxkFHnJYUcdhVEwuFkybetSYORob+kWb3gUEvb
+Iv26A32JeVwz6GbsC+76jlPtVzx71gWb9Wt0Mw/2EHUe5p/9yOaXJ1PhZz91yai
YLhECAYpHIJbVLQOLTcdnELuW55I3vu737Sea0RVbMK+g8lx+4VrWMliq2doo9RF
MDu5/zu6nElzsDZBXJ2vnzWXDtTwJ8EKgi1awqlsT8EFlM8Q4iY473xRkun4ZrcQ
kdDqqhvkPkCJV1DjNh1hTreaG6mcfwpLDfHdzuaUJlQGA9lH4YCZlFJ0wNJWr6XU
laU0TnO2DLj4/nEQeaHS69uj0n6ihe9D+zUsv1R6gufWRHHI+Gn4aumnRpP1uPia
h6xU4O4qfB6la2Y0wS9ngH7bgToAcZRKqNr9o52FisvNWCniGcaR8b1qHqYp4d75
F1Y+i1SFGQ07IFKTnkCRJLZLBSDwiXm8fyzAZgWRl5y3cR/XlaofZv5CP21kdXHc
ru2FtYOIxrccvM4mjG5Izlg4ZF3+PA+0uskMrur0kFv/wQjtBQxodFnIHjiLMN95
G3JpKWDXAldwd0o91Mx6nx+FxPB7BAI8FPR3Yk55ZPzWFm6BGNOMhZdfFMACyGB7
HtJ7UW3/cfnSM32c4oDkZUKijKjqAVjQ0VBb5uoqa3L+1JpoIq8FgssKS+B2daCW
RF4OeKGQZ9YYPmqHBSF1gjgwzuEGAUT0l8umbwX0dHzf/B/rpUBz3xJ9TrFszXQh
6LNw4iX4Pf6R/s3VM56iJL224iQLzjjIVmid0b6L1P+F7roJe1sVy45xArBx6yBC
D0EmjU5MAAQnFGgPv2Nmgy2gtgyj1m6boPmcjRCALPSOV7i9iAVgTkTTjwwwLCcI
c0gNeyC2w5Zl1vAaOvT5+Q0vTwqq8ivhd2qVmHraTPWweaNSXNjfq3Nry5B5Xk21
rILl+HiPiwH+KpCSU42q0IOJ1OuHkwZrrR8jPN5+h49q0L9i897mjTK/C/2PEDyw
0VzQ2KBk6gRP/ZGW2dl46iRH0TtI76W305YLzdwAGUKh29mNwu5Dh6yarAbWlJzq
HdGudukh9y1F7k48uhF3qEe2lgTT6aJItFa0SgFJSADnC9qywRgkBg05gZ35q+JS
g2MVbtmXmUsiXV0McBMHp1CjrLi3O0kDBQkrUtizT9y1cfz/6+fEiUONoFvGDjxS
FOWgnb+JmXOLA3ZGLn/W8mQdZHNGz3D9I86VYs7DAK6hTy3YDxnODzmMF/sT1wAr
aRnjPG9+9pn0MOucYLpsBg43WDr4WHbwbaXGDNmdeke0bsgaSHNAoQXmG9kY3i58
AK/FcpY++ioclVJ3O5ontLJbRISMdV7iN857mAMhTIeCA0q6R8TVWA8UWVL8jfAt
JRvKS7Utzu//Ca0+X57bBdfeXok6Nuddi/SH3gTa50nFm5vZovwAcLZ/XgC9HyIR
G5P/kfBkS9cQUqv+W2U2wMXwVuxpBx5zT1mLqHSmTqPC+nSac3R70KQ1u61E29NQ
U5rTmLI0zfQuya/dLRpk0dYJQ4SjmxLkzcoPppAuAK7z3q0VgZgC7X0DOa1cMK4j
tW9H4p46/4lpGoMnZR/x8eMmVW6RhSF5rB3ciBR/ZsBVtzFSgM7F/zI+xuzcl/8P
mbmot/Jif/D1Q9tDJZQGvME/3qmaKx6/k+ejCF6HznI0NTAquYPdUvl4e6GkabgZ
J8mLFreyLyzVpwdflOpujVu+KrDSVhmvclnhDNXHEu/Wh49pbP+zoMuZvzNHQD15
MsLVwKnjgtahcxxus4UmI1WD7epEjyTXwdBILsZGe/yGg7zGSs7u2S+ANleO3m+9
hABEoDXnp6IpLjtQHxI/Ho8x+xA8Qsf8s/q1VPsGLVdtlKmvcrTKHfncgMNmLT4O
GhloAulHd2CpLQozUy++2XJReiSf+hKnlp4031HPMSxE9dvR+2udRHkipIUOhr05
WWJVY9jU5aWzNNYCplMKqT2ZV4eS416wPtLdIuR374YSM9FvRE0HxFBIUwDDKa3E
+e1t5DjFaIV+XXM95q99P+nQ00S3Px1D9vJqeYwXbiJGO1DfPC4hub/w0EBwm4wc
0vE0EEbquGQj8Gl1c6qgEeMShkX8dG0BJ7raHwejCw6PAsIGyJrxUYCwFxi3pklz
xl+tivI/2ucEwTXTUA601TtaLdBEDV1qg9XtuWnSA6Q+K2ZjPieV7O68o80rRNz1
LHFmlLzcuF6asdd+vKbdOEKxdor9coe5gV3fZeqRz4dhC8AHRv7+hx8C6RGZASXq
qVK8zbKvC6Mi0JNXscMJCRZYH+r/TFeQZf3JatQmLmSYJUFWITExdDZSli7If6Z4
K6NyZDPXMY3jGwtQI/JUTNd+NRWUVdJ/2aLRkQFHGMHMoEB/7weLzvsjhMkpUfiQ
nY2CwDNiZ9JPmAHDCmrnVDaXY2tvzNO6kTy6PKR5iUJOaKKs2gG0tRnsoes8u3yZ
jxf4qxqpbVDwydxfJMvmkobbtjI+R6j8iDsnOR3TRetasuJDPdeEcwQQbp/3fMKr
PKXlYJdRoXj0EBBHGdd54NzRw1gzCRPKF94YnLmIJoZ6+KgCsKUSVmsdfSzT2M2C
IqSgB5hqfl494282IqMii3jSV39ikqpMYgWqDOXNzZqJs3MGOSgeKMtfDXdefRTL
WlNILDYV/6DO/p7zlRiTlO7sPFmlDqK1U6LnyxfpSqJRcmGFZQ1ieCbfapwjVnvZ
sHTZ6nl1lr+ZWwVNCX8F/xNeOG4LyNC1zwzqOM9s8YNRH0aBnp/+Td4VsmSZpuZP
03yGTb+ro4OuryYw9QJ8+CtPB5Kobg7WUTAhBnFh2qdaGPzVzSPWP6FHGjgIOskA
N+u1kEwfPEzFburS9hv+UpiGuxCqqvyJiHCsYRadV+RFnNCzaoyJnn/CcSBZqz22
f7W4+b9/DNeYbtj0JfQSmpYAFtTOGfiBxNRQdw0BwltAAb0t+YV8IAEnv4EvJIlI
SNsPFzydX8l8oy4eeJTWtSiQpgiL14daHKGu4pyvLFPwWvH95zrzUeOEPf8+vLkF
OSnp07yK4k6Fp+zmylLRwu0xlQkwZ4tGlrw7/SNIW+0+8sFraOhLsq0qmjVyAN3L
qEIXtwOswcfwy9O090h4hmJeauAOr7QiSTVVBLdgB2bREyk/JQiaeR307ezCTISm
Sswl0jN/sCTW17clwwTXDX05pa9aF7XOrf0h9GMlVpFuaKTd1NyCcaZbMLWSqt2h
NksiC+4Q5V1xG5CjRcPOAy92buZg1hvODnMpqASxHLhvM8bLlb2N2I6Co6j5HP6s
S/a6OduZeO7Tzarf7l1qypC6xuo5zJOnTNX1B9p+X6RuHQBLrNXHh+Bu13+lM//O
9py7/lD5zmCra3CyVcBsEamsrmb8/mhKmpp2XQakaeIBd2s7MJEKLQNwjNQ0Vh9u
tItSUsh26iJa/skortEEsGtTDsIb9fgVk12gAnGeonMaCRRteel/O31PTQEggX8y
rxeTH0dMSjQsu52tOeqttKDM+W+/OM1oP7Xt1Tm3euBgF4dtsCAHQ6Xg5hMQtc9t
Z3hZSi3NDnok36KCDJcERoN7gMH9lJzaQrWm6vVNND9GXdZhyouacpk6CwDddMdx
/NFiLWneru2QDWzAhEFEhgjYPNFXNgsbEuxwAq8k2c2ttWfOv+vJLYbZwrbeFb6I
/DVtF54zwWHDNMcDQAziBvkHu5h+6W27pSyp7P6PuM/edcsPtCYHM4irDuNuwBTF
HUNrH/MQegSCzKf7BEaMDigv3qLXL8AecNSlGHU9Dobf0wQMk3IdFiSAPkpXgrYf
GyhChOXIL3HDCySuMXmQJY/TPd4NZuUJVe8G88HXpRuwTOyTLm2XjPo9vind/eL3
xEpUIlII+jmQzZ43eBlrvWD3ZmeZk9+ElJ8/L6/M40RsgGaEBmY3XpZZKbB8O1MX
KRp8yb77Pw9wJnHmGVo0EOugf1KGfD/Zh8bWXD3Bwr7Y22d5j1mg4N4NNjQTTRtl
y0LU8/ef+9uFSW1Cgx+EXruc14P9wrDOd1SAx0TqhZ03xZpQQhtdmsJLdvw4CsMh
WjayKh8/rNSe4W6EwREhW9uoXqacGuiML1t62tqm5wd2wDcdodMe4k7QRHcp1aj7
AQk0jcax2dMZcI1S0MfWES2oXYV3Ld3MyQFHAkmDzjLyj/fxISsOXl7G1/S6zHPe
E0T7TGVluLrTfj83WpqvzS/ZE7kp9vR/g0UL081TUizTc+jd9plGX6THRrvL6cdy
6+84V5cMN7b3SENup4bIRYWIDErQgiahRtcvprW8Cz2YNpqfkzbZWU+o2FjYxHox
BXHG5feeI0kJ0YqsboBAX04SB+gVC8u/ySvz/a4ldyZQtmVig/Bv1+jkQEYyQ7O2
4S3jYFeR4I13tA+kyFjpp+KXY8/pVCZGMtZEETQZdOVvet5k3A9DoCoe9yeDZuPA
O+HXoyBTrW1weRkhtZ+UhY1Eq+hNNF5hEVNSZziCVyRZLliJ4qcUViONxEHwf8H2
JeYSqGbjQOk2prEq37kvN88Uj3ZpSpGmPBMeplQpLIp7IzL8lm1vOA+yDWpkVOvF
h6ndxTr3DjQMRZP0eECW1rUejVgCOyiUbe4Nd2WNkYrmJaleQu8dG+Jyy6KBEMOY
H+LLJOwul51N1I/iucEDFia3G+MuqPDmuVyvbzm5qYuthx3hXh9vg6xHq8iDLJOw
2vtHgAxsUZ2cH+95tQREJR6ZTkjaOIgqdH+4JwyfI3ChIcQriZZ+HKOjDVnpHHes
UOnP8wcE2oIVNqNRh+zwCDqOJtXkKyv+ACHVY0ArAIKSBAddHELE8I2mpmZCMY3T
fiY3uW56TLwpjX9I9btB7vHJRQbKIb5X2oJ6MTm56L0e98uuT4IZwJuhr+vAl/zy
thcck4XNLMpIvhH3il2zU0jL6AloWSJk/uEAWoUJS0ZRZ4XXRPyWQSUGufvuxEwn
utWqyMu/f32Z4b3jXKN5zwjRKKWrI1GS4lxaPnCvYzFyWf478XRoAOy/Go8fXBgA
9DcLs5av+V56bthNV4ciJorocZQge5xawtPmny9h35Nq1Fm4HEE/qgSGbdeSI5IX
+2lFWuIqmY6I5UJu94T83dPtnMm+EIycPjmc8CtCjIHabP1ZZgFf9+RNy7jqD8tq
zqYAyV2ppfyT6LMiYnW48pyyICSlj6lz/fDR9CLsnKV2agKoYzhrJmxOfpSBTHPW
lodzgXCCk+82KeukRD/BY4oiD17Vg8ejhvCnW8BKjNuTdv3vfvgH9Ucml6EwP40W
XHBixaj/Fk1Hn4tyj4J/VJE6KTWhsYvK9tV0MhphBBIticYylbmLh3mMgJcD+aPF
W9eMi7kGbsY8PFjYfoUyhAq7QaIa7pOYZ5O7+JUry0SiKpF/hLpDrSFwJZwMxJrn
tPgsFJRISbe1rU4Kd+cSouJvAE45y3hzLqzNApW+4OlT4fgJKu2RS7ZbzimvX7Lg
x3LT9xFmM8d6XIqIa1RKYJQoaGh8O1yliekLG7he/d26JWH3K/SAu6hl5hWGamER
sUF5wxbDxrO/K9KoyjhVzkClnNlRWc2aQwdvNC3gjvbXOBKComRm6gNZrMakZ4/f
o1fukqi1+xYJjDwcPS4vsKPY8xySil7myjNvzSUfbfDX43y7McOEfJurg21gNQY6
K9wTqzi/UGo/2P2ahm00kVL0s735Ohn0H88beDhUtuvV9GLh82mo+SRa+wXpvUEQ
YU8wHK45f9Ifuoll6tc4GV06Hvd8hmuXu/ZqDqGjWgLs/4HXDTsMeca9c22jJ7B+
sF7TVadjGDFcG4H2t0+6s7H87kNAsDIkdb7N4KglxTPbKvixF0aE3bbfQq8m7f0D
goquE01EY3lLaXJRm3d2Ppqs/tVzJKLfsfTq4AlXOGhXV2PSlHxbIhtRIs6a7hYa
M/elLDPW1iulszodawMMZBLCGSUx28DSATL3yOKspN7rFBZJI15n0srIr4fkgtQ4
DJfFW1G83qf+h54v51ifzgcxPZRRmHatkcR1RSZGa56zNJyrUOlk65/UdD9cfenA
G/hIoglJbHCHoc58AltL4rvuuXQbRtwUbcw1p1mCrUu6I2r1QWciWSoMKs4b6ePa
4d4asAfg7WxkKmKnPwdmRtX9o3Ff+p4Q1YGS1oE4Z5U03CkLAqqg3Q/8eBwR3Tpr
SJUNSykF3r8dPQjwxA77B+Wlh/pNRFGLZpUJFspHe9No3V1mxssGv+XXtgRAp1Jh
f0vSgdou6Qc/eQuawdSrmhaf2bey0mtZXK6da2hiAkgoISXe4LprBoJcaRBGbR/q
iGpgSpKgKzi2vDt5Z8eXXBKCRh6EKjdyagAycHjVYvL4FCrIfZg/2OTY0I5EYP87
0964VGNlWZAU6KzVn0k0djs3kNJZi9pFZozt/sMzPFfj3m5ABHTTs9pXTLXL1+OY
QRCePjZFknOa8QcVGe1FegegNAE5OjkWmBRDaljsHMP0cuZml3PaHkCOQ7IDa0zP
uP7KImfyNhdsoYrtcGDxauPWJaOgnrFV71y+AJ21J5kJgCSQCFu+UROFnCGIbeZx
77mxa12LiA9Wfy4OrLIrOixu2eRFrHj8DX5ecewbOa1q1X8qbKJ4uQoCXxPEq7S7
qhr9WqGAAs9nikbbM6BCzAwKi2eC9jxNgLeg1h1xbdl43BBvcY8Mx2WWAWkCqsGn
V2waohy8hx6fjo5I1PPK0ElTJD9W03xMjpZNM+Siqc5r04J15Miw88XPQs/zzfV6
VTq6RXHF8Md7HkKkuTjjUula4VDWiUP0V0+gcG4MHT3kIbLQOI89pshMeLk8vYu3
N9OEzxS+wBlaM8Z5Z2umKplm+OSJP+XZXfFA8xjN+CfLrVnr73TzjE60aMwsKJig
LyatrjjvaDQeTIJdBL7mKvzM2YRf1mAz0vAbFvtSf/fci+odGMt+eRiDmMP6/Shv
KW7g52hJnHOiiuI/f85z22h6jU0mSdleDuYZYeuKKDOG1WHfibd+W0exfJ59gF0B
55JvvZyJ8NvFwSintEGqsV6C4mLSzUX+x+LupwICsTOBlqlf7QhOkkszxJIu7MMa
5VSLkYs70cPaiIHTTUSERvcYVPlA92LFsycdusCdGZpwuEdPslR4Ub04VOHI3m7o
r/Ep2KeLSx9vSCYoELt3VwvXHwIda521pnqe4IK7lkk7/uJUg03aFRLq6wxG6Ewc
7MfvGm8t4lSfI1FPKeAULQsCkmJMt6+uWaKvPCyYgiHbvJQYiz1IfAmUPGVSu2cg
3kgZbvXNGGnNm2iMMnlSdMmbluWETlcXNHkn3ZwVj1M1iQ2T6tiLgvFIau+1mXYD
y9u/h7N1OGi3ebU+etYubiGKJ9lb6dum8Xq93O6cgqJ7+MoiDrrQ0xwMlJQCLzkO
1/GqA6Y0gAy5BBdZPloOPmWl7J2o6uO1aywFn790JKr8luXeNR68HRQZYxQkKxk8
7Bi7PSuCiILtiahZAeMGV9f3Ooa2uHXsHFAjaXs+MU+im2JRSfbHIbmZZH8KHmQ9
AddjYyXjDhUTfiFQT6ARAR5ClyIjziPHp09U7QZRqpiCsBx11xsOd6ZCGOlwzhvr
PM9YGarHPWie1ElEOrDncLdiiq3AahjHDXbRBSFlynFZm35OYIy5GQMiIP4NNStW
kTYWrnWu/DCZf2P2Hd1FordDkfTMQrORciCytwKLbN3VwHXpkz7jFeU3N4oKxGpH
W3fpL83+Tgrn3CknnTZ5wQwILeVhQDzy8Cj7GRx8QUkXKixapQJP8agaEK4YDaBC
zWkURYGG77L3hSuzbgnVhw/ReN4iJshugPXo8hMzUkwBaxUhf5YPAp0GXn2rHOS1
OOd+HUa6hXxKMfeTNPGsJuIK0YCExS9wLvbfwi4kW2VLh7mPhc0s9iodnhi9KpVf
PY4CBamRVSLXyUWwQp+c4mUTLTLfCwvAt3tYDF1LKJ4ZQMnkVlqSNhWiYCFfn7kH
gvavjzqmnOyTU7dNuATG6LbzNEBhoZUwzD6u+sejeN5JMpouuH9WsLt3Gdxdp3qb
EoOYAjasgKXooGlc3wyuc7qMZb6DrFbGqAmjDov3YkJdsjftaNzf1w+Avww2PeX3
UseW2/7fnu86I7p5NBUp3Tg4RteQYVEm5LdxZjXLaGxQJivoGTRVdqIjSzytKUec
aeFhXn9ETigWTE1iQhq69A7/RIiPVJJyZjW2ma0oNl/RrCmjL7dCqvRsf4XoOkJ+
CW+uTPJbA/NZym3LYbfWMYm35UitN0VN8noMF7dPGMdLUg6GwgxcdKrsOEuXc+L+
Udkq0ZJLaxq8AQyZnLKCfqbL3c1Ip6xF6Q6chbp/Wkp+XZx5GvUsooAdoUau+Eys
z+KSl2xNXG+tt6F0xKyTiaJC95cnSclHH6kAGSkDrzJTYT+R3vXqGxl0BDfa3NcB
yHmnOj2D2Nbqr9l/y/lWXFn4xJoO1iHDkqGzlom5JpJdyuz1W4y24RsfJeofqWWA
S22409xAgNMrZQ+5+UXzwW8Xv0rNuVuYUF/sHRnFEMaPw5tqhzwOl7wtOGMuW4ji
lDlJ/4DCiXDfBOUNdvg5mT+qMBYAnaJwNV7zbQ33ZJvVaPHa6PX5EFUvUKzpU2lc
emh53q9KvIogtNSVHJ9MRZ0W63TAlZDtw7wnm8Ps4B7bdnT2K6PFnKhjCcBqxyD7
3WFHxka5Q7NLhhfLg24dOU2BCQQwXrX4O8v0z2WOy7kDIUZhtObpeMH+IhcdNNkB
E63AZvpVHY1MFpmo5M3ZI6U6ZpT0UxgdY+bT0hATMojiNpt+QsDYPPaW9NsYuj3c
GJXvvDfDk7SHL70vjrCIyeP+0dEEQKIr8VmBwVQGz+C8sbUbSg8N75ifb1PnctS4
VbrsEECqhFCEme3BUKxZlyXa+SU4rH17tU2Wk7He3T6NpYOzqZwZMXUbp52fq1Sy
6oare4O+W7w3Yuy5bwxM0ii/ygOtK0gH6kqjh0jX8QC4hFeIS14Q9hAMMu/4o/Ks
vGKmhOQyyGarnXi1F6R65p2yuPYYaiqyrv2Ah2lKX1PunOAeBSfHa8Z5UoFdKjzM
krBEptTTp3gZrqqLaDnmTQ1YBMn2DqnbXpgIiX+RJaCjklA4qhUw4hTSdPnbhT78
w1gKsechRT1Qn6ItaLB4pXDMRCI/uif1xcgaFFDXYp7cl/egNyVgAvyBjpyP5dS2
6RDoTCB8LoW2fxyBz7j9MlxVvO4krLxM2wDOUEDloQDjRR2aSU9cKJyXQ0AJQ6uZ
V3eBrSGML/qlzfCpe5DQ2MHOpygz96zuJ3p+WJQanJqqTnBIJ2GCIDttCRdnz056
qf0kksjHEh8vggmNCdJbrsMMRi2sO20l8oI/NvNbjKq4lBLAprh6E7KVieQCuOEI
vcjE591a0q51SXjePy2kcNHNFAY+IsahoKQiAkUVLnNhFv00ctSee437afbNQ2nt
pqVpRXx3aVgGEItRQPXHNCu73Ega6gBUj5cJrfFBw7vr2ParEVcUmZlEg0fuOVgW
e3kCMHFD+xVwd/EEYQLLftEARM4NNyWmRA+UN8DxmQPD7kVWGRsNOnO7sxyl0JZa
iILCwKriPfWJlppgKJGwEAlRMEL6HN44vAnRcUn569AaSRJ6GwIMWXzQATKFfpt6
iWRswjCwy2l8aUXOsFGNPkRKeodjB+PWOrh0COxkOB43CC+9S5Q27pTlB9tQVBx8
XwdCdljOE0/oFYaQCdeJ28CRt4fL5xDUUMF47pMKpB6nmb3qoENxd1FruVFUmDQc
fL7mMTbir3fQH2X7pz6nXw5deFjEAv6xptxVlQq+PR4efix2CVXXyvl74ZI58D7c
5/HgpLu3dKICjCwMaHFEDozqcdc4vUsanWs69GkjaKoYrQqOvaMeZX+aP23T33oM
bxDiB4N7D8ano+ekOnetIkHzGWZWWiTnvLGsgkCfl1OBScPjylMTFE0Sm6BwIxvH
iEgEGpewhgGUl2tJ+hUjQzDfbaaL4ZNDpKx4HTF4fsTaMbu6dtcfNy/AQZM4wtRh
oXQRrgd+BzHLBogp0+ce6GVsenvFLhdSLAx0R+jyKB2nhwxEKcaUGSkFzHXeX4my
79Zoi83ygpPnfJ9RrvpVMcNqvKdrEBqQAc5JqgCwqXUnU0JTDNqE78Xsy0ru+vn3
YM5WR7CR5t4wGpIGk1WH1WPX5VVObqZyJncoqyWV4wC5ko6pQL97PSQ64v2O40tT
Yjox3VjqDMxSDz2yVw/n7t6ab8jbKCmzdVs5VbLwl5D6nATG9v9KEf/yNZGP9CPO
TnrMNrhtZ3Df/6+5R39UzriFxv5fphM+fvI3x3XrPecOVCy40rMqbbgl2imU4+v9
IOyESYCNOQfQB9EnPdlMFPdFnH1VXTiEmimlpwXRoDYEoe5xsfSdWYL4cYr8XUHz
gOtuNJ+1HhIFmMv7oP63XoWNrcggdR6eHWCXLgwIM035JrMfwfTfIFuLZAfPuao+
P6ZmbLGHZdFEAhCAFUqL5uo5vedSzqWysdLzyIfNnwO3onyMsGtrppRS7pq21JBC
sQiFKH7D4y1wuk2GwhCpt2fg2/pMDAcXA6qLgLZM1LCCoVKXJ2tNF3kMX5bmQ2Mm
Imj7i1mXXsKsYKuc2jbvooTvtvlkHsFoUB2vTfKfe4tqOtz+XWidkzb7wztfFHFg
wP/UH+i/P4wD4DE1InrhForv/A8K4KslgIBPGGuW6ypzOY6dK23RGRDq2AH0gzWy
n+9QRky8qHuxMfjRgogSBNSU3ykZANZoIMeyNGUEkcF+EDOx7QHstHT6PwBtf8HM
eEkvALBiw4UcaXmTPHXk8m2j1KKmQmmEfxWms7W8oZoOvwYN6AqkxAscfJA37c45
YRSanvrfB9XUBV9uwGJBQsqXeSf8rF/Svck6cHWjbhxEQKn8SJk7FIGXlo7q1X8J
jftiOm/1A7wBaTHTFP/6jqwajvimrFM6HOUM7iY43CA42C7MzYDGkFAfDEH4uBz0
czoIOFSG5bIpHw75l07QuENC5ZaOvovq+4t6aRoZpPuyP24mXQWKiW/78RiCivb1
fdNAT+8W7jwNpp/2bItRiAu7MzLGh0djv2dcRqgeaPVxycam0j+jkWEjW77TpZMs
M7/Z186X1FZIrw0nvC7Jr6K85RNPT63DFxBSjknQm3OqaGImsLGdFCchbUfLguYA
A/QFzT6us7/likssbetT1j3D68yMo/S+sCWvSsmgWwgJpV0QCMcPUiWGb0Pa52NO
9Kl8ebQJB/QnF8tcdd/Ft3xzwTLzcAgqRGKRVwG3CZxCjsB6R0cFCQGDm/WyKU58
M3CZR50k/tbwUuHwWXza1UDYq81EO7w0g0smJrqp+yE5+Q9IqKRxZQD3teZ5wNNz
ktKtGX6N++eADQT/Oe+l9xPT6vMpY9fMjN0A2OPjEzwDDmPzs1e5ThTxRvCS7jVw
AKjZ1FNcTvrgSHRGEfqP+pCRkV/REEUhG0ifkkYTswSuYQKwtALMDKmp0fs+VPEY
LOuJyt0y3dU4+ikno7/oDTSPbuj217JNmrWlkjyq2CfVOqKJiGNZwVgoWEJ0M3k7
rpaso0BGY+md207kAC0AZyZZ8LLxvD1I5vmU9tTPkbjFE8TzDphl4WOJsXi3ARPB
OYOD3h1A/ynHDIOMPgBCmyohgS4wQdlFW+BX/GEjyX2SY5KKQLzEjTEwza8xTPbK
uNY2GgRri0CuLT0n46mUZUZ5ILrWRFKguQFpY72chLVTcKQqbDXC0qsGIRGIOdpX
h5erm8bcRgtsGAyyl/jdHZlhAS8Kr0zj1JRIWCVBZJ1dGAT0NDOa5nVXHkBYd4cr
MsXn4/4JJvdEvvxqC5nvW89l9tE2wnVVx4IRJylXGyXQJtX5Vs3awrxkIKXMq0wx
vdECo25bIx2zBMSGqPf4nbzYAFMHwOFN2OMKyaNnr3TZ2ubgcV5I7UOquymikW5Y
FczX8JREeWdn+CzronbGsNpB0Rq6o2aRn+AdD6uCl8n3fbVxajaaEA5DZ24zE4iJ
Uu4vE9w5f13IbseRR+fmV3MRUYyxUCtReAUnTLe9MoXA+e+k363WkvebH7EKyizg
oma8IXxh+t95/m4ukr9/nu/2NtDFv31hgFHnxEdCBS6Q0HO8Lcv5soqi67n0/FCM
8E5k1QMvXhIMY7e97ygPOeK0P/a0rTZfjuCFBH1bymImQd8RN7u35xl8MbfZVc0i
0Q0oc4k4PgXruVHNv7BfkDVnKaUbFDfahDueCJvA7ji23+6qjaqoBCOUl17/+hej
VRSz9goCisefWV6nQk0zFKgLRc1ZXIU5y3WYfqjAFrjC/Xlv07MdpTnsIm2IT70r
zn34DyiYNP7kjQn87ekEQ4GgS9I8suO54Re8AWOkEFGOcjWJCQpuRgnidzZp+JnL
tCDCvyOVnYFmia9zI4zwkCaw1mSgSYcD6qi0gWa2XvOM9iXWctoi1RQxXzP8m4yh
yhi8O8niYV2Lm6FxvCT7vAd1a3wIGIxv8SytA+GEdD5BCLruaBg45mb79+94vlbJ
1+SUGGisU81b5skZhLdvOLG1nqKULVV+FM9LNffq68LptFKmgCZx8hU7x4ncwYZP
8gJ7YkhSfmw3ngxqwafJM5YGw9aEY8wzNZUdvcEEbZ8Hx5R41mGhrWtyb+yOIKJG
iZxy6BQFSMAxDqJ7qce61GcuR6oeq8pk8oLr6EBSwQjNesMiJZ8NWHV8hGPxrcyI
jH/Exsbbfj7ZuLd8fE25tV2YcvfTRZ1CmOKHpk1KGetjNm3n5Wpf7u6LOGtuec28
rs6DlhgizHIq4KawnchCcSXx1jSwEILT67dyzofips+PEiN6JTL80/Z8wGHgFSXm
dP7uVDVv0cMsd3dqKdTqUBARsMrpGlKFKLmtC21jJwF7w+AMxm7O1cJNVq4VEPal
J3USLdgnhmCa0bNSnsTjqBuYG2VxcBR2KM1kryVPVNCsUYEANfXBV7+ejcDHh+nJ
aNuz2lWiOgUKpT5W70LPa5I0YmdjxIwCOnzdfDZWlGj4vpsSbVdxsjvPqwhPZ+U0
B+/jYUQwdjDlkqB2upsJY96PTtOze/AUeUARIxRrGI8sCn1PtZiRnn774hNUEyTj
dcc3uaQc7F6spES3SdIibw5xQghUzI0ZmBoi8HZhLo0PmMuXm86KGe7mDdZDWH9I
tB6CdZl9UxcUHHbj3ctq+8mfvhNfhvpyRL0GJjdEmsr3KRDjuisHfGr7BwFdDsei
GzQYCAlME4atDssXnnCHJRxXHklS6jU3wUFadT/9Wt0rHXKP8DkGsapJTczX3BIl
JIio2HMPP1XHUI1lfUC64jpVR/TsHef0J0vr7Ejof37B8L4wKZMY9zN+oOSosUDg
V/jo0l6BaWdi4qzqMBPg3fb8e86XgLl7KdUaeETIu2MrH1puXE3u5O98LhBthEdJ
XLEYOofWxaFoE+wEaTSR0dM/fWMIpO+6IyB7r5Je4IkSermT2+eGhYcvLiS7cBiQ
UP3sj3GgJT/clAqjw8vsIEzRhfbMD8F/w+IQA2LffA6Bhv9X3NO2LgkB4yGdJDEK
zsXAHWw5ABgC7a23P/Xx1WTKxqL9wJCKpTJ6jHWGq+giCZCB73rqpfKi53/BseDP
9ENk1Yd/hjJQZRPQc2JuOz79ToZ7CUXi0rgCrjd1353YUknxlNaFRIcFZNBQbXgE
k9rymSKiueG6kHLAofAhJ3JHPf+2G//SHZqgNb8RXm+kRNHb6Cy2vi5kaPNzLXeT
pwYQJK0q6Q/9l+SFeol0R701g0Roc9jYkPNg4/nlmn0o+vjO3IjK9BNI+07Osizz
vms8+0aBWwgCp5+81hScd/PgxtzoIyXqQuCuO4F3tPo7gXPb/mw3r7W34DjfkUnC
Xqc52JeoRMzDc/Bf0vZWz9CprN3NugCV/5HE8feY1rHa4bUFyRCJklxzx2XXL0ot
5/9cFfLREF9oSHEGn9AyX/v1Sh/n9LYEBILM9Z2NWi6W3osQOKPjPV0MBG5eN/ce
dgxinBcElXhxEBGtDcbbeuGJEGWMEF74XCpn7Y9BLTv7hEWABzGxk822zPS7bbzo
USQ/Kz/6SauaWbKNMmIR50mAIqdsLvQ0gZncqOPlFLMPHxPpl5aQQ78jLtVtVHmZ
E2yowTjOH2aXYR7avJslHZEWurlUA7qIlIjP25dCRSo93j225Rx38n7qq+o8HYeq
jqh+oDVLHSQIY4KXyseg5eBU92U13jPTTJ0AGbgUyymAAZcL8PPNH2JCs+s4Jx1k
z41h1/+RWadgoAOlG9Jm1dl1fHXG2KAV20buFQuHz9ODpNna1BRYzGKcIixT7BPR
h4HoL2aYghfWo30KAqwRgk8NYWKIdSnn1YH4jQBZUshU8gyLUIGzqMxctuViqPYq
7b/oRA9cW5WE3hQ7ezEuB3RBXB7DyrR5x1KuTvmcdpl98EoE5LgQtuLnUxdoJ5rF
lzDUkheEhlwQdsQb/pYCankSeOjybSSerycIkWbpQo86fqI1kU2IB78wOar0Neto
dDd089Ko+jEnEeCxPzPyzZPC+b7TXUVwPCY9ZAWOAyF9Uz3NYjizvkGgxmcgeuNj
6cU85BwbKD5UoHaqAA9PdMLsmhtB2LFehjDSPU7m0IH2p3TsbKM18skgVbymy6zv
vRJokoFrzwwgToIjfBs9Nict9Rqmjml8515AXDhSZqFUrg7Ysu12JaRR153SPQZ6
kLuvnI6d8PBUEuk/Ohp+Eb3AH5e4dSqleWTHxaNSbBQBAHZEP9MDGMsEY2rSb4cH
kUdg9ief+YQjZ/nKTi0cJ08JiaACzkRAzkaDnBrPMIqGl6YFFdb29MQiXw4ppH7Q
u0eTOiLaZyv5wQym4xqVM7l23xGQVKxQ4L0vdFCvSED/k23U3qTX/n/qObTbO/ul
fGYdTkE2e7giRwCTNOLMWHrMENaepkqQNCZpMv/DqJsnxFWXf7bGH5yibCoj3oVG
dg70/E29eICBdnoyLqkKwwWzUJ0udiX8K1nJdyH9vDqarCnbpiTlRzuuRQRnMyuh
zRuQV+ZgJHJln+s7SQFCbXCbyJShZDM5DO/cnKZrfzVkq9MlcA0O3K1msBN/a6dg
JpsKLfC+UtViVGNhTGaJTw1R4bf/87uN85mRzKZaVFc87ZQe2QqgSXy9t41JHuxB
TtX0MyccJbs+kwL8WwFjGcXfzdCjJYCCtPRHlRJn0BypappyIIrNGUFMySxTzOpf
3o6VPp3iA5qeZoIGnlh6J+6R8Cdr5Hn5uW5X/VmCfuEVfWHel9lN9uIFbgUWugLA
VGZb2/e3i5yK4lQnYA48D29Q7a1U1WTJa2j/wfpJE+y1cx3X+PURKnT+zvy+1UhL
cHVS8BAeCi0pkb4B0ucC4CxhXGIRgvj52W+m+iEyw5ZGSvOKz9TSSqHtQk65DKmF
rqXTj916lccppkP/G15bhD4n3omwAWzunoqBm/zlcQyjcSA4ZJpEBzo53Lyf8Z3i
B/eTAQCgS7TK1Q6TtSvDKkwE5Qwqw9Rs/V4LWYYKP3Zq5nHRxUf85zdXC/G9BtD7
02i0fqI4pb9Gd0Y91mSXVTbpDMl5tELiMe0KYwUeu56CC7KxxmN03txydmJrcjcd
4V0TVZx0JfR6MZKjN0GY6mTjF81SXyuggNhqPbfgog+hYmvCcLONFxCdmZerDk6b
/botZ590KjvA8ldt5sVFnFQynMag9EK+TyUoPZO6rIVSfejdnMOCzyV9gqHTGXC4
9AkqnTJ+lJVKqoVDf0uaJ2JPhjASCltGUwSpYQB9N79790HOGKrGxTH8S4cCZJZr
3y9lUlGWs4grypG7gWBCOV7kvUW5XbrHnbuCTMaTZemKuF/naQUvP6tFz4vqxw0m
qAZuIez1V2F1qf4L8HyhOiTUqRLM9eYDiiSNkW3i4QO0NdNb0Qv8mNkO+Wx8KENw
X0f1hSB2kMz6ZQc8+CE0rBbmxjFBh/gjDYoyCH2/U43QVxbkliwvHZMgNw2O6D4+
4xXK4OXPbvMeuNTUE9feP7QJeJm6tfI1tSeRmiC/42Enp9vgJ01LKeyzqwhbeq+z
1E3liQ3A2gl7KRjQgpqwz3FwcvR5587LawPxu3r4hqyTdArJ70Ztn2u+l7kyXdJ5
20nIS7RywV8ZojRZDzTVn36W0h6+MrsFf/3Uaf+4fmk7aJd1iXSeUmXhw7ANBrpL
v0OJxrsYi7z5rYBCj94gFurMaUZ7vo7i8D2DGzOpLKHM02HS3ZzwqdyOyFmzmLP3
pJbR9ARLj3N6kzbOGV9c/NVeLL0mjqQ4+kk/1ymdktXpN5PjUbon5h5nJ/0Ibfad
uiBJagv/cqlhfqgF13x95e43DHSq4Eltn93mzH8tok7Q6NEA2Wdvei5UIGxQIwak
mSBWY7ehSmKZ7Bm7BYApDaxwFchAerO7UV+2AiPbpWoH6921QqxhrqCeXJ4v7SxO
EGq6zzBzjcEWRzTboIRGRjQR7AbVRkrMARUaNmkjF1HDp19oQaMmLiuR9cg6TFHK
Lrhx/jTU/4XEF+WYhbng2BKxCtAPCMGeiPH4XYpsvBkH1UHSvDEREVp8hZUBW/13
8BQCnUOm+9Ftl4tEGMwmwuch0jPu+s+KJTwWpBOTA6bul4Vi7X91xZHFUs6LsiXc
mrLcx8bOza5XMhJBApag7PJjinHyts/A1WDFtJ8RmWPdc47m8y4/DAYZV4lOysUj
2SNBVx/4LHv1sS82NLHh+8Yh7AeqDEcQRn896V3mOv3soPEQa9sbz1F36ObV4vSn
+s6WQ5Uxa95pSFy11hjS6rUMjpMj5edqC4MQfM9Z3QapUY7JRVeAPFu8eUyNeo4a
Z09e3yVf7CdYg0i4N1I8P0baXxkx1dNjfksGHkF687Pm59VMIjrRv9pcSTHvIxpK
EY6gZIcoWmLfjBtsN7jjnrdrzXgIggrORe3XjMVsURi8m1n/6W8JsMsSGv2NAu5Z
uZeI04wVQVWL1jp9MnbXt7M+Te892F7bkR/3iIkoodpNIlmIZJsA14tXGo97ZZ/u
f1haxAq9z4Gr8nJcqVV5Mts3UqgM56D5aDJR9OFN5xp4SGqgX1zoalJQjCaMSfMc
CN+lmV/+4S/xWjt8Nt0mhRe735geCfzpGyUEvIsz1uZgZWKiSSsNv6HsVz6ZPDQV
It4msEk3w7oyIBxgC6twyhszJCtIJnqAVYQ45NCkah9se2a7OCYW8pzIbvVIkEFQ
bbZA3YSMq9vSEoyIbRRUs+7CsrFQSE3hObO0szcm4APjRFHXy2BJwyuRarz5IXr/
qh+HvBiRmGEv9eEmMOFyQY3WG4yRwRttfNO7fbbtRx8n1pX6ovvILpVmT+sLMPqt
m5VTrMxKzGDh6GRlNic8ubhkLL96p0UZSVSGkPgipnMvWcqFyGQjJRc2H1ZI5v1L
YOktq+DO5thzK5weav08496BHk0F34+uRrehV65KR2TT56b0gqo859o+yW8K4127
dZV/INhBR/+kSuaViv5digjmf660Lyz0eZlVgIGgz0eSGKVevbDKsR26eS9Noji5
3wol2re6POxxsxsMZ2fgeSRrNASr7gejIPLB3nuxEYYNYgClyT8Dl4RQi834XhbR
DDjQlywG6vZu8ZpYXb97zAyJVGVO/3IR23aWx6ZF097fsM8Au1g53oqD9S5ze4me
DrCYl/uD3ouKH19CCEdQR2cQjoJ//ioTAxIKdIuuMOILBpbJ8U3vLpMtmP90iGFT
1dNFKBrvKxgz5KbcuJ0UYgAS5bumQj2jusiQX/08BGhogYWa96gUViTtjbagmKAx
SGYWawvaWMMRpJUOBflKdfYff3ExLZZbsgczMgsKJc+SN+IMW5KB4lu82dKNLxfZ
uKPk6c8MWIUVOdtv9VG8ZUJYPZKGjmAtQ3uF4dXP/M0dmyBMKxe2pN+zetoQCTJM
khN3kVf+odmPN8Aq3CY8hW6/C6cNrsewDtNBk3PpVfYWy5PtDZ6IOkl24knourRx
WsaBjtAgS0FAdaUCvGH75rGmnpMJpyHUo1D+QZX3DVwGepb+LoyLOydSO2syA03k
ZI5+wcXToC3SwNtdzHRRUB7fj0wVwS2BLg6+VOxdHhIXkGRM4Vy9s8b430tIgSks
OLHMdn0MUoeZO1pJZMakLocdNk3rXJkOi0EwCMPFiF4kyh9GNbCNZoV8U9P30hoS
fuGp5CfKrzdnMd1++pzGF2/Ws+Rp9aRsO8Egdmr4eU6RGBpdnM0040nzwh9JdZE0
OhuKgprxsBGHIgViymIAp/u1H+zYRwqvKCeMPlWvTL8K6ovPvUOYPyJrcelrkjof
BhsIfemhXNL1d5qfSUf4GqSxhgHqyiu/RrZV4cXOrnCTwByL9mla6z7tk8fOb/TG
Cw+mvpXm+LeekAZHv50pe2d4afGJk8WccBAMaXXiFFla9WYvzh/6WQ7E98RMswhu
WNzq7XF3FE5ru7KBFilcepNA5VNfUQLf80sYwB72MMBQfasxnkmVjxFb+MyTOH9C
t7cEo/yFCOf8QHHNahg7YIXCHtjuMvGznZJbSg0XENyFsOOMn1Q84XBzcCbzVjZg
29KpcfPgOJOv2MbZjDipZxvpdl98BKLzV4gGs9ZdGQEZWdw+o3GxhmwZn8vxqqWa
xCeiZEMbcYqsb2J5n1rWeVvrq7s5FcqfHIT/afEIBUi2TW79YqFj89mJs/1qeMle
lupVWncbiyyHSgiT1FqGyd0RsuYqlBmcYfGPHW3Q2mjKtqohmCPii1vMUzO9voap
GXXR1UEg4/x5Q6J6jXERsm4V4ckwYM/mf1yxmYmV1SjoLk+dzDK/oJhWenJ5qv2F
ynxvvVIzPUHymGfKq/cbuwbpakVQhI2g5nYm+FrXdZwmG1yzwxOL7JZR1M5DrkRk
PWySirUTs8lj9z/j31SPLMaz3T9fb0LHZwaDehdqRp8C3zO1iK+F7UD4uOhL9kdM
4nRpBn+kVG6Fogtdfmt9vJ3j78NKkKFhVrgRtL+2HsXYeOlDFkAleTiOm8b3aVqN
LCvTU4jdbikMTDZQcIHQaeobbyyHqYtjXo94KKpfk16D2EakZISuZyEiWzZZHbiy
6B9TmdGkvvYGKHg0enpfX+VwlYlZkfi9giuEmTpwkDHPthJmGwhDNp1Aqg3wIazE
brNlfgrGNUSZNYRBJ57sS8FEhVn/5K3If2qG+ndiH2wOXZqDl5cZ2sZoWMpFhpqo
nOPIvGpBQC17GvbRzzOwJcr2JemWZZSySJ1oQvz/XUR8GQdkOY5dG3CxAM/DCzVV
KL8/GgVLV7cQlSQ8T3JHS8n90ZMajdaS0EZGQUGznQHTusjC0g5cj93Onhcp4rth
SzqJToC5vObBmlf0iIhqXaTNJ+LuN/WDxsyQDWEXxJmsu+4NRbPszO8BCQ17Qege
9v2cRkFxJ+b6uDp4zV4h0BrfNKDcSgMrJE+aFL5Cj0lago1nn33++TVgHYx1Cw4J
CKCBv1yux9o8znBQ3aqnRo3/NSkAQj0JlLW8sXVS0meZdh00GBLjVeQmBsCQ1Mks
ZihyVw1ufzHtZuJrVXN3B0DccO6F4DHpm9OvPxeODPUbsHtGDOLoBPHhsJ8cVyCc
gqmvpMLE3sNcUD2sY8iPsJbVo3bP+6h5iLcQfRGxgJCalH2K/z7CBJk5C07rmnfy
GmWN+UBGxVh4y5zHZSYZqSp9D0yfFnIkdjFVAGNVX9BNRgmlyI+CJT62Ugd3hZ5j
7JGFrQ42CMs0Pebku4+1luuq7gToUT+BYbBn5IZ8O10/Je58Y9E3HQH8Ms6LhAoq
VAikDDvfvODU/6UEg6f/CWnMl9GNFVKz4NefkTRodv9yBeONmsHYAPOZJ6keyraW
KIX89m6pJQWVlGqUpFmu/9Q4pylkbjdzy+BUtv8n/7ost38xoY9s2PJd1sjfNqZy
r44qXu61fcV/EY+6zKseX2SJx8jr3ZAkjZ5NLLk08Ut0TR9evPHLDicobZCoUciU
56fC1SW/C2MPtROqts5ohVDRqeXDJ95PXLBFUtqOOz1NiNqeluE+b/9BjKe+U/NK
daahxLD6ROU0vOJecmNLVMckoSi/Xmg/DXAdaYz/d0v77Reo1pKBIPpqrVORYBS/
63YSr9BUD+pHBiVDm2tUvE/XZwxgBt/1B4JA5uLbUlAVKoz1BwGxrtJJarIQyWYI
nmifjEnnUI3FJF/rkdrY9bUdRzsJSqR6r8v8QovjxnRuzGp1AIN8HJ8r4YZuplqY
DmGylvqgkNZU4OIGgX3QpAYAfmPta7PcHRL00RXGSkBxx2AvnafZ9V9eKX6ueQ6H
7v/drwq8barfU9p4bEjT831QC0UM1ua8xuYEFeDPct3JiFSKPqhHPf+Bn09pWXgX
Qp3hwawHSOw1TwUB//dehcTJZILqgb8Hp8Mlxee2HFoKer6lsmDUdvYVkoF+xdtZ
akfsjSEciWLsHLBjoi0iOe9qw9uCPR4R2FJ004hZjW8svw2UK3Kjvzz6RvfQ4EuD
9R7G6fYEL1dAAOuMH68t1T4ee5Zwnzz5AlA5jQE2XSXQck37JAxS/FZpR364yDBX
0wzHObplt0RABMYT8WPA+Bl4gG7qD3pG5+IB2k6z9jKryot1oI7CpPcHZhCSIu9i
SBcvdr+q8AzvuceG9ZaH52rD8VqggsqUHQtQwIV1/OnIyaqhxEL0GRuKr5JDJ2i7
P3KF2ev62sgBfuDgeKRkOyVhexPTpaNlHOWVhuKEf13wddQLkR9TDaXS6P0SUPdS
QYXUn3Wcwa1Kg+Ed8mdnTLR7eLYTyvrp5lU8BIeKdCtByHKukvY6lftKz6bhU/33
7DymnhzLXopsZoeAnzJ7J+ViDwJdOf+i45Nol03GYNIlB2DNsTmRklq80Dx3Pq9+
VYfSz31g3cpo/rqdmp+gFTObfzQ4fEwr/5C4zvCTm/F9na275pN6kZtqYwSKljnf
6q4FZ0LaglJQ3X+23y1bPEgifVApsjlASryVqVXDi7JuMOR49pkL4xmjMsZ7eBFY
ZszpJHu/BU1OF4fag/cSJQaUz3OphapWmePk7APphwllrB18T6wxU19lI9QWM5G+
7Lx5ahkBP76AyUGpyK08zt8Weds4f+vyu64eCF2TURwDMBUMVuWbSNMjMQotnC59
wOEJ9NbBh8aOg2lmrDBPLgcM0+51SDl6pLYaO8R6SPtL50JdwOxKT9nXWIhWrmLE
hlzH9CgG/vZRiTw3onACcjX9gPRpwpbtbA/n20WYIXbo+jlLRI9mgYqP6vRY0xwh
r9COD2DnyoWkr7y6Mi6rcVpQyHJQcU2LcKoUpvqDUa4aqLeUbc/X9vWIm8MQ9C9s
MNSw/Y5eCp5TUrqG5QZMWwaxCOHmwKwwHaq/R4QqcUXDOTjatWZjXo+MuP9bUHgO
zgzD73Gaw7EXsLP8ia21C5JyW2BBELNZkwog6Vg7DCwxr8Nu2ku2ZWs1rWExWnjz
Yqj3fIXDwhpPvfVgbpcZCBNtL8eApY3KWo8SoWpdZzaOcteA1PUL1fzM9otF0JcS
hUpLBhTyXykKTPJ5h3GXw1CA6F2PTEWezKY5wqDda5zE5iY6W9vUfwILN6piraMy
UOwQdbcwwOsLqa/KK/97m5F2Px41LcUSRB6WHcfFLqT4aIdn/teC/EsfhDkM6x/Z
GK/m3UvdQGHn0LT3n/cKeYDBUzQbP9uc83szuucjECwGTZ8CX1g814pMwP/aQ6BS
fWMpTr9FP5KmDhltqLotC8jVkbRs1aTZSm3SPw8f/ewE8CHwrgzUt2NJkvCb8gcL
Axvx10grWfFtQerFpDJ3h1xtswGUzBPVn98A61FHXgPrBUf/cL4VzzLiROrvZf1j
xlBsY7xWFGnNvdy+B3WLP5clr2CjDBGiGIGQo2h3USmBpU6CbTDSGS1QTjHFIaKq
2PGKGfClsPNLVXX86yeQaX5fmiuvbsbEfNGMZtUKK6IwGsTDSItfHmYVxvpwtJ7i
8+ISbB86ZrGS1dr22uzAuZkkT3fW1xRHPPTdFq3MJKlQiItDaN/WP/gMcLbI2p4k
if7j4+Gq9z81HAI1HfZxMtTj6NsoiJ6KdWQjuREyK50MxJaYRcHl7k2MSX6F4J5U
ce0M9bkBpsCg32XSk8+54ao/weBVZmzkOq/9aNbDGK8b/tkHndk0sOx4S498YmHs
8m9yj2vXsOUUglxx85FTHD1RDJ3AV1OGaThySL5bqGP2YqD89uRvu9moh+sQGSme
IomHDMDnnZVFAK12JLbhkhY2MZcdHgRB1ylYedmfME4Isjw5WLYLnZlHeAyI1IGx
DafkfjiVMflZjU13uITaBhhyiQxn2g+kZ2tmGIeqVonn/nM7kAalbtFY7eDETV+6
SiGN2Hug1x4fUbtGfY8y6naEmrMsQGmDlljRsjvp1kYEoXYhKDmDVmaOYt9G2PXS
25SUxVEqsqk92WY7iJwdno863kmyJPn+grWY8cUNymQqPc/QVVFJaQgZA/gZ5azO
cT6GKKntSKYB1Z+9QdHnvdzXg96McNxUF6PW4xjYvV54GqnvgRb+hyn4ICmuZPJe
+Hjyoz9+fOOzpcKaza9ZApQ0RC+b66IAN/QgN6KqTrEhHtReqZy7sDkf3a66XtPv
7MBYwk0v4BZJGO6/5QHRGK0Ojj3LpJJ8tMoorXSgmWMrjUIdiBZsq3oKGkUmuRdl
63sHKQCj9C81gS/06/QSIUOEcswe/BP2aFF+eLq2R3X/CvlbtbaB9zd0KrAOGF5f
ph4dG+dJrMGnDXHkFumynT3jBlTCVih+4l3Lc+g98EDy5aVKuMT+L98x07N6tkwe
bEGVsLls1Yp55N+y53KZ7gmTUcSiv40+MoVXaZrDZNbr2/8Asoi3LdQpliCNGC6O
7mRGSWH+FZ7BPIbaEvfBcQ30GARahf0oUV7MN3Kwt864fnm4MWYxC+7ol5lv/8E+
Kdv8hpqrPp6BRX/GGeDC6C6LdzdFmgb77uuISidX9ZBPMU+oQ+oGO4t7QRMDvF+A
TsjxnAs8RPF5O/d9uAuG4onf2wCCWdnZtqD9UOecshB9Kgkou9paythVxX1cADav
N+/ALRFECiCwTGdxokoPpUZHqzkAPBsKnWqwBio4NQHnomB0Hj+ndcBNcTu7j6xr
T2otBcJuITgnPjfV2C53CVk/1tJX12DOa7EnHNsLuNsMIJKGlotgHfrRcMMk5cjx
VUxTowq9FQvBf/ywvvRkhC9RiaZ50UrnwiNtdNH/ks0NwbKIbzQ1N77EkBKwAYgs
v2LIthMvkx+CLsfTCORm9KyoiO3UVJ2g0r8k2ZjQ4wmWkofFEcuI0visi+zRolMZ
CCU2dKqZ6kttbF26R2wiQjWs0BXozqX2rHRE8l4z+jebEdyHKOV6U707qNlyfecT
2bZ2S6f/y0F9jwE+pEQ/jpMwy+XPWAjKbk1JbjQ88QU6Ln3B1G6LlSP3fWRQX83c
1QbkDls+3DS39aRYg6apMNcUoOuZYnRYOXV0t5WFviVwRQ7vpXfGk33VgFw/K3b3
PcXdxMSbeBXoFjvxiwn7kH/qS3KQfFfhC/GKttcGuHWi9rSK9S9FYsJzF/C847EX
mcfZGRvBH60myMPrY0wpG08Jp82Ia8YZvF/DuucIaubxgV+DkJjo03NNI6KpTEI9
iko3KizwLoh6AXoc5x9i5fFgSIqD+WcrnI6agM7QuF/tsvlcozAzHYxN16k1l0+V
XaKJJIlyE9spr/Mf7TNQRCdyeSDAw6fYRroZaPYp+Ojzt8jyPuxVsmO8bAZMAh8j
UJ4c72zFHXSg5kebTF2FPa9hNYujuEIkUsIpaVqMtwgWwPDUBqrLfOG/AtK/dzPC
HV3dhbCLCQ4TOe9scYyKKYfq25tSX1Iwff5zxnUUsv3agDv4xgIeN5R6NrN661bO
KaswFWj7NBECKvUmfCN8vagnjHAz9TKnvUdh241aXF+Ql2dnO2dR3lEeUfAfBotd
505AHgFevlR/kFxMdtbfTCPE/76bCnupHbx6LVYfKooTWUj9WXoNVdWk0dCMm2Xt
jtMuYS8kKIILl2DrjGpJTGXTYV2SLMyKN0arzXkCRdabtXyC1F3uxTT1ZJB1CIRP
f/KrsGH0LeL3fMvzVxQLj5yjozhGpfd9naMVSIHpK+yaYxh1HOvBld92oaGNlgrL
HIQoWnyiJccaOMO/EKe0dhdsXRGBF5znrDQi+CZIaZ8zyLq9Rcyy1kiUShuXeqi0
M8AnXNqpQucNwC1B9Q417BgvpjetKzE+H4n7EUtgpxJl4Oc+4i1BxDu2KIBOU/Cu
8/peqNqMkr+QZeDc43r/71UNcGdhlUaK++LXVB/PvmuQvOURGj0Hr2AJJ8I6HqUV
EUhRenmpy+5j5RPZ2waOziGvLTgrZfzAO3Or84gzRrH6OkR5ohWqGwtlnYXs8/a8
PuCxEiJQEIIX0WC67kln8AFXg2v2dRyTx6jIC2OpIlYkaL+7XystB5yNG3y7PcOF
pRxxyBhDed42CM4OzVpJlYM0bCu/5LU79EjTieV25EU0nQAZ+ZVRjBNDgBRe6EsY
3upIGr4LI2h3iPuKy86N9P5JBkPow0ix9qxTEY5567csL12TDyYR25mbX14mV54S
UW/MVTCb3v1fe46nCbI/NDyZYSLBVutoeua5AgDDHFKCDKUqIhJojAWxQMG3zeYC
XeeEUfptxb5F/0aOlzkY7Rlck2rcK8NyeRE8p/t3rWyVx0MsOwmGnM+X+x893t/g
L4epyLLNkOjAdYb+Ijg/5dTgLgcG7v4Vr117aB06xRzST4oGdiLBLD8oASk3E+2Q
bVijsk9LQbV5m0hSY2p+cEntqJugNdBYfDccmQvZjLDwYqXuXqUT4jAflvMlxT5e
+kXizQPrLbRlroak34NlUL/3T04mftDDr04GqLKJfGeuMPfFoWmQ2pbd/XJ51Orx
k6BUcLtGR7Jp9dTO+PyJ34Db/xKvIpTjKInZ8dEUxwBq+4iGvQ5pRHPI0lYhzWKr
8/+bMmw++6iWfGZ4rs0VnD/eJqvmPYPPGN8B3cW69Toi170vE+2/oVLy2ys1o0mI
Xz7+CIC5/TCGt5q9HVEk/ioICxauXrxyrGBrCPWgQ/xZVRgC+6kqga9P6w5SE98t
4YunPUxnpBSvVSiFq8An/Xvp/cfuL9X1pPMBsXDEywhAfu+/hOyDqu0Fgi6uQfYP
5enNAIxCyty8DeZ0ySdo4cMsjmg3bhSYXCOZIKM1Taxlv3nPymFhfhcKicO6Eq2u
Z6whJ7OIMQgQccjdXFimsfvHMcppC7Z5bXHo9UIwMC1miAzS73uGgm5mXir13ogz
UIFsOeNe/+Jou7I12zjX/AAO36MfPfscYgrcyTh5ExCcNyLKTxvETzfDAXx2QTD6
duHGgmrIgUCdiZgSkJqgOaxrriyJhEykiXjTurXmmypbwClHSDdcA5Bt8Tq0U2oZ
HD5AAbIKeaMkuyrBPHahhRDSbY+pb/d4U3iDFp3V1kXq9n3fDRB5Py7N255/FcCk
uiYtP+ylAdAsS4OqlQrLq08CzkFNb0zlQmYP3kR2jxkaILBG2t1fIPHM8srzzEuV
QA8QLw45CGriwZgcW4t+hEvRZLgOwTfn4Dci5YzoR59n6QOPTNipa3AmOji3cU0n
TQe/x674pFgsN3FrmKmpyAqEYYzUG/LOvFGIEgv/cGBbFIZK/9HQT5TNcCpfTmv2
OeoPL9mECz1R8c050lOGiwgZh475JNZSH2jFiIkyptSNIkNCvkitwzUYRZDSfkTA
UCjeo+3vpSoKnaOt/YiIPz/VOcIGqDPcjj/uET+vquZ0UZjoMZ/itdMkLlFkgDsb
XKMGBo/wAcfJeJ+AoODeC2It8viydppQdhdEb6fKgbfz2tL2GtD6G2VkSUOVigM/
cVewKmq1lEmMYGUJPVeZEcgRkqABJjoWZjxls7i69Hev0uX2iUlO5HsPe3EjljVK
s7q1deJe9STmE0MeGdeVo7hHqC73LLFeMniokAJ2/AHW4GXl3gKKLSSmGAztJsIq
08mJNy2Xh+idse/YinSsml7LKjdZ/PRWJE/xBPHZN2/Q0oAB9NxvMJqujYrQpCez
qsnvMh98hXtnOrUt9l5r7ymt4GYiqCne0D+kmfdUzUmy2QYJ5Ur92QIOu/D9PiMD
XVEpFkWFPfryCiUtRt9nRjqm3o4pZPkBlXNuw793+yQE2mIpxIbyCWHzildiEaFp
/9VIWlTSJhoS579yB0YQqVM4ghz+5tMDKzLs5CbX6e/t0RftjsYOMq79FYtgeFcS
sj/Zmkx8vu0cOXXx/weScBhkHV9qUuWMmzSm1HAmyletxZNDH/cscn01HQALRCTk
/KzO9JhHrt9ds8cUmYTCtAeMWPJN2XoXUSNLERjsdQfIXk0HTxzdlFFU6EhAh8FG
w+RXp1/ThL4g1tr7F1LSZG0Svh5hrhL4MhmcjY1dj99FDzTN9hEp2SQxm0Ciz9E+
ObEszFeaTVaPCwUpJhwNFEDnMIpThKH7QonUgfAiyveW1y1JgnjC5F3EvrmnDSXK
aaUR/bGPYab8ycyGWXKhQu2Ru3iL3kZeKtOLjHT4otm0K+lAHnGpisNZugbKen7Q
JiUhEFb/H3amRiDFGjx+yOwYLSll84dxMRZjyobjMkTDYiM//JtWpRhm5iI7DeYe
ddSajym+KVcRNEdv3XDvM6qWzCcn+1tQrI8/MPMMnpjZWcom/oeDC/Bx8zqo8NTJ
1ATP8HtUar+UdGfvF75/ay8BcwMmw4XOBF+93AhfjW3rzwZXGhNmzoZRKkh4baDC
hR6vzvmHhUAb10Goc7PlbxaxcPZ10hKUX2O2mRTytssIPx2mNFu/FH5vJDmj1PlE
upyGijnXvH586fY/xfdafUSs3BfBZsYiYkhn1aANZ3lulZConYLtjB0IaczYPveb
Vl3j52BomGyMhmg09Bzjzk+EncjrzWeZ4Vu90/4AUcg8es8lhKNWUH+jZR2d76G7
kLme9EWWxOHJ9brcaBXgHzE46PVJ59EtwVWLSm/LvMNRMeQ7vA6ybXRwf2Qgf8Xx
MBYOZRo6S/Z+U/Rtc/6/Yhd4qVEX8V9C9+sFr5S4ldA16r1l4KfBVc/OtOvZO4Pd
Q1LydgI4QjglzMlsDTe2nT8oGjYGwBGCUeF+cngnyRUwJehjnyadN5/qZ+erLtFo
WDKvuEo9BIbt4ELNLWuZoFjh9wF+aO4xU3vfoUnmWaiwz8LMD2F4Jc7hG6MZIjmG
f317zJ+HsyzbYEN9VHZgRm9dG15Ve0m4l2fFCCLY8tAYJ741X2EmO6qPaJ1x8lYO
9TXkkPxRmT87+b64ogET6u/E+DMnkjrjMWfV+6QU8VQJ88rNg4kX15eWNrDrNnIJ
ziDwIliT+o0KVS01yDsmqO4CxY5ojyapOb+r3blSh3zrSzfVyDIR+bBwOev0nX6b
wpD9jdMOTYD6WZruBOHaQpgjzQswfau47k6SJPOBc5kKzn+IlivrpjagyWyi/qmM
Yxb1HkcFpp+AdQ/3J/XoKIKAyCqRLiBFMiMAcp9q2P/zEmEA3H55FyZzbyAoqcJE
t7MlixXnMZCvU3DWjDyqMvWssOBjX6ZGNjqbvhLagDkUEZLd30VnGk1z2v6iUOyr
1p1zTc/JMT7NauPW9uplmmlEWeIpLoAQ3dPbYl7z8DZtOfKpuCq+4w9L8wKYA0a5
JOm/dOsLE82t9v8+jN5PpKDnJ8WFdDj4zH1qZ5ZzRxK83A1UrmR36DO0ZNhKJbBT
EmiIP9uqJsoHknbE+3m6aPX/8roGTu44arRPoGUt3H7T0XM9yti1HI17YdIH8Hwx
SdxanuUA9ekOaezzyMSKLcngwQQZwZ1fPjtZGv5CBTjToismHXF59Qc5bgOu9zvx
Km5wQ2GuL8w4PVwoIQg5760R15qzRS8a9xAqOMIjV56FmVKeAweM6SVBJ5wMMQ7b
f1wkaTDAaebPsQ2CNsQu81gRdNSB8cbazbY8iDoR5yNiSbiUtoN/NdOsSAayYdWO
DEbrmJqBkqv7eyC/xhZg5v9I6wK8icLB1Z47dI49JCXOls0h5m/0WJqY8/zeAI8C
2qyQlPyPQJce4zkOGg6K6ICzaGGNAbvS2a7CQyQNlZMdle5NGiB0h3PrA5gyDRBa
ATmRKivmJJ7Okc/OOW+orBjFEnKRPes4WtceDCLV71ceBcEqYtNEygNQLJ3rhDBh
jZRDjjxdz9WBfa9UllQYU7V+06Em2DZlHtxXXZ7wpbUNPU3eIGR99Y0wyL2RPOrS
YJRMdlbWS495ZMFMxgwHdquEu9UFHtjUIl0bUZZd8dNY58NGabZmSRKWPPX9SEgl
0XmtG/oy1NADZ5w44iIZwiHVup7NUbXY/WCPoDnOIFezvfgmDHoXSrD7AieGQCus
AEk1Q+71YNxLo28/rbUvMD1ie/5azZkbD+6PsdO7rlwwAUF25ij3+owLz/+s/fY+
Yx4DKwUB3EnPZUA65hkjTqlSpdYK28RqNazrxGOrpwdDpUy+bm0PYHDaOk2ilOMw
YB6N+CmLM7eWU1j0yciCuU7fYpMnPB4u5YjiO3NQK8/L4+rCiGUxmq0s7hLkLQ/R
+pBHfAlUHHpFXVpflfj8/JWfO976uydcs4p+09iac5wBHqaXLdwFYJd20/pX12vf
OiMH6Yomanu3KLhQ+J4xtkTfARyRhVb9BWJMJsqDx4nWE46MythChCa9/sN7t5aK
xxBMSw0pNsvXBcV20hj5hnWEhVA97dFEKikXN4R/ddu/tI8LoGvF43KyX/a1yNK3
B6Px3lTyElemRxOMlStACPuc//nTAMrTWaGKFTh/W4zzEfMHDDcqRyC4FUe3+5KL
4gKDVqPATEaTq9gvuc2pGbM79uYuceA9O3f4YXd6yGX/A9pi5aPGfRtjtF96nlqG
3oAx4OfaBKBcKKwRyR/wlDXC7DUp6dkWemuSLW1MNGYEQa8+00K9VPQaWX1i4Bl1
93Bu9Hq22Bk4lNTj1P89r1RwRib/AkHCRno+vNYTSy1nIZjmGbN7yLkCx6I6M+Dq
YoflLdtHr7pT5JLPTmf7BlnNpcCzb8XNx8tFXWO5sXnAJUn9HubVvG4JfmJZmmFC
tkl/RcXsyndUwNlmFPnMBccRrtaySd04kkWRgrQJDEqOXXhaLyc0NmMCeDGK/TkK
Ky/tzS1vEntg5oDA4Zgxs6+hUUTd5NnlPP7G8fHLi0kFSYKFEt+k0nyDOt13pWp4
/27G6BETxQNwa97kyEwFk3KqGucDDbyCT/TaHEhG/dLYbuExxKYOSzvlZVwVKxo0
vyoG2jZqOdPP5k/RiksiYYK5ZSHZtMewOgVLdQ+T9yIi/BhSyLLwsfbsyXgVaMz8
JITQUlG/IYJ7mtQzQaKxt4qrM39EeakyIgmvDrsF2f1poH+dbk6gZu3HyvCj/BF6
1axkcVbQg1BLYATXw3RiBSsmGrnPFfAfhFyD8s0gigl6jD4Xjx2hxZWBBluC0iG3
0q45zRumbM27qCMBQ0i9NhdBeCo+///kC91IJnkTb49hyqSyEgtS+E6vdcJWoBnJ
x5pfJWRQXkdeIopEvUyKyynWQsSL5sNco9DZVM8aM2aOGit30EILwARv1VwQ/aHv
dleZJwIUhSelY6lApDl4ya15XXR3ZJLzkzz9FnB7W1LwlJh97j4be4G1+Feb6mxd
XSfQdySxz2vIzk9eFYWYtOS1RXiJcq378decx1j2sbBYRGCa7NciFkKZZCokaK2n
oQyIchQtmibKczbMOdDef5yykF5QXjyC37yfRDU2Z1x/hTR1yDKeF9aTdTXm3jWq
lfAYtNH0RMiTtTrZRGMODqpL+dmOstpJVWI79AnOGmo8tLrb5G7TNvRhfzt7QN/Q
F4RLMf2IrYORMh7b8tvSQNsPTnAJmmtbIXnRAKkNFvS6y9smbqnjlhOnRJ5lc+Ej
2MgRwolAO9TJLeH/gy2A198lYl9d4/07UOoeDofSMZpvjECGz50vShacoF+DcPzW
qB+eexXckzYlgSe3NLtFUEo6nOM4V4YaTaUqZ0U2OSJtZcsEZHTH7HIbtLOmHBJb
7erF+XCTTSpKqPn2wcCtaxNwLWyY6A3g/27Dk1Ywqd3SIgIWwof/uiWDMszLyx+N
HAaahdlZZLqSTU/57qYzbYw4IrVLp10DJ9rPsoToyp3UmmMEk/4QDCZuyOMDybiy
J11Iq9lBWzWqPS41lr34xP483pH3bbfAuSpMJlK6jiajIUCUa6UIqh5ZwCG4GGnT
7+4VRb4DHNCI6gi8lHnvYAzeT9X16Zh3vGji9g6ozVr6aYz9khkTEUTVpmtRuMT1
DeZbfHOmZtcrQLOBPiXDKJOwJq5CDd21e7jOGYI5FojpWLBlUlBVY4ibKqESKWNF
JZIye5+sqmAPjY7uNhnFjCNT6rRI2VANcIf0XIszHTvnq0sSDf4wT/nN2KGQ/YcL
HQAo8hXO/dcmzcwHLZ9cgA9yQFbRaKaJtQ/rr3ZIEVETfSfgHwxO1YKby7muRImK
wzMTBC/pRkVMeKHU+EkrzddlfbHzstzLnw3Sc+2wq9RyTUuiPMAut6900zLEsMEi
RSLUjDLHb56kxQYDV55hfRd33Upw3hcebLgNJOaTX5P/waZcJ6ovbWyfMZoaLQQ3
Y3j3tOt/yrggFl6ce6SlK5hQ/KclO4a+fsPgkCCvbjtFBI6WBKt4zqNmrEl11tO9
GWq8iBS+OjhND9YQO+kU56HTsZAb4b1PzdLCMASRqOzKZqXURW2fQgMesgT5mOhV
BrgHydh6lUgIaaQGX7PmAReUTGeeAz5SQG7vST8Wf3nkc8mruhOKWI+2CaD8jXie
NM8FJ0pkhNyDRTbsUHzhugm21PF9R/ZhvHzPM9HGoRRLVYRqxLgCBALwZ+XvV93p
apvIdxHVWG4/Tx446mPjfIRmyxYrBW5eHX12QYuw1c/ZyuSyHZplOibeKDptxRHI
bPGcrL47Pf6BYjb/CPstj9d48MXpRUfdyTqkH0CFckdq6CsfG2TL9/+FyDuOB40F
KaD2cRp9p2m6cp+OoTbLU4Qf0sE9KsxCi+fxb0b7Dq98GhCj6VOsQux3qC8M1TeC
ZM7m6GlPFDY4lndMOZu42iP7KBTQBqcWcVS05B4Z8bZtQCv2TVB0UzzweEGh7HGO
HLciB0vSgnSdXD3QadGSp0Yb9PDYx9N13/FH+XrNxugxLkMmN9VRBhYAWl+ORRdv
kLdbG3svF5A1YTboMLpxuUMxVKxHtwaiQ+9RjaBiG5Wk8zW8t6rfqlWmfn8ofA1Z
ksFxG5mnRGESCKlrIBJkyL/bZf4ui77/ON9wS4hZs83a6DvwE50em04jug1zUOjN
4sD3pc7441vIKMmcvbkNFBKQL8uoZcbIiBE5cQapeXcSYn+SPhVpT9h1dhAKLgH+
pNgVMUZEhCH4BNU3tyOUfU0MTcfxc0loev+EyRQUTWgAN38XeiuyoEQqa3oEblSs
0dBknmzjwEvCkCvVFtLcxklJsNKzBU50zD+ZbReJ9/GSJLbg5MqjkS/dXSpGfcvR
60740h8K++ROSUpxM87CQ+zx7ou8+tKtljNPrBzmc8/w6FxZ6xOvDx7AtLBjoqLV
qIgqkL8dSaI8ZGdFe0To0CoYlOmRJ9KszlenNxmVPo5mibXA19ui4O2/k2VCafHz
QVvtG4/PlVkhoKcr7y1Z2KPbGcpaSgm92sn1Q66jua+Wnkbe0iVgVKxoHDSNx26H
OMHoNwaCzPfLS+qQ6tK9CtayMaH1JifyDQi1HindVcmWFe/xUsqRIVqf/KPgeVdk
PIAxTgO5i5d77tKfqMBvl2PvVoYAlhN/ID8WGpIC+tZutuIEBX/xJkCyyrNA0BpZ
V01wQHMZMzfw2SZpDxX/C6UmuxPvoK1reXKxImsal4zeiO+TQjsSiX4mxCTxZpO5
FZR+w0Yem1kEQEu0NmAg5jQJLJ84D1LI2TyUu9O4lEAiUyLlgsUEk7CWy2oHsRm+
nXODGNA19aPIL31QwCmlJQtKeAA9nG81LbNnCgoA6q7X1C4agxp5J1LxzP/wsjke
i7JLYTiDP+5MO0wOIl9uqKUvMo6eJu5Ltf1iciraqsNwwzu/kCG0IBJiX4DfrAd7
SyE+w9SqvLZ6rQRAnLO4pBy0ndzmffgdH05tSNIG9XcTIuJ1MfEBjgN6wQxi7NF+
T0jkmGyxftr2ULLFeLMo4rr2B4cTg/eyJOFOg5uIYT80S3ZNHheV6otIn2SGQJx+
G5Crev9PJ/GskQaBD92HdnbU6aS7eFaVntjLAMy//8Srm8+o6NsOsnKwT8r4CVx2
sSE/H+8kvW3ALQXdKp0YaAkbACtlFOOprAHfcd+4DsYrjy+FCmHAzDw402+qYjQJ
TW6lUY0fE0Fs5FTCLVg7NhFGCOiwSrLRDuDg6pdYk8+VKW/bHXpVUkPf63GVtUSG
os0qiE8M8/sAUmPXUzJyxfD90PdSZi5SKcVgLQwwEnVR6oFSe+YqusR8+/1IVZgE
NkBaaotLiVbHPpFHP3TN5heSOO0aF7LMg3t7ctn8nUPfZ0ovePRzHsc+zk5c46JD
ik4qhyNjDFX3MyVONdR8S3DHPOYBOjYOXkXKUbo17pp1Uc18m4S9qlfzmvDJuJL8
h3Re0T9oAxsToL0+h6GnEwQkO83wcT3jKOEXxcR+G/GG1LTdcAkwPN+bh9VIJVJR
N9Rj4Y0OVYzim/8pE0V9wVXYYUQil+harosp1w5WTDI84yNiS8O/KBNztzsrDuH4
oqqip3kqzmyVPm2939a/lKBTY0cfLXTyHOT01jOh5LVi6JqN+1YWkMjRmNXQ86di
aF0Rr56qhQ1F9Bo/qkbrdlmtv2QBqjHqO+UG50E/fM/n+IM8iY1bS92nsq0nTGC9
HX51DC7C8EPwYtQk4yzaGLuiSoV7R3npACY43FZJP84UlFbtOsK9VQGwAZzdEY+D
XzlZynHGxmKfyzXXZfYgOAmEOS13Zs6MZT8ZjeWTqsQl6C5kqEVjufMC+S43vssP
pq1hvIkiTd9xPOWz+WcoQxDcGkRFs7hRGylq32Jnk1nonIDnNIU2zCF3X8ZY19YA
bvm0XPbR/o33OxZRVACMAQGfqOmhu2tMdZh/GdxaugOYkLDhw9NiQI8j8eG7CpN9
eKk0ANpTNNIroZblNdZdQLwYQJDfdRsqr/f4AQoVk2yhlGuryiXL/XYLPf+9bUAF
9fz+c/N79Stbc20jrtlI2OoJ0MpwvAXr49vCYQ/7q+KyjpJFa3gU5aEDvfzKeHS9
Nu5FswLjaZI/YBHchFAxsgBak76ZSUxKXcmRFhEtO+JyJlHh+/0XwOBy+/GCgkbc
x0GXUqXEh51syM4zFE0xHYT6PTEg5nDSzbWc9eYfFu0Y98AUlw/Er3MzUfEdbIi9
duBASz15uwl9Zcy3qsn44arLlAv8q/Vw2IFbwU2VRiA+yZPAoWBf2G9TK8ryoS5Y
GkZwCefSnr8rn4gTm0o8+ltWYWfFrviBw7A35UFPqoRH7zuk1KJ+im0yp23RQm+w
ZJzAtlzVUpaDHVa/CR9yiLxEihvMRklOSTgfQK8Wegvsm7GZXk/TFbnaPIrMYQcc
wQcfi79eT14AW7csDsStAJa+KZ/n2mrwkqonbQOEiR+Hn+G8nDHwZlFQTbQ3Sz7j
HsjrvW+U7eLuFPJ8gFNmLP9Jrbi6wIcUf4mdk5N1UOywVBItMfc0XbZNXlGy6t9U
PpZX0RRPtAZtWC+oFYI3GvnlNbfqmgMSlIiESWT3cupzhJIdg8Qxsx6QbatbZ8eK
Fz+1dRWKdpfzbTvC+ugnrgTED8P8nbJ7xvtjDdCBEXKiZyCINQ82zKh9FXV8ls79
5lrCQLkZNkfpRF1BvBhYzwg1/DDnmfYHXP9NRtQOcJrJGfboQKgNNptSN5NqGZJc
6+/uYTydXCqea5jYrb8TjvCWPMdQwTBzMyTSu4Hcjtf3aAOeLU8nJkpXjPTbgyyB
M8ho2cUzVFg4FxL8WldzpskAoVrCVvUZjLqh9MRo9kL9cLaKuCx22m5cH3rugtpm
9ROatpB4M/7OmJI5c7V4FKGp1OWF47SlKkx5+3Q0rYPHZrzhnVrrXER9VvHlhhcI
K4IYi4GqrvB12sHbF+gl7kWOYRn8rDkFJS5mdoV6Kk4/jTvakLNiLcwAZ5JVgxLR
KaJzfzOXUTc1CZSipWysqctq0vWHCS0JKporn6H+hGB8lZPqJCYW2cD+5EfTCl1H
yvUg26afNnEr413yC1NIqpmCGe+kZBiQUEVvAU9/yZsjYKljuJhmcSIpyUMJ4nPi
jE8giAR98BrV2BR3sKF2CBkKyqzjc/mL207jDsR3ONlR2jWWEhQmvIa9W+Owjx83
fzCE6BuqFJ65hNDiD5BXGKJBgdbE9bUoglyDZhQT33rtjxJuwDe3flmK7tQgSXoz
kxzekErwzfsey8mFTTbeTLZ5tTzBb1AiWXZOIE/kurXaUVKYyB2x9m7Zj7srBbqy
BmtfS+rzEe0SwpijOQVJeAk60F7KJtNkQeSW7Gx2BpdlZrj+70Axz21npPWIOeDg
GiAmcj/3uYbIWC3QX9fg6XDRHEUcsSjb+jkBpa0i1OL6vqjJgCua1cwu7soor4eP
MRVsTDweuREwAOoyQT67yhcUjsncnUWQvJ9tqNEtXylcNM0/F1GvX0NSDATQ1d/2
rFSBbc9HBD8bRy6AHEfKNusSSrLFiB5FeNxWr5jfWSz4oIeNbgOBS0Ce0kC4ynyB
Ww+wwIap2vNQPQzJrFFNWV0oOaDZNlvc+UJ8qei0QfAlsn0NCmwHto0fX+tUKYcC
ub/liM2kOGq3/1ezKMyeDtUiKwlfahKK3jzYipoTRLkcZmC3oZjZ7NdxBobwHbFE
BmYlOb5mkTXcQb+FECc7sQmEBicNrmBlO60y8CA3JEbf08rbBA+44+hUUijAbIRB
tDx5WgOjz47nM+tUO61OsxPT1cP1GmlNF7xRpzXYZwhHhdsQzIdg2LwGOG1GzhoB
FUrHt2lh4aT2Ciq27wE+W9IdEQ3EGGsTP97ctoPYEuRzozidUgWNVM+eevIHYoiO
EZg3D7wAG4xmuES96nJi6J2zGaesNfxuv6yshV/wBnpq8lT3aa1vNzrafv3k+dwM
Xvq4VB0XJvONZtASL1nx8YifAw87JxvnG/DfvLDywB/JPElB4dlpJ3JG8iss5ac6
cMlXGp2DRhCstfKJvWYXMPpt6LzKCUEoEbBZwdm24O5fa5kaz7JjRxZV2Byt/0KQ
H5RhSynpfNKPkcFqvrQBjWZlyEQGXzAcMphfXOJHqUo1cvrgzP++r+e+gF1AAGJK
3vsiKCUyI9ryfFmaV8q1gqPwl+5k2R2hbO7hYNLHviID4KyPJWZ2W1MMl4AaeJLh
1sKehSyvJqjfUMyQF5d5odCV1uqK5vl7asMop6vVX89+MjKTaGSSqsC2qfr7CyQz
XZHzY7Q3hOk50sn2qR+g9x4FOqNcg7gxDH5fEkrWVjiET54V3zioGYwc2Kiuah2h
zdZHUx1X+sg7XCFx3e1pyMMSNj/PWNjejLjIoIJ58w9moW3PVwjckT7YTFNjfbet
mRx4hEYvArEun7iobfxaUHpV9q2i/khenInTgGlZzKjoFSFnhwLEPst1q5ZaGzI1
smYhMovneG1P8nsJSvQmk8qTD6WpjGQoachAex7b4yaGzMaSkPMSNU0XmOPd/6EE
KcdObm/hfKBiOVAAKIyI9tPIq/s48DvgXS2ksqYUxYU+8Wm9HNKDdI7V3ynAQrT4
Pfn4EcowVqEU/IES6aeCxOHBsqc1S78wQSmqXe//R0Xtv9B+A5GI1l9BY/Ay8DW0
BdLAYlprVPRld4NtJLiRhNx7Nu3XsiVgXt0E6HOZqHXzF5IMKuZVhWVZqm4yPCxk
Soq8k54GwMo2Hr+2RDx3nTrpBPP1MmN/2FBbhrSdRMhoRavqsLA42dd7X9/3N7bM
hu5z7xHg2+wvlmTDZsYYECkDi3RHt4odiXZkuzVeGNMaCiaM1ev9vOcCEvNaji1U
teYfITBmMrPaaEMKh5zvDscxVezypJGyLmutpMHhVn0CkZFMWNPY1d0vDx4qI06A
oNOmE8i4A0eSvrMEUTzr5ISGPQiaLD1i0QIxQIPpOrpYMxRCyGcq8gXjhkTA/AfN
u98OsbiVjc29i0ykwiddYqCOdQI19+P5I/sjzQIJgW20QBrHNhJYnl79PTlxNINc
F8tcaSejaa3yBL+g8Xy5WZgl9vo7Cttj0XeELh2Y1gAxI+uu1iByh6xma3h1qakk
KaxYdaAG8TMFw7mB0jTSFcCeulAYVmi4K1AZqz6Mw1n0gwVWxJIbf9ZBm8gCN/Ar
nTAGASBAclY9LGKEo7+BMZ7bfEkiT9H6JkAEsCqayWnaJcZu4UFo+xpUNtPjx5Dz
4ftVDnVbyE2XHHNZIsolLAhLFTetc3xEmIdJH45dYwTh8TenCWhPPHc2aV/Km0gk
WebkF7ciRsFdASENtFQ5OwP/aTfuMrdeNXMCgTEJk3FYUQ/rHxyawPOtFAIqsdEY
b5QwbpCcQ/Syxu3dNpFaE8Tz6C1MUjYQE4a+zSxWM3L+hhHY/d/868OOjGmhNRhl
twl7ZT+ruU5McdBhoiu2WduOA6mwLUgTsKrBsJmsb2EhGLyUH437jR7JOnkCFaJ6
q+lm3g1kPXQ/Mx28nR8Nu6+2+bOcXCwU6KRpT7SoeV9Icp9KkmDVgBNCKWbP8F7f
MwCv6jaHMInBSkNs3LFWqHRUfcMQpRp1a5Xvt31UBf9pg7jPjSNKOgOfkVvg3erX
2m82wbhCMH7JcOcP0sI0/D3588YmVI8RZNwmzsQeFTJfvqSJoE2C6WktBKyvy1fD
F5jTmGB1AnahOaA4Y811HmJzUegJBnGC7vEJUjTEyKrUYkYxYthghEq1640o3nsX
YWlwm4VKIENNFtHgQKS95r5kME03oBVrRHukUC5kbHSVhAvpiYFls8N7fCskjPs2
uPtovPmz9lD6LjV1svHyxbbwsO+rGaqbN+vOhOCF3LsdJ8zKlsLTsFWpPQXCb/Si
h78UZ6Q8qjLH2rP4U/0CxeBxnvrCAkoelGsvh/4Nxz5N7ELREcWfhbZ1Vo3ZzNTc
cda6rrFVn40RR1C6xn9NpsvcsPD0BDZwbk/5Inp/eOK/m5iuiYljSoSevbHGFPVw
m9ZalH2UKpA5HGUwIUZUciPSrBKTj0YXTe+bORORh5JhlUz4XqLZAPX5TmTc9zls
m2LYDR/bF6P2ma+ttXN9NRqgpoqHo+ViXqGExoPmDDH+7WsYAe7I8gV31hlUAAjh
Yh/eUWwIjzs4f6UKvTm1spTlKt/GlVPVxmVJD2zHuWKqrltWyiTAo+i4kNad2PS1
nLEPtvtxcRH24Z3WJlCB0OtZWIHPs26MPAxBsQ1q7RdZfJMW9nfFwNO6DaLkQqCd
MauK6kMIdkPKsqZDX6t1J2L+9CSTmWBJZlCl+PakAbmN1IcznI59C1KYPubWL/Oq
3gPIc/AfMDsvPldXlJksiN8RlMrW3W3ut2s7TlyX06zZ2f0qlQg4XXSTCVZsHIdL
PY8FJs2N66K2fTI3PzuDepNYDWorP361YN7p99nnwOjKihS3Cyw6n/S7BYqDDwgN
op02J/CjjDfMOD3wxkBqFHHPOJ+HwhSnfnytvE1rh2d+jE51BnQr3mN3fORNz923
rvfOXOqkuxF3ox6mTnbORJJftJ+cw8oQUnTTTTijOMnTrCRJ6OAsZ9e7Q+piG6Vh
357FdyAm4u8NpoZLYrN4S/ob47mKzJcsB4yJoKWIXfmZYnjkIUaiHYPw6rhf8nam
24S/stDd/Y4TiEunybxIMwDRu68wvS8gzzu9yFcuWYGkWmiYK7VNYZe5rv+YcJJX
FEM3+NNWCFTK+bqTMvvmxN+N5ldH8LKXH+h18gLhVWuGJ4atsckwQ1a1vVb0O7MC
RdVCiLuT79yEaceJ/9eA2Ci27lyn1WZqMPz6mqcxh4T0wJZHiNtvRtryg5ltBH5k
9wPo5HhyHajCFzXte46AbvAQKNJ02oiwSY7HyYb2E7lHK/yOlSOOxj2PW5MPZmzV
5U11Jm9RYQiQk8FEt1n+TyolSTCt+pLPZumCo14GyibC+ZUGlANGHQrZX1krPOtC
FDd2cUJ0roysaabjr9QhYor6Qch+efbswo4Ct4XLwSA3Oimxt2oBSpFu8ipUUtbs
QnX2J7FfkA9Z6056tUKHJC3mcB2tN7eEDom1ZZfNtucR2ELKF3ihmhtPA3bifpg6
JSXzKJK+iEq5GToe7rQV0JlgAxlvZydRddk3qx1fpNfiaZODwRRow55fADPzGvmK
V+xSvOL6zUQRaD+mlNRl1s/RYrKcXvan9jtgFuYUBjRAAu8Isu2O6xWkwqOJ99lR
QXAr2J2GrcAoBxWal5yAJWnXGh/y5BUm4bLVzAdMFMCKJOYvZ7VYZkvbTD2hUaqF
cPqUR0qxBwRgwQu1V/nj29VYrFAiMQuf7/OIKaglKLjiODld+X4at0s2tJypvhV+
IGRMC0sWeOvwKxG1hCZpums/px/eHKRMOtizowQYOS10B/yT8mh3CQ8iQdvXrEYG
ZAs8YZFC8P+MfWMaRiaZrt23tgHUu829yDy6HM+F1AkR4PKM9PLm+GZCZc3f9OIU
6vUgxy2TdruCUpUSG4oN9P4s7lEKyZiT1Rrtibo+/pIBifwRGR/atX5ROeokH81r
tDr3QiR1836JSa4327KExT7UURVgKBKjkcBMFcOk5x8hwA0sM/g97v0oR+JRe2M6
Jeq2K5zYLUyjhLgjjCLJjpimq+HflO2zN3/Wfx8ZLWlvceLnmgUexnJTHgiu0Hp+
7wSfStpSGCgqV3M39EILq3aHiZM98pgYX79o8yAk4QTQdCrXAkiuweSK1MgJUmd+
3iOODdLmhg0/6y76j9j2P52Dt8be53VpSoZETlkCujuv6l4R+yrDiN5WLLcV3mu4
HZk/Qa0fTaDyNwCS8mc9P195vaYusJAtEouizMzNd4NgBWSWsjhEa1+VCcP53tRP
kLHoKwR1JyTlUNTtSIIr95fDCsSazDCJNVDcEtRy8m56FmS/GINhQzWCKJxW9L56
RjK1jwT4HY0D66VDNg1FJ+pf5kI/Ty81xk0bbqB26sGZf+bd7VVLrt/OGO77Psgb
umnY5UR5qx3MrGTqtt4Uj95e0L+J6Xea+XrrdrPI0vxuBIw7TKR6YksqhRFSaP4B
KVKYk/WXTeUoA7Gbaj+yFT9mWr+HdcJZ1eaksIZ2fYCx6c8M/O74TNMgh2LCLPgV
s5m6J5N5zATn2JmUMkwQlQl4hbou/yLRSD1vNnbviBy6S+q/4I5FjZ7E1mg4qSAD
JYZPoZ0C1LVTjF43tQTKpsNmvbFXCoFd3VX5MaQA9W8Al8ZWSKppbXDZ9pwK9U93
Yy6B45Y6u/sEgw0vqTc17aFBG8bKjla7oJ6V1yGhjZm448InYZNxtMSGQajlKI7k
1lD162fX+jr6rcCnyrlu6+CHiCUdfS9Y+2+4W8aUN9++D4fjtbRe5u4axbmymWEU
wAkZ9cZa4S7nq4uQEo6iB4bsRDWDRriOS/9lmCNMSH+kyF5jCY2kPxEAjMICr3dX
vWHjHAX2qqtKqhY2Yrt83xQJCGVzo+pmk92KEtxxWox3TtZFLDDhd1r9pvfCH3pu
thdoda9S7wMzqyIRHF5UN87rLpv+86G1bgWDs5n/t40TZXMWOq8y46pe/eEH0iz9
xRB1tmqiHeyJR4FNF2k9GVzZLrT4B5sfczjiwxlvAqWgD8cuWdpZM5hgWngK3t52
T6cztvutn7WbaAbYUhZonVohTHZ2yabQeULdAjqVzWMJBiFabbCMWBZZz/nxskt3
ttaj4rEKeqnr/nJ2r2KhGvo2pKDrlKuDLPZBNcxrs+OUFyAYANw4AJfzMoltgYEA
wezBgTPDgl9sWPakiCBhA3SqGkaqNS98bGGWBDyjIDfcIgGyUsslsyYtoj0IGqi1
BWaqm5MM+DwlZHORf7syswF6mRKBHTI/c0JMxICiRypzo9O2Nk3qfH+conGKmrgs
DIq7QSW9RTiFEyurXrWb89oyuxPKMehfpdZGpgJsegsK/caTrY41MWxjOb0Z3pcK
MrV3zeEFUHIL/YJjH6pWg08ksON8UKo+xvIIjCJ9OEhlkQGTUXjVIboHlARH6LSD
cklTgqEmMh02hsMZM1okIc5tNK5uRfbxtN/4A7yTIRn53GeOXsCQ+oTLxgTutaCR
fAj/JTXUijmZ8NCzHQm7/nJ9ORWIZi3v/vhXvaLjqVziYwTgJMuO44GXRxjgCTXZ
58Kr03i4JIlzGElq7M4RIQyOg0EP0U1iD+C5Qq5tmPw6xr/QU9tDic1zqMfqfr+w
/yhut8TN8mXfwu1flxJ5VOQMihqAxDGFJ5s4WhIM/X30qyYJG1TtIZByyhUOkVB8
X9yuLHcSgDgBqylN+3qC+wgvTkfCnHS0ahZiUv1SxwU+M7/mj+oWRNeaX/gsq76J
w+znNuAVd87zQ+mFngcX1jtCZpL99UmHebBtfFi1JO4jvHkZI08zeT2BvLbqg/yu
TWBBAiX+yrVnp//CBf+1MKvLyVeMB5j7wO8KxLJ8CT2dcbqnl30oHADEguEZm6xm
xC9a5+RRkTRVlEWOFiUuNbsH/9pk3kj2c3V6ZQoIjueXwIdSgMdQuHYuHxTGUn1P
L37E1u+MbLIvBQh6MS8MovhNkF64slh95Ehq+3gbKnbq+ddLjy5b4HfrUhIAsuBo
iNIDDc01j3jp73HYOLVbX1onVydWEzqx4e+322SUfNDlJl/VRyQtdgNsPZugZE/3
/7LiuhGYpiZPnkHgRpj190A2RIpJ7P9Ce8ikg+LS0rqyI0U7VMQHe2WlMaY+xiIs
g2ocAj1kVCXRyKy599Z1v514lE8NomaewHDzRNzPO9gmoLj38q98Fv48ixXQdTsO
257sfRkqZZnGmGk6D09DWcgAi5oveDHYXZYg04oTITUz3lqfOZUL4Z3xV7AjQW3L
wmQOAAw3EI0Bv9sAgU0dLmetGGamKn4D3CF/pnHhbmWjMsVqGbbsdPrqBhfsXkUM
Us9bfw67g6QcjAIMJ5xHfysYAfh1zJ0wKxeMjAHFMsF5MGIj9VO2dM3JNhYC1mhW
Ju1bNQA2GoFRhFGbNDRRg8J3KhTzMEAYrorbPgTFig3epdxbsUhyqvBsgV42lJqq
zu9hfD76A+04P4Ml8x1vsocKbXM0xh+FPPuck9qm34ER5acERTlI63JZnoOptP99
Mo3bQ4XtS4CtCdo0GIpkfHH54ularbwp63R0ANc+p3P/9d4KrJDGTqSNqHfnRXhF
IpGcymKpLln2wCAywRGlOqt5yqFAdbNpgArvSWekLG+2QpzzTFhBU4no3GI6Mzcc
5RmbS9tRdf6qBAfEzbePEyFrm7iy2zkRartPAPcC5uJndkNgayzwUIOItGUniSiC
56wtWwzKRa6ZfVyy6issvvlJaBZxIS9oHmWZi8VWHJAsH4tv8V4NDlI2SurZzxrW
q3Bd+1flCq1aO9BzwpIlq1c4erAabAHg02LnhMxTa+jgZwP4ZvXoilR6WOw1ruNy
Ry85ndcP6rDbUK2xbHFQ10cXwEeQk0vFPmAegKD1Zy0yKaypg6mZ7hz4rQSBtSId
hFtGEXWhEPehNnyPQmcSrjXALoBQ2QmAg4PPvdYB+gPLfzJ4AP+VCRupyUZ77hX/
jt61OEpTGXfi26unNlSFkgbsoUy5dngC7FECVimhfbht2FVZXQZmMMScmXuFhaTK
plhDwtsQDhp3K3qwZB5FZWSw940rbqtlUK8Ih9M0eGJtd9b5N/SaSZClN7q2SzSb
4WfmVIw493t7GehGp2jAA/X84ePx+I1NhkwzIi6ncqaNh6Zff727ZH25eHjc1GDA
xYruMKDeueoa/67GFvNOykKb6BbQyMULLS37z9yL5LG9tgSf9F/dHIFCt/HUZb/3
pVa0K8KW9L9DOG6CH11csq0ixygsSbLKE7/pqSc6ZiuENcFgnbfWwLPPb9PyDeTB
P5IpVQKbgb/tyKY55Pdjwi/OW+yfjYrXuZj5NU3hwHVSvjYGAkFYGz3FBuf8QVbm
gZfi7dxv3qmWoR2q2oLYPA7/PG3q6QXLLR5a/xl9lOef9M/HFgF0R0IV+ngVAoV7
y1NfQwBy2N9LJgXA2797ilyWgtyZJY52f1jcNlD4+crI2fiYn4NNa+RejqPmW7jt
aErBh+FebyGNZ9SR9A9YukPgbL2IBqx1lXbF6hzBlnHdkBLxKXydl6ZEhVcHr1WH
iex2oZlgECNonQnYR3T9KXeveW2ENriS8i3sJKSQYnIHAQz2KWSxcl7k7LezXu5T
TU0H4DO+Dgy2x7qsXHVSTd1zakRg3QBB+vHsn7QYpLGh3/Z/xIYpU2OQih8njtWd
8Iz+g2aJKbywfkVbBEp6ZGmjFLguaVkQja1w+tQ34swbVvHpaGgZLJsfqasVBVFk
WRg/teoWSqy0JNDEMHmDg/W7lLrYMrYbWWJlXrm0JbaRvEFETIsZty9vjVhOFO1e
0EnwFMW+1+Okv6gH3HRII4h5bb8BFQyJHmW+x51TrmvJVq0dKSnmSW33ysgA/puo
rsIjvtZsdJA+6Ml/w+SdAE3L+GcjBM2L62EG104VumvLhA9zyS+x7MNa0kzDio7T
pWQrsEgi62A6y7bQouxk1pKpmEedUyeJvTO8mHCb2Mz2UHthuWPwJLkrJbh+4DKn
Sl7p26YboXwwr/J7ir4cSZesBPLzRzjsMOWHTXi+EUXKBP+spFYqdJyqMhWeuGdt
TvjGAGQmFaLWZQobgGitwCDCBsFlgF1e4lCo3Gjx3oxd19s2qPJMOOn4DuMTT9MX
D/3m2luSXOsthGcqPyqkaeAxT7XtgeJe08p0qNgc1dgoPePQKi5AXSVOvRq9Z2tP
vff1Md133Yooa4oSZVQJV+74vPM7UGh3FM7Z0FuqMTfEc4Q5LTJ+/DxElx2XxmrS
eqpkbqqkTxt4UzU/2zwo6KLx6tI9u+0t6s3Y6IpI3EUCKAtRd0J/vHDbyG5LX8kO
tEIOkpQ3h6uFl6QsEmJEro6xKiZiCU7enfaXmU1NXwz9pSWPlyWC+F9h4URW3fzK
MT+c2Rf5506envgqJizfetnN/qVF8Z60VVoc95ohOSlli9iwig3Q048WrT8XYeg2
90UrKhTr8v8zJknH94heFeP9u4zW0hYNfnB0w5rB2f+2kMkYJvmomASzp1CQogny
gSWN3LftELEgc0dt6s0KyyXqTYitEtDeK8fFlIhpDto1fNPudb7VY8rC2PUiP8jw
JEDV90BkWHfgp+JiUULS8CZeq0KaAWRXXJySIpaUNxU9z5x3f61x3Po/Lt9qhRhp
bUVn4B1j96AQCsPmnd+TCNNwE5VYZnuufxYH1BIinxl7Aa7FLFH0SLTMlTvrZG3z
P0SJHyX49W307d42nPHZzHWaK5Z044idCzvF1nm4S1peOST3X4r5IdH5hw/UWtlT
waqicJhFkdQw50Y/CvqOH5/6ZAEKSmH+/CdTzLFi0SNe6cMl4w2qkQzECdIjW9ud
Kknb7C5v7dpPZUUDvJzoX9BnhCxNvt7f4uGL3XUv63bk9ui8w7K17j38xEF6vhCp
oLczTuZ1/Dn8BHPzDJhs1EuHfQ/bgDVsz5guhkcCqPImUJ+1oUHEnZLY71zCoG7X
1PHuj6wSw7YZh0s3S4udyZbjG+lYddBoccVn1I29nPS32aTNavDU/Gq2RGspARv1
B7veuj9NC0vEEBrRc4vmOQDM1/4uehnO7FN2KvBTpNUUB0RB1bQNErSQ/OOEMWVv
Jnx083gqkUCFyzZFMmeOqhI9uGyI5GkUl9s3Rc1Kz40y9SRU0CPoXHye+u7eBVV3
AUmMcxQh8OzPsRr6uFGeoCJxeQKQMr1QqZC8hStfegKvqBhYciLH35f2rN6xbZoU
a+o6/CQxKRuJ1P/B+CCNYx8Z1UNT06zhbH4p4MFLUgU9mxlx3XLpmy+D0bUD7sG9
h6qt/L6Srh1nIgkEeG+WMCIJ6lxsCCkltazPVxxvk4OZ9+vGwbKK1u/7o7mgduiG
m3KN/V0wpRNULlbDS7bGHck/vkc5F6m+m5RinJLA9XChgM6oI1wzZz0pmpwUw1bf
fnjwTRnx7KF1iBMToy44b83eENoFUGAQ5VZcPX8juaJTNHlg93RZHbVZ6v9IibqF
+/US4AtA0t/4Y4tBHyjgHI+blTz2c0GyvVt+fsW0dcOLHmQ14KUX5shVRLQThdxR
QyecpCbx8cxV5HmVMwSKWnuGChTxd1mCVehWgTaIHKsarbZxtvkf+tGZKZMMmVMv
tdXdQl5mAK7Y2kaCR97XnzrvE0JseWdGKPp38c1NixD81cx8nc2drh21zQSonQsH
CGdP0838zMiXlxnxeA4jzCZzuZeyaMHcEKVdYduzvw8FlV82VxSMaPVF9YA7DKD+
3EWaHr1uPhAl8AzDIy1hK7NDkuDge/Ky8KcgFHyGB4JhCYQEA93K1664PYHrofdE
FiSOFQLGiGozDS2oABzwYiwmdjgWm0XlZBeUSlUQb8dletbZaoleWQcIqL6NYIE9
pJ7yQajELRPEPN7rsqlaSuz+eqYyL//LfQMRQC9oYNZbZFc+bUhQaAx2dR373/+Y
BbxtTQmzdBaRel25QNQg7m2ejz5gWHa52QALfR/VrzfK/m/XNGIeRP2VD8RK99CK
14RU4c3t8BUhOAbGrha13o1GOZ3dBPBgT0cy4jlSXPi9qlkF8aUdDi6rcr4H1mHv
QtdKUHKpvwH3bmQmtUvvSOBOokkXZkogZCeKVAqJkMqQrmb32xcuu5TRrurJWkoM
0DbIiHl1mZYV5BAnGeAnPQd7visCekO34cZZg9yqhF/NM043fXLatG1ObZkQv5BW
h8g5H1zVXiI3waWCWO4rcRYUg0YRjdtDPCrybtkNBcu5xivwt7Ogj0po4lGhzDqs
WbS2aoEbKC928+ki8zlGT+fiV29LSU5074BU7CsNLMyagWDht+YD7x0QzHjWcHZ3
HNab3UQEsrxg3ANGFp56fsFgToxdJ8nNXsdVPc+HhzzuUOb+J7NRerMQ+pN8CIcV
NX9KUs5QzvZ7tjyg3lLFs7jiViS65T8U/a1wSIf34LdO+w/lLoJRmeLD1XY6zwyE
jW1qDptIzz3YNrLZR5KnY5AMTNG4ytQwsbSdKV61v3ZybGyA52kFMYFLdMysNUxT
SvEp1fpgScoyG45Uoiyb5myXr0oQVPQWFCCKtt06EXK8wPKj0wBlmJ3v5XgOC8qR
4z+aFaRDJVJsOpxGXnKBE5Nm7w+CQmRiJqeMJCaqyP/p8VW4o43+GHjEFK0ig+Hq
A9P8lUCLSAZftSm6pDJRJfeVhCe0Hw2cw0olqNUxDLikaDmcPGPpwGaJX9OYCZ36
Wdi1Ekv1ddtJx7+LhcPXOJX5uvI1xETBdkxrvdwmzWwC4ByOc+oSVg3z2LXuPd6X
fqLdKCPZF00gFw3nMAycVFFz2ciDY4iOae/o1DYQvZWDC/bt3eMUWWDm8fWaFhXK
bQCTXLp6vBcNZ3dDtTeSsYmhqE5spZgv/OUevtPu4pymfcjsuAWcyusfeAEgm1/7
yzGgIWyBnxgYKX/GjJBZXa8XSKfUhPtgTByhlQoTcRSbqoFThLEYQnqZFx5H91Us
F3JqYl/T28672VB6nJWjMINlZjf1pkl1Vpy1hhARKtnTP89ngaZMv0efDVllAsSO
KkktzKWu90PqpyZA82ndPdfILzBFk+dfcg7GOqms72APYKNlS0ka1/3ueKnQTgcr
cPoYiWgtOTYYc7wULF/dO5A88Nm5xe2yo4V8e2x31q4i61f9jMmXT5+uhFTqJ0K9
bxlBMzhFjlm614zU0yLbN7O03FkFAeqCTHN+hdd48MY/+JlsnQanjYoV5515Gc1m
KSgAaL/YgmpxlyY4jIHv76LOy1QPsVNFUKNYRtkQdu1RZ34DXx2vbZLmTiqo6ZKX
drukFyoy7cWhnLCQBQZUWcKkf31OOl2K+HgfPAO/3LUMgixFyiMoeEoCgLfsY5/O
FWST89d53tkFLOUU3iNfbaMOEXVQHUqTxAXSbTXzt+rd7KpuhuY3+Ntr1iTW0V7k
8LPveLPdF9fVwlYCUUDXPZFABJJmQQBu2QoI+B4romrdTn9RiztiM3eGveXVAgJa
WeVq5wTeBbE8EfbW2saBQo3/crPZQPYBEi2CBAM6XSELF0VwCBlxnS9mznNeJjdG
crMzeNwOYqYDUYVbUXyPWK7ezm/S+fVqUSUKtCTWLvYhr9g68wOme9DshPmN1bg+
uYMLkcn8poDXLCOOApUY/wkmM1Ajx9IJa+a2ja5Y33ue5f9mzaRKM9j2FVMg0H+S
bAYkP3WdyQUVlEhUFikyHckpC0cCDxlyfyMX18hDx+DeBQtKjLbotI0cEeYhAIod
e4PDRaFJmMna3cOwA3uckiWoA5AkeTG71oTPa/i8c20k24Nxa2E+d2UYSnGcku98
7zGWcJOdHi6l8kRsp/amE6wWJteWDyrjQlDvBWknG18w3+EiuZpKtxHOdZOqU6fz
xzsSHgszFyahdUHuj1IVU0zuojfSMwd9YFXYUX6+j55zlpH5dCxJh0JS5vKSbbHq
+BGEdiKIJsmIugYPdi2imb5GZjdgnCFq0Qbg4dH88VQd0PR9aoL0p6P/x566pdoK
uI+zduiHNpuvXg/CRh1+B79q0UJT+ZIvaArZUcvUTURJRlY1Fyuoedo2824EgPsj
sDpyXv+jq0ngQeUcDpQ7yzimqzKdt2FdvH3wWSWqnRiQdihJLuzuZYHumoRLDKjc
WkZrF/ibEfvnSd+cGtaEGJz6QTgwY7D0MmSBzc29xQjJaw4NMldZaXo6EfXqtoCz
2Iuj5oKy3bhv891eLde6C/oIK2Jn5CtEwMRSy5WdBGR5Eh976oR27ABAkDVS7U2t
PkN4F/BF8qUaAJH33wR269i2Jifs9evFlzZtpQx5Ke6xQA/Qyh18W2NJ7BzJ37eV
csJ/wImp3qPUUJCaOR4GoQrYbcHsq3VARVBD6VLc1BgIhJ8l/04vWwLmjj6KUkiI
zZAhl0ELeWMfSVNS24xt4sQhig04is/NfsP5det+WjGHXia56UsVOVZaouHQqTr8
NsI84gTXPgJwxNSmJFzPZRpoEL68ahOU1pmcRNL8nRa7Lx/XoGlohbFUuZxbVBId
Skfoaq+/R2WqpguQm4hGw/eBNNvJIduQdn45mg9w3loRa2pc+bKbd6JsJmgnc3nM
foeWgkFhY1IaNfWtumh2kmt2iuzy/PRrJ2EiTLkiow8/9hEDolFBpvirkqFtJ8es
UmO8tOG4Z7flJQL2xu+pniZloKwh185RutSvpXFrlJDZqVMN+YvkJS3ts/cAWNgL
YapGEeUamjwxWZnkKns/6K3PQ8yyyQeQ6jx5oNfyjtgbIYK0XV8JrrPQbkFEumN2
7MBYfZtwn3+pUjlXW9KxC162guRQxsEpQI0Echo9t3xUtiYRMP4ps+kPaiBALvXZ
7MEBKNEqCXKbmOfdb6Mode8/YggK+khrCzhD+NS02RYVFtuUD8ARmFVVmsKtmUiJ
0lEfyZmZKIasNAFUdqFOoruAojl8iyFtEMdK9Hsm6gaMpgs36gAvvM4FvNnFsge1
dgZf99cSUfu4mbpTe7mj1t3qJv482s8hxUfkIyJbJX5w3SC3YS1m6cgz+0t1xFhM
9gGRca/F68Wl0eAM0YN+fCf477OfAmWjEl4FOIUZde7mJyT2KKdl9zKJo7JXEbDe
0M6fX2NTWkUPssLh7m8t5TvZ4CwYvvddThtFFiIJ5U4CgJR5BhVuMg7BM7ZW2PjL
Ag9zFwnDnvRVlabC61alOp3rK/iMAfRRR+FB8Mb23+1Khj/sFmNBBSxsTA04d0MX
FU6W+fGCrPgwczUf3oWISnVGlzQc8Ijrj8YjzkW+2mAHMrOhjfS8oNLo2wCH8Yjo
RwDW2TYaH4Zbaj90QuHH/VnE42u2ljzqyr3VhnSsUweDBqQCBofVpCv6aVGRgMbl
bfTZx8sZQb4rVnoq59xmfAHTKCKll0grmMhLdknR3/ogf4pKOfQA9kC/m1fKwOnX
+bjFSV22tncg4Tz9T1CyA2ias5YHMq+/oSvhuH1l2perWeAFhm4jF4vmM71TgrTS
NNX0yQBvu3MHUCX34ON8puskXUbGR0g6JSZLdDIPa5+/vpE+kMX792jagZBfmcT/
LXjcmYeDJ+e8X6ySdNfqYgZPQALinz9IlTtOcTEjbGneaQnYSYY9/1L5mJHeqIaV
pEOrx6liOvVg3hdCe7aeKPjTR42boXHr5k7LqdE00E0yrgmtDur+e9i/LDKqGYHY
Ubt8ZaRt1/4/mTMHc1TaXW5yJnk+javLoK3fdvfgCKRklXqkbot6lQy/FeBfduRG
gxkE3wZjysGLSrv3GVMhP23Tetcsq289RPmd8V9naDAmywFs/1yo3dSHx47M3iAZ
MbSSmneeY6sJllQIgmZDmZKsL4j86IScmSux9B7im2rsBqHHGDMgGUuD7D6lZ3UO
0uQm9LO4/XuT2P+gcl3aLKGnGf/SRRLsQXqd/waxAPzUax7L3kRivM8ukpz6xKb6
CXIHnAziO+miUwxmwHv6EHODsPguQyACvase2VxpFY24NBBNHvBALNwoJuPTWr7V
F7Z8JfaSWi7w5M4bYfuN/QS2S5dqaBDJaSB2HhVDgIxsK2OetAdN18+O3S+2Sokb
thFt2JJ7JyER6UEAw6oQwe8tqsDjxAb8SagjM+EFexxEo3D93t40/S9fSM8cSPO8
dBrzke5ubYeA1B4/zpzeyZ/3rMl8pdeQd7bsbfrbBXRpI6oK2QT9g4kkz6vkKl6A
P96iA1ym7jQV1dhnoE7lWhd5/rngMsOuvH7Dy93gFhLYshp48KcJw7uja/AgnP9T
aSCv71E1TxwFbXPz7hInuwkqGSaWTb3ZkRQfltK2hsvyDMDWQkJ67tyRuExcR1xg
3TLDl6gQwnBG5XL8YF3Vl9Kapr4fN5g1sYBa8+uXci4wNFw7lL3Wk/ZWE9jHelCD
0dFp3oKPo2Nnle5CHyiFdkFL3WBCbow2r9cva6954YioKdYhbTSHcxKiCbnFkWvU
rsRG077C3CIUFigKrf/jD82LnmRm4lQBV7rmgKbTfCrWWjq9n2WbNE/Ry2T0AeUC
ND3+cSEWLPtWf3f6clWgvO6ytrS4J4DYz4BXM8GHMfO8cgstaV3oDoA9pqauY0sN
zFsXxB6dBR44q9To4P68DMnV58a5pKbTh/V2EDaXxCd2c5VX7oOXpRhv58DSXm3h
MFuiGuduR8KE+gwQbQWWxLi+t0JK+Rolfa+Btr/axe2c2Is3j2VOe8nfcQILRwGx
hCIAiYTCTBVmwLpxBwvFEhhbeJplGZaMNmb4zRGg61N7q5mVzUtyS5ZjVrdeZPNK
BqIRbJB52vQC9c/vscnyYM7mr4W0cyfnR2D1W+1M+kA6vCVic8Kj1CGhbNJ5ICak
n4cVLEq/qpa4FZ2l+hMbS4x52YLNNvjVh7cFCaZ2xg07CueKIRR8Tf+gC+0GGCmp
N0jYn/UpCBa3NZdNrk7nnEmBl7hhDmiuhPYGa+0UnSgoG6GJwPai6qx/R3b+GpF5
jRp2Du4bGA84CVoq0gRHXN9biu7SZaWlrgIHoINBp5eOmke2wuxpC4tfFaErRZb2
mZsCVz77xl+xQ/vO3kIfT50KxqHQZbtrMkpbbbba23MIlRkwvYyoDmXTLNiVXuzz
d1yYDSvlpWB/xPXrkYOjfJEitdsRCKOH4NjE+3KPI5UoVQCIYI6HGyro1YBFfCEv
XpclmBZ8qaAQAzmY5alntvGT+CT0yosBFD+MuXbSg/V74Fk+k0D8WjuFhNn4Lmle
KNpiKtxlGRLlFIQGP5saPlf7AfJ8FDR4/9cVuL+SGtcDYlCp7y9xBjAKSJFWTQaC
1tN2iVd5VYXuw6+qg7eJ44c8Mk/YsvGKlwWg7jV7v43EeG1hT+MhRSXTTknLYIPP
qopwq2PKrlvuGG8ZO+/PG7YBH9Ie766H1TSef1VpSbfW3jsrjvebnV09mQIeexWm
xFA1L9EhXytlfQLQtPAyjFglVOjhrLoq66M0VOaQMO8akcIVb0UpQq+Ya+2fkUpd
YBfFk3xDbXC4UVty0QPUZKczlLkDReZEP/O4HvBHgQxaXONfhn7JH7UGnqxbsv2Y
vj5/GDUqhZtrgvmc0zMmFIx8lMMUrHsXQ/bIk/gaKF79JcECrMgAwtG3RCtTzhXX
xzNpdpZk8MYny9WF+exkGKqp6sDpeEre4978MlluGFWow/tce7Zc4tKRzN2v/hqm
t/6n03/rfXDRRLDH7QTZigKRlewEeiWIRrJOlpIwWmNGSzABBTT2XlSaZKX78d3f
SestwPurJjd1gY5tdbMJHWgYB/xO1iHQAE7CxMIuHJPvAfoy5yVNWPRJ1pqcD+Wn
inmTMa0HN68rfVX2Sy/81ruIrnLv7LLl5s3JqvIm45GHplBz9fC99OlZlWaMRu8g
pK2rv1oPUg7dgdiMEXTuaXslo/7tpGWhLD9oGGWZNaeE9HyyqYYp2pL0xx9ecw5b
AWdsrZ45ZF7OK6VqZ3mT7hYtS7t3XXqT26YikoOhUdftNm5e8VHek2El6jwOw59p
x2lqL7kQfLPpSMhRP73pKCtFuoXi7SHjNbA9bgnKUVVyjVTbUyZzN6khthdkevbW
vPL8URZu120vXyQJGLmJ1FQ/RhMhgYPidGkgdEt9rsbu6ij6YX9bICbHXho/rsxK
IA9DslYRizmqKqgHTPMPHRZcuxyWYe/8CneusbqWL5YHdtxK3IErYKn8noggot+9
UspWo7EUwDuKMfs6x5k56LwAtNXL8Fp5s0dPzVoS7cg05KSsMxE/0ErfeFvd8sTH
bnLzKIGUcpQ2MhNIbfcMqiDoB4PfILW3EUcU0Hz4xv2jhCs9AZ5yFt2xjvWQ8hHy
NjljU3NDE4DyVA6NYY000mh0K8pD6OO40fQDOTqJ/QrkpiG1n+Ls3KcrhwtlPRZS
0QU2vzXD+8dh4DLtpDEoowWNFvM+AZgfCX/2JrrcPruzJriqMsmlIdCxG16DgwIB
MT4AWvUNnmRRnMZOEbFpD+rhaLpwNDDdDTUHlLBkH6obIjRj2B2w23kVBi/6RzgZ
VJTf3zpVM4Aa9y1rR9Rp+v68CJ0qlb6D5LKAtsGPx8gfx5nY9SP56ktLxdPO3zT0
GuNMhlRjrnAd6Vy0ZAQRTZEVrAZh8mjq9F4PcMC84GRMFjh+QPHuRLXwdKoPgLX+
Tn/3+Smo3cXqo8zxkzSjUlCaOjN3W7DOAW6HagpHAu0Smhc/a7DXCpPYT8Sp+98s
puxRyRY8frqqA92nWuJC+YGi2oljF3QhwRpzIt83I1SAeyxh3hI6EZUDM1OBQ73n
+d73lqOK33wqt8ITuOH9WB8CeD6w2Pvx7aAVQ5Ul1aN6e6ca3aEprpSEpzqX9zPR
GYdHWG/FHBA8+4Fm9Pu8g8F983nJZQ5uhYvMvu+/2u57cortwvU1OT0xh+SpsvdD
sFxtxfgGO3OBeh0QRlp19LJwP7dS8PgfGRFlY9tH+Wnrjnl3pyUW3/+fNpawj/fU
IhPDyvrkf5AlyE0F9h0u3nCbk0awL+OL2TB9Doyp8EDeJbWJISSH7BHJLKu5NNyy
8eXySWVcjqIshe36PSl0/LlonwUaX2YAnS3w3kCjPi3D67Mu6L1IjeI79u11oXae
QsBnMdtxCATaGVZFuuLrNTYKqk0fvehC4QPlxzXvGX3gv2Va2DknXZoWagpK6WR4
m8ufRAEwXFh4wmE2fHiOB/fsslnfRZBSYJR/qZUKm/aPzZoBBCKrUSPdhTfUnMqN
zhzSnzPQk8ND+2p8yfNocLmM2DfxWG3JMORiuT/Ep8WglMKKPOcUvL5QcJmwXCHt
b0NvEP/UczKDNZnIRlnCZac60G2CieMAkiqhVTJhZrqi78tjvYHC++8ickqpVRDw
xASaFyu4hmXrN0DbseYQhH64RtK3CvlDwo0bprfk2EXsvyUopVE1FKUe0rs90pLR
W7bwQTlJqxV+T6eEPHBXmUSJMwN0AKMgOgn/mXYtsZ6mk52gGfwLTExZDoJPTOdC
FvzPgb7WsdlmYflqyAqIEwKVyICYIzhDJAX4aWheTBZhv0udPc7wZrDN1K4w9dnL
z5AgpSec1y0Zsd3BzHgCwelzDlyydUzOTE1JxMwI39g2nS8jxBTM3IWfsU5A98cP
Of/c5vq3miyEM4ZlqMBv38VKnmUKPpMIDpu8UubRbDx0az0H6AlTPLVd22EqjWGk
RAiAkOLiNFYWpZHxODbkeR2DmlglPyH0SYRuyGVEt5gDzEEOhFTl69SssTexcUJO
3wIbWZGiKCRumm/OZHmnCMMG8eW+IRV4aAeXRRKnjaz+COfbD7TEb+xPq6xl5Iav
GiM6kAysMkDqq3aziUq9ddVgNafkuLsPia5g49oKH8CTSOuaeTBn4+PZyd2/Go+A
nojMdcW61wTXa/CeeuCipo3HfT0+0r0rvlNBFVLffFksPR4gRrLzXb0mVLmqdmbm
+P6HIS+3kzPHHRI40TT1D5oVdike8t5ruHFfqTCLFYO+wLmcUx5UZGfaMs93WlqP
q0S0FlewlmZWbWoUN7SGI/v4bP/O7vEkJ/uEyyuKcCp4U72+H4ImHWfPW2+VI+JN
BYz2WuegLLu4LADXEK/uPYfduGoRRNA2hPcJF0bCHRakB6zgr1ZBlQ9SakXFUaco
MUWeh4rDBDW1vhfaYjRWzi8n0DOZpAZf3BVEVuffdbtp7pDyZtoYz4b4quMlY/C3
qnNcaJP0tHyKtLgq4UFdAXGg4Mp/aBpDZJTlJ3q4HSwHC4o2FZ6orwIXJzjNA2EZ
5ZgIvuwW291jQl/nBoHSGI8XIIMz/DB0Tgsr3zPA997c8e9ayhP4RxDKMWXzLE5F
RJTtRCPuOvFx2bjFMbYpoDPcL4pyXT7csqYKzPD8b6KblKLHPQ+paeeG/uMM098q
Y+H3OKJ8I/OGR/wvshheqwkM/+DRpX6+WyUz4mPXLmcWIFnZKZaq+xnxxiP0dWc8
5coJ0wqWehAmsL8PxNOaMA3kEp0qYUrKtyVfZxyk7yhQUj+W/l29DgZ0neZ0khX/
AXUKpk8Z4TnXgT9o4UYxdofNQ8l8CcUGxexcj93zJNA4jKvk8pwYTag8ebsulmoK
MQ26yfN/JGnaGD8vvRURowxoHk4hriEWqnD/I3ynMzlEqbyg8iMyceamtUoUCh9W
o+Q+Da7KlqU44lv8ntkQZpDgBWwfHk444jpxZtP355rqKFUVQAhQ6DSVZ4WCDP4M
1FSevUqZqPebVwByJ+BaEWaAPjy54bjkg8MesnM3DKqHmIxAIZy5RRqtp9jR82Y0
435At59cUENjCeQEhPXf0wnZs408uWa2xNuRRrpJdEcaMxKO7PeT9bSb44s8VefN
ecEMsQM0NPXhpcOhQGMaZ+/bGvXF8pIkGjJrjfAWy2PrBz4oj6ntkYpo6NgzQI/e
sJdu87XYdwrQMeSosCIlXDfiVyV70tyEiiOBvUwhH8XGZ5iEAUwotLrCKYjygpFR
n3cHeXHMCxgkD1g89lRquN2tUtsy1rqeo5476BE2VizLABOErfVuKMXDlsLN3m1O
ibJT6UKVZnTujR4ekf33C617fZGYwudCtBxq7qk0h21cAIsty0pB/hp4bjurcsKM
9+UCANcBJtjTY5N0A6ps6aDPRKvy9ZJVRRpdb4BjYgQ5JHXbOBOz1S4ndHNI/fc+
tMOUP1Zzzq9AjBDXcloa+JRPAro2GJgFjnsEhiX31ZN0ZJXtpeaFH7Lnad9AbIPP
GNsPH0Raa0nx0Eu5cGC0nMLCg7tm/b81cgbr/uPGR9IJbg1n2eaRSDhhuK/fhz32
1dZy7mfWHr1RFD494LH2/kGEggCVn9lDb+wE5mATJkbE8OBwXLYdPvIEG571KynC
1RWJev0oFMs05dahxIIL9TRx5XYO9SQfAi2IZBwCoEJtuGzCaawOARcTPowiDQ4S
pxcfG2cw7LSVPrvtD4RoLu3hfXMjj9XA7UTRYm83a3rFyDvle6FxBEEptwhEzS5m
R7FDS/XcihBzudWKoGOXvYOhrqz3ygM/j6qv2b4y69cL35/A/lpBoLZ1cggbXl5P
Y/VNgxJW1lI8JRq3oMkP7LiJ2Xg6nW+oEaVy4cIuAWFIlkIv1VLUoyJkPA6AWgyG
iRbmJlRi94YrFYTtPNhGJXietdnXtRsxKsPhqRfgDOV3izYiRfwq6Ic4CIlnM3Xd
MXxGJX2DOY9QzDPc/CQk0PknPqgh10puITdk+uS8IIrAVkhG9DDGgZrLh0T+37uW
4uGAoKjHfZ/XZqpb+HGrMAPfhJcfQUXLDjv5QM47fntDDQC2KSiTjaBTMMd4IMkc
xROJ2DvdRQm2Wfr+I4GtfS5FBki6ujsNFWH4zv287H6Y4exO7gpIwwswI1uZTGSN
yn+ObvuypFyC0LuGaKSPFrDt3x1ULLBKJWN8+/M3wJ/GA1QVl/D4Wb8kh5gAcZgJ
Mg4P8fD8QBSC7gW7YYSD6i9wQYiOP2o8zGTdKzt3aBR/bDaVYI4TLePSjUlq4Rla
heM5TGJAkbCidgmEopeQcuyPKbC6tryNa6YJODDqnS7eN3apgqj3EpOwiov7BW/B
mz8qemKNDOOEgPawH6eBmHChO+XBBsAsJ4CNclEzE22wpf31lU/Vr4g/KDjmXMp6
Amy0uGcvPBXZiCvRATyUUqfCn7RPC0BQnraLtlzEtQ0T6aLzwj1KdxhjY1oI/9BE
g48PscOKgtKcUnQgsRmtJW9bBSAbY0uf8SimXsCbsR5AsFwpaZtaMF1TPuh/gugW
qgZ/iACeZcGTVKaNODkIHsYlQ674Vxt+xcGoGYUEtDODZAvuzRJVsAynoUxP+NRz
pOrgLFfYCLySflyx54niM2aoOV7Aw67b2XOLa5fkbx7/WpBc4Yizhq28qDx5kUrT
rIuAA7ucUH+nIHSaxEC3ZFEB5UXf+qf2vfi7Jczh4AVGaV8sXV15sW+peWrE62MN
lO2+cY/wvN0GXfA+Rzg6pwVe6gxT2G5CCZuk+N25LjH8jtGwYu0klxV4QrXuUIJK
Os0YdSLahunCrDtE+huDcUBvEFumExUH6UptuC2Me2hySzMVc46U22ZiT0+PoyNC
rB6L7B6gEKFyS9HJjx7XzPQI5mlGJ/5aoWcCZugz9nELQu+zI48Xa54DjY3S1YCg
CNywoh+Rq0Sriq2WIURachFOQ5scehb+7o6Bt6ezNtcexLuwfYjRboTK5uVDYHVf
3urRExeitwb//9prr5fmDf7E1j3eZt90gqpbPOr0vjM9P3NZj+cSHG41AbXxlsvu
Yl8Up9yQ7/ZJ+sZsov3VWZLYzp2JeplBEpSW+Yo+27rxN0qcz3gR5rLSjZcVzyJf
pZySgpquhdLSxc+Vj+02hL4kflSNHMlY5Jli1dBZf5DQkS9b4bCAzF88NzzwnSgq
2NsBeD1g9aBELlNlA9rvrNhAd0z1loHzySIIBIWWQg+UrUucEHQgw/5oXlL0Al3z
U9foxwq+NDIkYlUv+7e5n9EkLK8uajCrJIg43T+UIC39zARHZ1mGIup5uwCALaLn
5q7Z5FL2vbIp9LV5mwaFQfk0qThpiJDvEb6v4aogrjkZtL318PyB7vfXSKiwKQK8
TLcYnNOuXdnMc9hqmvrX5xO9vn5Sr/Uw0bnXUo+fWE8PXLjdlgd8Ei3ZnlVHroWn
PVcKBRbrLZ37rqP6Nmm6td+cjX00lUydG3J28/YodNJI2+ES19yvml3fm6SEUs28
ix1vyI0RrArFck+F9A8j1BEOXQXxpiYb8CUSZ1k0D+wCTLaqfPV9twlBTOBQ0jNl
uP2XHvY9qDbJ7QhazjU0DMorDle6Vjb7GNduY3DF6VUCvwCyk9PkG4+9mJ5rEQBQ
FZun1Y+8lYZQwiiffqV1XnN1kyGADahJiJOk3XVU8SEB4KSHQjAj7uC4PAR7wiYp
gQLOdYp9gD1K4a7GSM0oggDxTYGNQCJYUMPvMAjMTchbPwNdLT7lPYmt/eRrddV9
lCyknKbTe3TimHXDdD/lVsgQpyHe8J1bbkYP6D0vvVveW07PXtQAgXHWeDN+Hv75
MbPFk+DYyCuw21azcn9z6J6WM8Md60Hj1nBDZN7Zx+Wo38eOsbmQ1E6Z40RMK9Po
CtbwoqThKwvtxDZ7PpIIX6O+bYvfWJ1S56JVCcV8j3E8rg4WUe+MylQ791TiJN9V
M4sFwm82uOTxzG9RIPQpTAmpoDNv7ENunDlWfzbY+MfcIPDYtxXyJxfB/vfZ4W52
MqDbd44ifkkS0QTwG6guTymsD3JE5PPijuVBhfHStSOB2RDQsUJxcW2Lz0R24M9U
+LAd7eG6gWDzR2qeaDUII7yvRnHKF9+Dd41jGucg9thGgDQ2eUMe5mZFgaEGa4BC
pOrm84ySJIIFKCeMiB8/8Ql0Rlv+EteFff21rUB+7EwLhIJ2559982UDxaSERkS2
df1dFex0H+9D6TJJenJqmhWxr0EtyZGpWEnNPjN/fe5vqX12cCOPWzTP3CrVb0BW
YiuEoIFBGjyqYbsaiVtF5tf9Dl0jDhUhjm8oTH/JJBKP18WIyjvLz9RZVsXJ2PTR
EmM7VcH5IgnJr3joR4sWq+GaeLmsdOAwrdf59scfFlEjjc0S+icthRKOUZPhuMR3
oTV4NhTI6Dk2ApVSUMuAlSrEqymYuUsnL1whgMqORD+dOh6/8SsjW8xcwnOjkx33
tbUVvdh/dYsnnCXlfhm+3b3y85Zl0YXlUPb2m762omt4bJ3BiR+zrgFnP6HhW1Oj
Pkfqs0JjXEUi5F47Syp8hflKASpxYMm7cTEz14rAHmOJ9+dfJCUKR0Rf6PJ7Lydt
kBN+hPUbBZPQJqk8O+Y3NUoZmcL921Qv2oTlS1xS0XES3c/gGV4uu1Ol/A7uv4Kf
XWPkfJfziB5r3qRDn038Yydi7LBapTbG8nJ0yGvkzfnAFITqTFG3OaGfRGfDxOWb
tAcA3R/I8w7M0DqERxEMCITLwcdPGaEzRf8IDX7OKTylhjyLRjRkVC6KbbjtGyvp
eVnOCs+ftEJN062rVmFGDurdfDDOQcb/ZROvQ4RROdN6oIivEYmznUzb6Vuv9G91
+zQHlB2cnvhaBSx/81eq+3JalIM43gZBy6HMFtFy2IzijF81hyKCl0puIdLsA9Vl
E4fxjSzsRoWjuaUfSn+GlV5X1OTDvPtAUm9RfUNwaea02KFip6QsqhztaTdkUUeu
tXCAKy0s693PdguN1XzCjeYRr6Jxb/TuNXKxPvibcsddbKx9wdddXopMNDfwKXKW
mjgo3MlZ81+MdiKOcswzvpc4dWaOy2qYQPS/zliznfxlIpOrx3Lt7vEUphMi1Nbm
iRexMWEEAg/M5ZFbNpw8iBPWB7erF9h3JhP6S5VvrSe7xdNznLlweSsSmN8uYkWq
kESIf6rupq6YZ74tZ6EVRpBSJaiI1qlq4hHDx7OCEbT31Iw8wOmWL5R1yzL0/KJT
6p0bP05WY0xB/r4BHS/2qQDg1O1/cB5x56h/j+nhT700HTxRaoVQ6fPuj3p61sfy
+A5wF4dRXnCOpTZZtp2XcOjiTdoPxDsxoJ818xKkxhvkoZcnkP10Zmv1ueYCw3Gf
SMk3FCBLcDXW5rwz/bOhxSL+I7QsYtsd5bpzvn8EMDbaOCFLzQm1eAAjlv+RpkZR
uLyNCFVs2B2tHM0ROB+fdWn+w6pKJInguXoX1kNihZhIkTGdMyg4mpQphZw/H7j6
DPD1XD8BAjjT8UbP5NFPXjviy9MzUCkKxmGN3AgUtwSl9crW/hiJxhqURqVSdyFg
WNOWNRutDwHV4nbizV3upAfc7LJWckjxVIQ2MzIVY78A0JFgz0DaWjLr42nc++0E
/YTcqF95EZW//dgYybvFji5SXsWH+vBerxdW4sRLyq/6GZqAIfp1scdn6SdkLPdy
G+Kfb8SfSEqoTjz7pCZaNgJRuE5U0LzesxIvgzKYiH0Tk5d+H3DYajINc1r6lbHT
WswLqIy8l5GAazCaS/jrq6ZtQQmth+OLoSgCctGoccgssbgp6za2wZ36w7WLdllq
SJkIOBUK8NT2CNSno99VYbTCf7BvV0WsJtLDXCFl8FHX1bEceiJXszVpWkLTt4dl
UIlBsmeZF/yxCAsmpV/2XMzQ7WvfQk2v2RD1WbRJztnBQHajCmWtC5EnM+HOHl+j
ZPYIuzrofYh/WPudwMTC0MeUbgJhGIFkfNlz9hJI276wbquhTnOcILP7R7/2KteW
Ad1EMvrLgc96zQ+cpYwfKFWwbmCVT0yYSnjRclhRFQr9GfCFznv3CNx/r0/cy+dV
QAeSkoQYVMyx5CUmWPdYg7pLDFZBSh0mUrFz8qsxQNZdHJLq8PQaPtWDJ4Bf9Q+Q
EYUWlMm1LsFhwWV7RgpQfg3rh25WMnZ4+mPfRXbX94+JKvQsrCO2K865BzD9pzh6
Ng3pQVbV7bwe+SXpHWCiTmu2P8dDXcui6tMYktIE9Wt5QnIrYGnpCUSlVRvclTat
fia5JoQY5y4cQGk7+Y96DrBHUhllMobXkSRqaXHsMKdRRw3kgSbPX4eEKCXA78nN
ROKc6IFtGFkZ5diW0yoWVHeqWBdNPb1WjRZ8JoyxSaxlCkxFBjx0hiaNoszO0qvT
dDwlRjJysX1KYe7ZstcIu7Z82TKc4IiUjGb/F2q8pjKwe6Nx1ULpcErmapooJ3rO
Vh67Itz1l+GcYHkz75gf2akueKOi2TnfuZcKnw912+nfIP2oj2DCBXFukiMvx0pr
ULmgmvaVpSyYY8oh9MqlP/+Xg1FoY6QREw0Dlb8EmWYYzAZje5p/V3xJ61U6T7NM
C9T46oocx0oEGOgb/yYOQpFRE5d9oKye1Z5amhUKfPz1/4Tz4n10rcdccesBeHt1
TGxIMcNNuFRw2SUipfe7arEpCgdb5xsy/DCMj6pYB4ppmmObVmMjCc8LWVoDKDqG
DdW5pewQ8Z7ymTN9we6jTF7IcFA7joi/i8EIfeb7D6xta2/2yYri0hHMGePHV+Zv
HMGCnuTho0fNZrEj6ZlCL3JFthH0cCfy77CV0VKfn9xVfF77gj88grywcgayvxTn
Q0Ynp7go9X33jBkKWdqNkh0MEddHmaeXE3TgJsfZHJcvoCiu3lodF8uxK/ywH+UQ
2lEalwia3zR3+chMJSt6jS6DpK8HoG1XbrkMilhKxPSTQ1JqS14fiWuS9nJxWdCC
GNyM4rwTLnJh44S+vF1i9tReH5mu2zFPjOHivRaeYPcWeEXPgdLbyNyf3MVt+e3Q
tLEHSVnb4Vpm6jCf5KizjBM2UYXhkPL7yZuPrW3dnE6o1tP+mzqEpjoxWdG/R4zN
eHSuyETgH0F7Ngat3crW02g/kNJ6EmJTa8eK3GevUaiE+DjZHJWjuKnx6hoKZtTs
bMWBm0fiHqKansXo3WEwlTWzfo2tQODExh7j1UDBzmAeFWt4V5AgxGiwgPD91wMO
+hGBg6IR5vJMqY4t5IzU2oR4E0WOG7LAkarlRswdTHww0dZMUVVH2yAD0lviYwNo
v+D8t8GaqDi32zRqO1i46bQrKvuW2/nxCrpFFkc95hMBgPGdK4ySg1kAHpUHigMp
/wZs0GbcC8mWjYzWXASOMAL38Lp9bLl8iwb1L2uNozUh9LbJbhCLDDUjXa5ru1+u
NsJGvikcmppPR4WfcMJxuppTRwXLySjyqueLWf4zLjiSOMM2QQWcCvZxzndcPMyN
X/TuMXJL/oZhNbh9xkiINZrgjbmabSxFjYL9n+u3iTUeJZEViFWpsalBh6Lw8z12
uMM1PbFTPHm+JGsDoJMB0hFTA+vMrmCN2xTf0Db57B7uMzcMiXluMwMnWxQtjN8R
TYEUfws9jwCokQ97dKLbOGSC9aI1gekbbbWKTzqnHEPti3StY6FS045BniqkfFGz
Bn4mh2ROCsIowCtNdBDP3c7AYzyqFLpQ0enx8sD6Hz6jRBtaZf7xp/vvJd/iUUMm
4yfvVlwbFIYzIuuD1Mjd9mz6jckON+yGIOsI02DsjUzdF+yB/Wmhso4T70E/gVWF
uxQ7diizlr/nXnpjf4dbmdH0OrsQPN8VEsBNWTclNPyqMkPMtCFeZZESn5UF7j75
0okPe+jZmzHM3LhkSPQjHEBgwAodh9RP8PQ5McLZG4/R7abnAgb2n9WbJUBkDwzj
jxlit+AAcy2yrHY4AMdrh85HIB7K1nR2H16mjRuNtGOzVcO0ahK1Tb8417ikyFh8
Yp7M5C2kmayzPO9xpMnJNXRewzKneFJEjE3rmscS1JoHTuS5kxacjDMlx92LbiHE
zez0dhvQN6h85QLgvC3ktW/UYD9oxpdU6xAGiakqTdCmpOvQe4lVcyjLVzR+KYHU
3VlE5jF68IwXt/k3xJHX02rE2PVi8Lef+uRCq8b9lVF3HZ/x6aC/yT8c/E+6Y60P
g010rcgSeMEqHEx7ULZvCrKp0qox+PAIWL/Nq8wblO6u4O/c6CvZY7JrLfY8jOYh
5BoAK0NuNHTorIdQLCmcw5MALTcBQdeLb5EhIVq/Z1LQE1uUpWLuC7tcKnmwNL3d
5xq/bdM28fbkY3jEs5HCrN9vZWJVF7cQarHUi2YHc72+LzYZEvaFM9ij+CRBwSxX
HrRAktWREwheqNbuQSrjIzy8naMj1eYcqZAgE/5qh38CHqwH5wjIA7eOn3o39+ol
iWv5omVe6QuyErUcbjLfJB84/u5ZyPUCATdy1H4VRYXm2Euawb6VJYwf7vydwz8R
2Oh9cL5JGnGU8AcEf37HRh3VZ2VPKGOHrUrTlBPjLwWNIBqOKp+8tsJZpe0b7tWn
CuxBSii3LakapZ6lpetZ5p5RZPNNW3OegO1sp7/ZmxsWVlV80dfsk+ntFanqDBYH
5oyxjnLXddRqo6joBGIsr4CDGua+Os30y3GzJQCevGPAciSZ3dtTmFp+F5PW7SpT
3L19QXyiq5A3uSFNcpEX7fFwA8tgsb6Oe5tLkZaZMx+xkRlD16nODTnkRBdQK088
UWh507GCXqDecL6R0qqbRtbj2rZClgswk2d7N+/umxoMvelabiuZTkvANHMVBh/U
QxNXs/VNIBGQH8HSACsChJqzmZSDy4/xKs/YpIZUOtIyWLEpijoWlxh2KLuOFNhx
yb2EXE90OwowWRYk4hb7eM41ekTiaZfaVfaNCfEbeX7BoWzYBmBBKRdwt8ZwIrjb
kl8yGHsr/pn3mlQRZxjPER7eG9VyiBvzRwuiHx4teEU5jErYNcAuxaPfOnXa1vPB
jo4+Mb/jq5PTi7akEQrp+GEf+J1icw1z7VreIlITMWNpjT1FF/v13PXYJYqNAYlO
cf75HElGgiYjIFK8B1OjJyRN8sEK4jv4fkBcZDf2FkuxYbrtlw5iv/CylNwbStXI
+FeYkhXRxOddWYTUNZArTHk6ScsCR9XbO/AiMwNZeIvjR/OF3yh8iZO9Oz7aUdM4
DyADNiL+2e4X308Ffc0tCQqco+wqeGcj+C4UeCBS+fEA3/PhQdjzqvnptjopXgO7
Kc+4Nt+bb/yiGdVWotBVaw2MwWpQRsQVny7sSzuQMP8187qjJ5VIpcEPiC+5c/Jw
oMYO+5xGMzMmx/SodQ01//E/cvUfmvPKqkLoWHsEALDUOkMeB7nflEz3P/AdqSRa
qqHb84YZ/dJVSj++e4X9+AeHuJxd6zQ8shdA9ALsXaIi7toEvKiM/CQVv3u8Ooty
/0mNy5Wfkr9HaOwRd4+zbz1pXVNscQ3zzyRXQPZbLUBybshlzFy4SsBTOGRIbjk3
XnElHzGDCZPOXA6tqzME9HC6sBCoVl2BIkUAOOPi7KtbAN6S5XJtQ0E7Vetxyhvf
gUaq09eJKSoVQ+pBP6vtN67UUVe50PvPypVa6Lluc1ZJcAJ9IXksQVhuimYq8RLF
24qdAA6/8s0kFRCrfNXsqYpTwlgj2qUiCRtL62JPQuer4F5iBiXbFcWJa6RxbMNq
RQjHL7xyvgC0VGiEHOskUURhYbg+7o1grvTWFS1VtDg+JBBa4RHC2xVjhKstmYib
oE/PCKGuOZFyyO/6HfgHTEgjRrB+vUMDxi1Z4gjmg0ql4NV11EWDaYObivtw2OOE
zh8asXoslQ+HINRdpJTbygnQSz+srzZ7BoOVtSbWU1FUaS/MCF0jXf9pSYFVP479
8LWKdHEAozR1OSyJnWVvougnsWPcic9Eb6m4eIK8TVz+61S3wG59aHNxJwaBZXuS
9AuEg4i8f0LALBo/jqpuGxPrzTbo/aa6ilDe3oQYZ9jNcfPX67XEgpEoGfDl9Ioo
S2r/ipv/l9DwU05uihY362ISf6iuWtdVQp4Vjmky+QrkgNQL/62B1BL0k7sGR99K
tzRwnLRuZvCNQC/X9b77q3R7P9C+Ps4RmGQgP2X8vrWPHP4x0v5Ow50lGOp+12d7
kTeemnu/Lu5tJ3oUtU+fwqgv49w4/kGh4/T4bXNJNiEgCrIl6UR5jZ94SVnR61h/
81YMEqWnQaOfpkKVYw8H2J4+NgP7n0qCPU3bZLXTSaTpOh77AFsQnonjt0fHTivb
KYY6XAVxN6jeU/aarw8BL+i0mkcSv21Ma24viXiPlJ0SynEnNATPJWCUxIM+A3O0
j+3ERA8lOC98wbZ6loyKpqVRZfeOhYOeW6xBtesKG4oVYxJmeB/fdGM4Nfy6kIEQ
p9R++UnBvwFmkCxbZ+93EyKuETz30tj535d45BqlYm8Rrd4gWcqYIWeUYQgJSGHV
INPCaZQlMA9TvI91w9adhFZN99N8QbZ6BC47NcOGUGpBbAK27FG0z2s+fkhudzBn
3pKeSdHJPR2rhX85pxj3Uf+u71TUAKW7nEyx1Ymj2UR3nJSgJLnbUOV2wzwmogbp
Q/HZgtb3ELHERhZS7LEaywWzHXIkgVAanf4CMRwdKVVwFhhqsOSRsztC86YXpYF2
+VrUZFwg0s7zz2o9I+aDNxyINU9THh+loss7rSUB0+mTTq1Tm6oFbMbOemG750zt
q8LGh46d6oWRZj+u+7EjazVzwm1g/E6y51SwL6yJeR6W/sM8dIF2o7KgmpSfTW84
4W4gcdFtPXSDQGhH/D4emQNI8XnjhBzqtW4JAk1lATcCjXu5vQwQZhCijuqxP9W0
6ChrU17MGlCGVbMNDI8WMbOFh7njPTanhnL2zgGvCd+n01qJmprrJc4ry+KLmsae
ftKi213iS3VZk/5g3iT9xfuPXHfLLmic8kvG0J2ee586CjQN7v+CktAX9cLE/84Y
1uN37V09yhtp47b3uveoHJGwqKr0IT57dgstMi2421VG71mWxIL9VDn14kWfLerT
jvu/U0+fulzPi4lUqeOV5KblvCJMvdPRz+dAWgPliGFGQZQz447AjWFSB++TTrjd
CmzW2iiHhy1HfEXuJBckiyZj9AMCIKeT5kPiUaSx/DfIh20HohPT8kBerje9AEm9
EUHOYiEyX2zJarcQ9Lm/a5SRUt/57ga4GM96QhYM3rHnawtDlzeqjaagFVnrMQ6z
wbsb1Mv2kDKdl4hieCl2rBVjHJNRwx3WQ4hLyZ0dXjnQV+K7uYvkbTeOAMY+UiYr
WRT1SsvwDDlU57bzNMFQ2V0Ur+xJthPHkvL+H04iTqCZJOhugZyKmorcny4gHJUO
o6ITpBdbViREef3AJgNo3zb1kgEPHrDfP5BcCdK4/kP7FJmyzMDYbpQNKnGJm+2y
XzDaUJmG7wGlPyh+EHDYFJ7sPJp7eqXkbfWGJzsmqnbd9xuQH6kC2mixKURe+rG2
EjhSCOCYX7bscsKeZibsoKuW4YSQjtnwFylfzV87Ar/m/nka6tBymL7H57ohKqCD
1h21n4Qu17VareU/6RPHU1XdHUKBOsCKyHrulnINZ3uylZKWQ/1fG3XwPAIl0mbo
PUboYNaBREzEWcFcOfxPgvCsnkgnKrVZUNvKCnB7AgmL35EovysnTX+v8drDrxJG
YdwCUTkjSwN6Q7D9BASXvnnIqPbrNi4Tg6YBnjj+yjn9bJMTaee31WCr1E8Cug0U
kYlMRdrBmNQIysreCW3Q4tsYZWfRoyIFKNHFkwzxQrRsX5XzCFMdCTPUIk+1nFuF
vJsWaXQRhj8W203VAi5/5gZ90EuYqJY8fbXfHvuYHXI3ThQkHGsjQD5ixpaLNlpO
+PpQv7Sd9Yfbw7CYMjeyUq+V2R11Gfy7s7WOmVQa3pzyLdCSzLOwrVsixUuGfLWY
e45L/lTBmGIRp8oweeeLwR8WaiJfAZsZ5dKmRW8Ve7R29/I9GZcsbr9eMGsa2bRp
kyPfSfciW23/yUxsYvwQpQXKmUzPScvpyqcCD4rehIMayex4IDk1V1gFERe3e/6j
96BiZklyK/zhRlwZca6zwE+QYrtfpxiLCVNBmdgI8KrW1UwE/wicL+F0I6mR2wnL
GSM7r9IAg0VMdbg+LXlOsK5OAtc13xC0N0TtI4S26MU/vigpZ1JjjIo/C/eELxkU
QA0jQj/u268p2ZOOnHO79+6cnJ26axdac+D0aTzszF8FvtZBOfbpcG728T9N7fHk
m1rdBvRQN193FhpsMfHHMi+6+J4FN5eL5fRNfDGiS6I7qCdRxJbBwtoEnXn9w/Ui
ay1s4MoEBuq7IYnL3uqG37ZQGg47PdpiaZwNtwj/OQu9Rm3Zh1SzVM9Ol5po46Ll
ab0gcWzYm5CMxdAMTN0KzBKYfAnyvut1cEiYs4xW5IkzDXATJnNBXuq+wM/rObzr
hfZtD3F8mGVOjESRXBgLE4QDPsvNSm0hkqCv7zx9fmdRPrLCPfk+ja+wvr0geHsV
Cnq/VvekHtGD7xR5hxkKUza8rPcpBkTRDclvjxcgMCECQzyZPEJ5Jd+IWRuac/x4
kPyjbQfte3nSEPxxcEq7K6RHRRqN7w1o6r1smj2kWu+XsaT/GS4WjAY0mhB3lPnM
6+GfTIbokFxIOrSEKqHfPe1ioj6RiGtYih9vCQMXAMsCHoh4mBQljaf1yTWzrWIt
emaLYE21mtoxkBfJwmcpMnHNgb/mn9o/xMByr746qBdZJn/oizgwNMQdTkfDiXSx
NrqpwKg9XDf5c1ALjXuigPG+v88IOX3gjTzeuBpNPIQVy8322WfQdBITDQhr5TLZ
i/ZbhwbtrOfnN3W5H96dQD/KUN7AXGYGwb58gvK1YdeA2kMIwsck4GrL9ii34wNK
41P3lrOhg9wZw+IQYhCtdK96+yKJ8yzEe/p/lqFh+4ryWJUsb9vs1rEWqAaxVVqx
hd2LNcZvzdd8m7H7IPY9/T8tAJ6qXDkKPJcXg4h39vgfxdBnQdhPF6Yn62POyqez
VEIrxxch/LICyDGqkBsLmoAXbbw8rQmwnzKJqZeedzBpZsMj84UEP4xCLklZfVTy
u5fBA4TBmuMgpOKpl9B+86/mCOdexoVYMSYB8sx8JxW5/ORWPiGQcjQBIlU7jEbw
snoR6WlYbYIsGABXFsH1oUGzAAuytrYDx6xvp3iYxBKHYkGX+VcDduWE4YOihGNy
CCFVqer/mSRZ7NLnrbOPgMhrXeRdo4FIfGs0iLSceONDoF4I8+FrmR20eADS7Feh
5AU5TwBshpikImGvlS3piJWeGLBovUT8a+6qSRbftqHuJrJxsPn5/IQXjYgusUJC
kMF35mcMSdVGyvCCIImu0L/nyk9yU72OxSPa74HTD70eJAvgn/e+bm0UtytJA2C3
p9FL222hWhKuHbEI0Mc5qsldJcnpkV0i5jqZpDpSLa+gi7Q+Lpu4Bj3lZ7wQd15k
zAWCENht7K4mF651kLutn2u2QSSnMW77LqTZyzzis+wTAWwW9QZLMnwPd7SwDs95
py2SQJcrZ7KhlVd40A/WqWmUsHHMIIFyr8E4cWGKWA4Ob/RpELp5X/1kRDAsOXMQ
HEwsDi/ymOTHT2u8JE8YPtF+lDjsRWXsJgEPBw/u5UPzhMkN/29J0OsvdHF38E7P
/OSTv70YVrr+ljlDgkTVlZ+GNtn0wB131YXb00VCchLKjkOOb/1vf0A+FDxQovGC
+sko0kc+C5yuHimGNSKPJ0yJr5kBYCnfWEGtAd9eGQ/jrmU0YGXLnGsC798u2goS
Tl6NeY7Vev5lQz0x25grH/P6w2kES5IrZZXga+CZmz2tase4QNLRdxWVmlMpCFsh
GAvHTBBMwTPwYKVbXKkS5bUKWEZ7/yOhaBeK+2CL0HM/IJLxNjZ557YATyyJCHJV
ILXZlRBMPfo6UARES9AVNCUzutGxZpwWBJoT53ZMnXJaRQvNqWZhDgYQY8+Mefaa
zhGOWNE8c9gwkTuoYkK+M+Ha0YF31Ec7NfaxHLIH8H15wWcckZJCUNQ9aMx29zqJ
rT+Eeb5NGtk7zlbspZRcGKEcQHdUV8S5OlYsZUsKZVaxkcTI5bzrnmlTluWavzA3
dABkVLFYiz0OBvGbwbLjuI4v0AhjUXCwxy0sJucI0bhk1QcwCuHpL5jGesxOJkQ7
LcU2dWcbkCcI43CziikbUPIAId9+6aJ88p4GQUZ1uf1aaXJ0b33jLzQdxnWVDgxH
RwdyneKyfpwRNh69HCa7h0hL6Tf+Ug9T/aXU0ug/EKHPylv0n7w4AKZYu9C1MqTU
/9Qx2+4/X6cMaMx5+R6ueqbCnBObMbLu27NO1g1ARJ6GbVEoLEvObRnsaGTiBnXH
GWso907CeL0B/3Cy5mbGnhtW3M7gGZQVHO19RRzh7HnqCNUqjNMf0frB8Xdovr0G
W00hnxEPwDG+AnVs7NaPPvhPuSeDxICqQvoCGyasUB5aH5KQDmfQrCsrSvLKclHu
wI8QIAj1NpmJOXHtbyZI0v62HgdehDna7TrDG72wnM1XHUZ8AJu40+lngQo8uCw0
McRWmndi8K/ttmidWwBPZI+s4wDq+JIbwUEgNQ65HYzSM5nCp7HeLawNZRtN52ES
U3DDoyLldYq1oMeCmOXWsKzNuPJUzT7JT4A9kMcrSmZQx0vMA68BwSjYEioniM5W
1tci7uW1Td+0grOwGDTrHvFJ2PR3PeKy5sqzOlKr12hC4vmAnW8+1T/S1setpMgJ
ptnY9iKWWPai/4XTzKM6bE+YiQkQeKcmjzLBwbtuz/YdNyROk5f8ci5bubHSRX4l
HP88udOH/XptUV2cyJR6lJuZKSGwV2A1DIshv2OFaikvDzFTxC7eO/GQQ3jQroR0
M7DFHhvKQJOPfanYVDcLviodG2eh9vWd64uc3SmsqYcQ/nImcG0zAEieIGqeDCRq
D/U0w2B3wWEPu7wJdMI5bIGFik1XMDxHdboXnS05TUSxKrKfA/84UWQR3VU5Gif2
w5e3UdPv5VyThRadc1M/0MtdmB/CEiD/HMnDPSXjV2MzEOuGX2QzTPt31cxQkhW+
q5deyI/wXu1mEpocz3XcGwsaKQR9azjOfNK6tt1TMCF0DbLIcgrEyWiOXVZ9f1Eu
W7fV3zR61mayGPdhtVNiAn/QlwyBnG5LxO2SDE12y3gp9byXsXmBH/0L349QiTWf
IWYN65wCG52yAFRZFDr6xEYsReBKn8Y0DTPU9GkpbhQhNa5MJuW9w5+kqdEgdD3X
oQz5Hl6FtzEgvuTpTDMwav6WpmfLnW1Aq9WvQp1mohFFMHTArsQjiYh1HDqx+EPQ
vToGgCiHOMlwz+Uv9Mn+Wgm/CJUkhpCswSsVJljzZiSjKUUgDTSfQP0qSMYeDZtd
iug5sj/Q8v8Lef3hC51X4HR16C43jGjXtlcJ8E056e5DPWKUZY8A/YChcbNwkhBe
ZzrtK/B93oy4JGEWRYxv5eyy4Z9iwUANZUy4kYCb9xB4nrF0A51i9YexDcxB5nDc
uDhAISBciqE9k3kYU0jg99u566cyMrF+cgRlJza9ZKAe/Jb85IdpoGZY4Q0n4RXs
KuFcv6NRQSxAzIgDa6utX8Dgxo8yYiDkqX8REGz5dO+0070jJhsfcQ3wPyEwxOE4
PU3cTil2LHoKpoCN8j3At4C0WX0aPTQHV70cdbkPN3/2M/DA1g/nT2jDUjdCH82v
YYeHfpEXhH6i27aL6ZGQj7VGGtwBTGil7Y1+Wa/3/qJ779f26sRUI3mjTuTirBKV
dchCg592bYBhAJOlxIW57HQOs9EJglyT6C/ah4hLTjnRJYHo4akUicMGUVmdIeiy
vsw2UJNY3gmu6bIbFRWQHEt/fYNv7/z1xrrmBARr8XX3tfv9OvZ/UI15kS04iwWS
1gaeYelhC/sHn4iQfqr+/B+G24UNMI28TT91Txz2mUiGXrbL9BFI+R3YY4fvOrYl
ynN9E9GsBai5FA/AUw5MqfhWie5BAQFqgVCgRFTZQSb9NGb+NURLUTGcVovyL9mj
CvI49ua4Spm9c9nIKTA7/taSyEtbwWIRdMyQnJyQ15H8ETmK9b5rKRVjhhfiTxSI
tC9zeUhpiCfcfowXUQvvy4dTafcNviPm0GZ5S8zHISX7Gskf0YHMAV31xp41WQAx
LfWaYQgC8Og1TfH/9073TpD+krqy7hMAlIIEe8pi0ZopCdy3I6KPLC1tNcq3be1P
mtIdAibLgoFQuGCrMsDuZ2WKk8oQu7isp4HUwMkjRnjvZUX87trusXwTbGFguo/7
+GwMKGffiYsPMaxmklVvyOwDAlCohQDNeu4E2kvD4HTYnD6qzc/eNnUdckRIowyY
Nll1TUxMTXsz63HqUDEk3pc57SdjFRX+ylhNfne3ZR5X3ncekFLHEdkDosVqO36R
16YLuRmN8Geqsr8wBWZxcM7kMRA0e5xyNQKtRVh7KVcH33NqVODq9ep3w2HP/ig/
RPrSZ0846SMsx610pZjZ4M0Yv1v6huh0hSnVfnNo34+qR8WSPqlLVaQalFpDVbDi
kGgQhY04b/VVHpdY7bp/qMdnx97knCc38ZeFNizlZF9B9yV7rcj2546tMHSzJuo2
DTaBBupho5W4nNAwghQJUkhoI9t6XT5PtcVlP0ht4/5OJCntEXJ/XvzzIP1bVgcU
zfNWNo5+CSqYfAg7QvnOD2uIypTEJP+W0rQAlL57/dMbIEwpRAghq0vZNzrrJuZx
UTTdpMkehh7Skx+ZF8l8aZhK+fl1yIvMEYqGrqEiGJZUPivt1zlirqROgrf0Qh1b
31RAT3zoxEua9uxKI8gGtUfnIwNkMvT2CLRQkPCAMpqdIFgyMA+AwmzLswcXdtZ4
BXEeUFQktX9u75cNQaIPFLFOHOt+sqB8+cEUjgtnX+q6X6cnU4ubK4ICdfo4TSwx
fB7eNYj9oykxlFFGquE4y6IxFERokyQN7SrVIvIMRYmAXcrI8SiF1Rsi9omKsvMi
jB7xbZGMnJgP3hiXGxLys4wW9KRJmfe7Yt4Qgq4txq/sIpuQRcLRtJVvA3bpSGTB
sIsCiNUmTFMuRmWlDiXODZdS+U55GJYtwnMKQIk03JoSGZ7uuczEeGvRS82tspYe
wDwr2Qd8ReJ5776YOkmajyXmzl+wfzZtq0U0l33NTISK5jsD8MzyVYKF3IVJ6ukW
jBkRn2LTFMdF4uOME1yhl+Ng+KFuBgR0v0H4klsVLKoNPQ704Sim0e4kzIFcQTkD
EibOx42iEq0oR+7M05bsrsh4mksMMEzhWPwj5RrHioE9RYMOF5A6cbuvLyPeiAMb
iX3yv+t73GqxVf/lqbvJmnXQdKl84O7fJbkvhPKjcotSsDOu/chUTbtHd67tAgfZ
UcTFUloHXNSDDEh4gCGN7hHpqXRdhReA74lSLdbjW/ckVsdegUUc69syRhuKXi8G
C5DLoo5PVzH0ZhnTFrmnY2s3yKD7uDkuJtkzKeUacJA+2LEtgys4jV6rsulh+a+x
DlwCUZGnue0SD8cxIRGyhd6opajVx/LHP6jIdahuEHza9EjUWFLSQrLTj+MnbbUB
IvmIY50F0SERJFCX1uupnOMdvbwCN8a6GkJgd3wvy7aKZ44t/sy8/i2MZFNQ9mkJ
hYWdrM9EeVp7NGiFsWRjYls0d/vU7OgrAV27C+snxznShAJ0+1V4cZlgEQu5Rrb3
Kf16HKppcQ3FY/U6QviujtChUcpRQqjc874pCTB6hUFCB4vmv4Vax2xaL+Mcp/Hu
H8kacN1tfWaimfm0OjI/Kyl9dD4Xv4X/H4uTZXhYmpH1oJLcbfc1eF+63x663zzY
XT2DM14f85tK2Qwo98B4YEB4HfICMy96HyTS86HCd8iMH6kBVaehZ+dg6CpVznQH
CwfHKBx2flaqG3Et9QgzRyr9mn9pFxzETXjt9VidjfU1t3v12anht1aWMT38IWMi
KMSvxPBJs1Y2ww4LAcPvDUcmPjc/mx4Uj0YCCbBLwv6bBxILSNobFQgatNiBHH3k
nQKf77ERj3sjHRGsTgRr4k1n459wcUM3gmy7+Lj0kD852OdhQog0S5BKCXqQAhLE
bHplItBN3oky/2Z8Fur3ndB36mXHk6tKnPR/iydodxuCs6jT7sIga+l+O6RIpBk5
ZysupivuAClbBrikdkv1rjiMDomP0Wl6ZvBw2xgGbFKQnL0Gc3YSVEwZFX7kHkHF
Om/SZpAWi2K+UsX+OJePbDLRAsWRYt5fF9WM20duvsvCO4elGpqGRvGPxG+k1bXC
0spVLgEbJc0/0VN2kty6oLkXVl2Pls7KKdE6Dbw5eTkEtx3y7IPgHEBuwDo1H+z9
kAp3egkmV2jCon0wsWTWivDHiRw7WVlQewJILf2MMUImhQG5i6DDCifHz3ljdpqa
fASek03hLRXyJgMNwy8kTBzS5yy9JXEebtsI8ztHA3HlDuf+Th7g5ODCb3QXEKxE
b6iLJu5uwG1VEgJx/KKHop/3RSidlcIykxQeG55fnSey2sPFbn48JQYDHcK8L12H
NFqkDb4LlQpprK5QwUFGI2n/kZbWCKf2q77NXlttUjW3xMDh6yVtXNMFy6Gjtjov
52HyvttsZ9piumhJXMHI0rkOZDdwBHdJ0ho/vVlDyVmqBJyoC+5N9Fvmf/ncUjQT
DLkb2kuoqvnOqNM5GZmxLTQKUgeh8HVfwjOGSB2UazsF7qH5EMQfYB7YqyyDZL0U
9aioJ0JmMteX4is7VZ83D3oB1HLmgK667jQGDNfS2O5Tv9Ytd/CzSVd/uCw5/7Qh
jjkFIHLWsp6uIYYGwWwnahFVhBSBCwM7Yl50QRnLnrmLDXy0yM5+7VCVZ7EHAZKq
GSyWMrFXGUIfwpPS4EeNDyyt0tg2O/Vugh+1xlz7XSeP6fneRVkJspofudJ55Zuq
8OQTPxY2E6+36NyKCr3a7ui77t5MelHQ9AY7aHsxpr8Y3XXwUNSdLlq0XMMeqhRo
SjwkevppfQGZOHqdC19vmS8ok7I0Imi3zGwUG5A5YSPIJ/TV758uxsYKcdD4n/GW
F4+tx3rmUzJV3YXgkjQeYGEvV6wXbZJUiHrAmmFiIl520KZUkStQGZL2EMpcwYZc
82HvVTiH4j7Io5Atfj8a/jFcOK22Vm5O+z6U8Nl5Sar73ZNMU+fTTY5X/dZusqY1
F9fF7zUGqf1wJ1+1s4CXaxQ3wzKsv3gqLRxLZgG9HTtJlSPsx6Y+QiizKE2bYTld
0fPku3b0AKFCNFJKFGhn2f62SzxOwmitjsMzR9M2a09f4XLnqT/srU9p6EjHRiTg
ahuT1rh5iAxZSibr6Pa41VDOVGInO8/3ByckcXlZnXjyWji8NSYehS4MVRljvLaE
QCsA5P1OmT+hAnQSCin4Zv+sbzThbXC/YuPN0S3yDDeQPjNqfuKN/8ak/Xuks0Vv
HRV5IwzvgL48oGkV4RWj6FD4JXD5LD7u9yCJqVopJVDGWgU1XoSDNd4Rrtkn/FwH
tZWFC83pwiChcbB0F+zvlJTUeGLhl7kdm4eg0M/0IqCmsRJmAOuj56PAfnsxgQ1e
I7nNPSVUiEpxpn0PukNhFJr07wDBNdoMAmjBseR3x2+so6Ols/T6qWRaPrWIf9ye
puaduJ9Qq24RXB67hZruqMYVkAPfhmvVo+setOOiNLqA/1ymhin0LQngvA6Ny4Wu
rPhCYugTggdH8iufHVacOUXM2aCqoqz8MUKScFwSUNobxBOw+NgBGaUxr27IDyO+
Juz0itLl2HRaUg4iGiE1vNQ7u935JGltbWqSrbKDywGpKlBeE/cHBjb0B7nY1daG
pOXAYIk81NNKHVDqevQTH5vy8q3VO8ZC7pTMzRqgJL95pX9TgfFKbb1ap/Zi7oGU
96FYdPCTgrovVtXjEblogJAiLPPWAMK8sep3QI47a0EFFKLmi+MdKXGvM8/mPi+u
SkwcA+0nE6VuPOcxFZpXiJiOFKaJN/0tF0SkbQkTec6gm631O5vHB18yvYTSSbq/
rNpsjI9wT82UyZGDbMOYOQSqWxDYUpsc1Dxea6tr7HwT1SD1/pCrOB5NSSZHlrKb
h0N6aen5SlzWhHBjIxE+imbODhxS4olYGlPrDQfj7ZNWEQE+AnHBZRTJpV8TmFJo
XqwdymsG8jrfzC1uL+AmZ4InDBTmSSkM2n7/AqFtwc8iLq47SLa5Egn0YuYrPH/a
8fLb1FM/XNPUDwHWDsDbQ3OcX0OLtgKbROMzqqDk9NP+jF+QneXZgIo058Ku+2ko
J7s8BInfykzNAuRMx/BOWmF/i+hSDo+qLMmYxPoN2DzS8u6FLXWPefyy3okHgxni
rWeyHy8ANo4hN1OLwgCOCnqxQt/E5oNBzoCkljz6aw88ui1fqA+sC1FRxDHV39ua
7/ioAfqJJsJ1d77SMocs4bEcsRU+YlyT7S1i58aBGhOcEvCSk3pWlRMz112td5x9
PYCHx/jzUqfnPUALkrBNdwD1vOLU5ufsCFgSmiHw516qP2qx5ieh1pV39CdUa9X5
azocGCP7b6wHNTgdbARbfgC6rsa+qlsQDacE28deKI+QQ3F3o65MOFkeTxF6MlzB
hP3zOMS2BgwsZxSmikY/J8J9HqeoGP727EjbcO6+KPj4+TspNicbwTW8V/4aB67m
RxqUpCmAcHrsJgcYROU4Nhg13lub4QtoZs1NkC4Hfx+tX62xKposZTeZ0PXBNZ8Z
B28mTKpLESlXqJhT/IvgphxuHL1ASiJmicIp4jeQ7X5IHi599FFReyereu6Iu0dD
DC8y1DVC9YJrEEa7tduJLh17eUSdC0Ajlxb0x0u2MRSqx6YWL5DkEzcVXQz3IrbY
42sxq77E9ws2IOQaseX8nCPozY8DD+XmWtf6rCBUbaXKk+iq4frxhIqHre55sfFG
bqaSOemEfsVcsaFs7w65BTuXQkbfMZEaGXpYS+CebE3wzZ5jp8FSaaHaqv/w9RS8
s6l2Z4J74sKqDoBiZCiO+EI2pxrjxqwxO9wgnjdIomDUx0rmyA6zamTj9AYsvrYf
C451e7Hhe7rC5f8KVtD71nMxzOQbQroQj2UF8LySOk/sc6xgk0gS8TtibU7Qg+lx
251EZp2LQf7Y2uWKcTJQ0G+4gG0vkWDgkmyn0sxFIeZhEeYTvTRpOGQzMz4OkYkX
OEeUc0xUiIZyofEht88HKn1xryu8PVvCg7J0saE3xl2k81sJB4xVqan2ul6gz4jc
flhCKO3djdjPU0F5YeAe+fD0Odxg1ZUspFoMwt0UOiZ4DrJbUVeRIecL3cwcT7Nw
UA2GV/kZOWUy28TfY820xKibBu2ebredSLeSQczlqoEFX6ltOvN9vpK5V12UrPhz
7ABTo/RQ71ZwIDDWuPjOwzRLonPIJP/LgH6gIcqCudSmdok8DVYMYJi3muRe88mo
gVnwDMQtwS465d7mRWVRaIzEK9teZqS0TsCSp5obN0b73W9qngBNcESATY3a2JJK
0VUVGgqOUkbT1AXq9nL6BaTg7Xvrc07zSSSMhB2xzFeBAyIOL4Ys5+MIuOtxGUke
CAzZYgS3lvkTvhb94u9RpwRBXt0lC8Hx0C2KIFAutfyNuCvd6V9s7ym+jPTRuWcb
zMy5BsHwJubEQ4hL5s5XgXF4Xp5t0sPzqVyMZ/CWRVGrNaF8HFqJClxfyr0cHcwK
eEzklq2cX0lbmfA1VVdzEatskDp9stD1uQ5BwhhMvKtqTxnInd/bEC+y6YE7FY+a
Rzkw7O7Zr3hN10CI4wnwXCKdrr61tw1S3/57mpgaAo9zu+0ciy1eSvFvKhRL25/Y
t1zPpNw1WUnT2ebLeTCIYDS7vArb57MYXetLNVtw3aH7FcACMMR1C9tuAQB9Y2cU
0BBgS+MaIPcqPZ7HMXwZpCYvwrH6/jTO0JjE2Jjm0f2ym+vzjK6kAvn0kVe7kS74
l2++8iLVvF1RtII7PZmwXQc4dNnSaxcn5iYweJySpuQyURf1e0uB5/GC6Y7GV7Z1
w+CzcBTlvepG9coFCKgbByy6QknYUCdXDl5amAY5G3gru+zgWTxEPLA/LTmSUARy
7ZCXlTK3VVQ4SNPD9ZENefsPRTkDWp/KH2PtOVatpQt/E19XH1+0ZNL/tssvfrCh
bNSiOos5xsuzSTOQRXGpNEzHcRFF4oZMivdESr9UIqA2HfJIPw2ymF+i9SVNAICx
RQzEPWjMNvhbXWS7sSl87yNJPp1p66Ivgrk+LGbid3YzpFwzkLmeth08XR7KnHzR
3kkZPSDbCtpVGvPTx/EDkLx0mUsIVBOnUb38pLet3aXUKhwO5Tg776X42iCvcuDu
92Gi8TodXdVfshs/eohOAxZwnwEgbP00OCDa/tb+F6+DiiEQd3EFo0Dx+5bYctcR
pzOjoIMIT86V9VvYz4KgfJIOU6+vZuwV3bSkw5ii0YwrzaGQAirOvH3O5vuOGDoL
pCAGX40ePU1gecfpJOryzBARSBacJSw39nByszS/HGJd3Rcf5qbdxKbO/3HeGgc1
pHYE9Li2cobnyyeNpBMUAoQWXkfXqsNTNhuIiUmd4zNXXA4R/LzWW51jd+CfByeN
b0NkYGVDjti6dRg3RUeWwTBwjAtx/VS+CR4BhZ3iWoM4GxksTWAUAOv91OKCpwFv
fNOR7bYchglPL3jrLZLyp7z1EBCFITSqkid7NWrPCOahhqyoHOuFgCYqJOH/Jlt9
jtbJmNFWKMNODuUGOrVHKiQGhxUqlnWsCHwRs1mNGO8nKB1jVwpQAvUVw4D4txo4
ysHEAjyBCEIYWuc5NyYkAhOZuetScXmKxth2YVVLzO1KMPqNcoaJSu1tDoJp37R5
e6tUP3XFNdaeZklcabnuePRD5cXca7zzZHNxs2h7Q1cPxkaK24TqKR4idLP0qn1A
0T2NzHzDMwomAN+924c+eWxqRcVMGn0FUt0vFbT6kSTocQWoTDaw8sti+ko+MqBs
WzEVGYeI9N4aFhPe207bOIGf78jISQPkJKNQ3AD+t26FZrLmqdXcNXgLegj0JCed
xPRIcdmNO3KPUtLOQRuu9zsdzf5bDURhZdqbnRMZ5BrxoB5289mXqnJZyoM7/hUN
3F2t3yOQ8f/ootwWIVdsh3BjdzNazwvcPXvhn2yJXpEJ95kXcEY0ECvFQPzslq/h
8h8Saj0M77nNf84EQQvRmWoO4FvsJsKnIJRL6odVh4/KVp9IFAxnt9kQmy+Vq8tg
EhYGNSEP45U+zUoba0FwJYksSiiMSI8iKK9UISDu/RwBgPoRjEtU8+/W83Uwfg97
3VI3amQoZrP/SSiHg/Qdqpe31yazS298nBhxyAZcYFgfwtr1C2+k1DG6uwMn+Gaz
MK+7yM14Z0FfY9N/p8jZ6nMAAUrOsXvSqQ3Ba6+QEO0B5Kz9LkAnVAsinqfI50zF
5cQr7gKwAHNNZNQGxJzaDYBjO921FJfOLI+P9BoZB/HyHzxS+Gb/p1YKNWIVe9gc
LvluKpxk2VZgugkrIwQuOFWopihOrjNaJ8B4H6wUREn3z64Uo2hkrZ1bcIJTdiao
f++eBc/os6gQJ0cgSr43V7kPDi3Rkk54nLr5/nzl2PC2/C+1XA+znTVaR4//JMNo
aWFpnz05TpI6RVW3qCfPm0QQ2aNrG/IECzb24mZVfl9irY1OwzBvKtwVvMEcHPlu
Sfv8oxjmAYsNGtH8JrgHTiLHPkMn0SbgPYmp1zoi33/kBIckQ3Ykir3fxCpx+6mb
yHXYO8yKl8/WlQW70DeyGGUxSSqktKcnpw8Uym5qCte5FiajzckttncaNApfwcr4
kk4i+tb+BTDq7HoJWQjXIbHkkMiQ+NQa5lvAJmahelyJ0aCvT1bEUTqTqKjL5Hpt
8Q93ejQRYUYDXFmph2izZhjILlSSrtmPntqRxqfB6OwLFS5z2nb+inrhsL9ALQlK
uhLK3crdwdnn1SNzk1pKpbMNpNIZuIQiJMigdtzHkxXG1UZGb5Wmf4dW3P3R3eDr
/UUtC68EraU85NqDS0EmUXSI6nidjbiZ1cQpf+/S/iO1ZBsFbpH3/XEVmJnt/UrB
LR5zOXrfu5vEtg7mUSicSAqUgy0grliookmy5dEvvj++fR2KqIjRxQa9jdqGbrI6
BrzBKPOH6eRcwSKzA7nvyaXCiaCzX7+8jWPFzes8D1olxzoSeNVwrTZf5YP9yskg
ugEJz/1zRzSJ4YX+U7EIknu78nU/9pC5T9EFMJFsi1oxN9LgY6CkrtEvqgLQVN1+
JYxoywbT9bJF1J9W9t9CtnpXILj8jKV4CzE2ALp7G6GQWGp9oLfrtQiEVgiGHvan
zZ3WsNqMogqEZt3SM7T9p7yGyowYOte1Juci2VEbSADUSwBtAgarbxxHo/fC2s8W
BZcngWEYx+Vm5gfb+NeszC5GnJmojzHwizVN76aSTY6H/REO1lTz8i73Y9eOyIi8
6CKAX4GHNbrySg1iKzvBds1PS4gAu3Z81CJSlyXwIqDz89Q/lBIvIiAOEhO44fkr
V8vpm1XQqRB36Xf7qjIZ0NbUo41cSZ3tWnQ5wdCEv9lgPvY+RCaSzaJ6IWC89fA0
LxRSMPJ/fR9MY95ST1qi4Jm0C7oZ8p135uelSqrEzQRa9SwddVKoge1Sa2jPAtEx
3U73GbP/ePlKN6SlDd4xo2kQoRmpLK3c7nb8FKDObpR559D0Blh9v4GNpnpeBh9Q
sc03ar4x3uPqyNBeRYZ2+YAqkRjmqPwyuKKc6uZVeraZ1+Yw0A4Ox/Y9JfqM31j1
3+c/FFnXNfwUOrjycIWenpN3ip8LappdATP9QiQlLo+NBEW0BrjIYOzp9TDyABs8
n5Bxxrn+lUh5aOIuRaSNg2429yapMcqJldRCNygNMl1s2aMMC8I4Cm3YN6pGlOJn
LaghSchwUOLJHr3cW7F4lfCXcVYnqjgR5uMg7hi/oMB+Nm7LC7+ChnXVOzyWKbC/
6VkqBfl3iqU/+9UTS/z4Li6nGWUY+nGnq9RrdcXUbcpDSzBdTyLLtyO8SypAraqK
7YravApxMmsw0Qx8UNToaOI/FSHmLg3/v/bbt1p++4lHEmNzF1hB1ivSlqP4Rn4/
VPn5JTocRWnnLUV+HM9BFzreJ+SBHV+hWtBcdWHMDZtUVQqq421wmQblOs4aOqSa
aPZnxMINyXP56e80KbVrfkXL+bjhUr6GRyXA5gFT5BluCpabkSIOBljbrIeY3b8i
RAoOXx+jCzCXj7SjeJFqtkhWjLw+hPipl0n9vpLIQi0Aon/FyUN+ga6jwtnlMSib
InUgAgUps813M8sJ7uebgHzJ++l+ZSsGbDMeLB++XGClD0yA82K6aJ0hgggL0plV
mbDru/fxfAsODNKJCaovR9UIv2/RQEMDUiE/EBrScmJRrJEcyJgZxZxyiAz7h/ty
BKrreGRwE9nDXbhGu8ntx6H1rtnPih4WLacyFurmWaXLqoleCbiyFyKKtAIPr9Lj
KcnD+oOblCPF5jo3J6wjBe1J+M+E0UHcFSU+rHJTz9V+9LImDhOMCGSgiJFts4Ve
uwWErRzEHclU3vdSCIUzv0whZXUytOqwv95TpEGBcqsO/c1lWZ//y5GjtPs8hpA9
ebkdMlIrGyNiPICZAaXYav3+vifP/8CV5CnJbZw4uqPC5gCVv3aPO7KhqUsq9+Ci
pxEsG5VaYlq9m+PbEurWtzWGQ9yFWaDMEq0MR2AV8Mi9lP6Xl4mcuBiWFjqPs6D9
x230gj6LTxPcAz85jDzXo+Lz7mzPtQb2ZxBPUpdhrWWf+siFN6TmxMMiW6E7cW2K
4IVehlLUcXnixxg3Ed4/GZi7Xinn+wzjs607JMtBBKCp+XLIg+xxcrsPjvcsHNUn
UgoNjUsSi/73IcGMWAmabY0ok1uiClCkcsSWovBpZSWzSHEhPkxWj76o0D6hBu3k
0+FJ2hwGh/JQ2QRhsi/AtlWYIUriB4T9DFRRHWzrTGVZSi002oYjyHCRS2WZdJ20
bn/qbxKUc5MtEYm+UZt9U1rWDkhU8p2ZRAg3G78IbK8D+BGe9+Gc8pnmKxS+11/c
N/RY7SArbJSZug8g3OAgDdiVEm4+pvYOQqRnaDLAu1X3dadjLtVHmLLBGaElW5rU
wT58kph4PC9nrWuxT4CGTRJvki78X6t7/oy70zOK8uTHdVhqxBczDNkzlvSkSNav
6hMaTEkF8DtPnXRCzTG+fsDsqU/8+CYptb4GRB/i5GGvFnf+ml+QKiy5lgLDRSJL
MrP2qosohQNRbXAr8IVxB9PO71Llz9/rlKgW3ZvByXB+vhnzRvhoCWLNj1LnrXet
yRI4r6tVSWYkVO0zXoIPU2EkmNkggG47opOG8Ue4zw3ep0TlAtIGFt2VQYXf8tyl
NtzHxtx+ay1BPhSaKirRoe2aYjfw+G1z3T8nj8PSeoLnyIgLH2tjV/2rLhDk+d08
AMjUGzXVHvYxP0bO6AKIhOqVE6vDUNaNE6JvmIIARF+afEkJmC8s9mu6zQfoLqft
NV0aAaWZ1ldZGjF/Xw8LiIUXEvcY+aTxdiXo7PoOrO0BQ8XijPUH5fsqvXFdWp3S
AQZUO+3gRP4MYGoU3oXksyDPTsVCYEANypHJw29VWw/VUG56mHedWgyLNEDBjgXL
bwYQKmP7znQtVQZy+l3+l12FTfYDK5VyHsqQRP3VIg22MG+0EeSguZN/BvuEKe9K
veRs5YBsbeocKBuTZvsiu43q6b60pN2Vqqa9OVpdByrgvkSws6Xw2RCK6UD7ORwj
oIxGXiUv0DfZNm30/xVyZt1n5sUhNdhx9xvSIeDepCb8BjIXtzU7YS8569Xx1O7Y
XITzN6GnYuBZ1dayF2fWWZalfD6+frL18YreCoeDvHrHIlFP26o8qYvm6GOZ+S06
JJLgMuaaUhhPrdsY5FP5hj3xyJndTKv6/8YZpSZ3HbjpSGrGbPbiUBphS0NSjElA
I8eHZXNZaoW3Qas7KSh3yF0UGru3VxGh+Q+BIf8iy59vouGAXTjaB+mF0jlNzLve
Wx03KVERDhAJ410vhNZeX4HHNW6Ys6XzyqecMcVx8X54JJfxK517Eq+2556qWXY3
nmaffVbNSBduicpvWOFux/NWFnicStDXn/dP1x7I/8t89Qod/AtM8cH+wnUYBLBg
Fy59UuJ67JpGE8QV55CjEeuqoYzDBocY/M4N4B5HLcamIYVgfUM8MzeS4R1H1xFK
7AJoccfTakykCFjROQuIaCpyFuf34hJCPSK6VsPA5lCrQsyCNMo+8MExz9n/eMP7
dA1nKEtSZDixx1Jrdu4X1EY9K39uiKe4K93BDtoPk2rkUx6B4ZOyosQX9Sts0hYs
wa/n0sUXOTlzLHnF78lR2jVvZRHXaGb4Ywzifnnjzk0mpTQRHIRDD65V7g21ik0N
NGTwVJ/airyukP00kno7X9rcLLzFd6b56nFlvPNZSQLulp/srWvANwrc8e1CJWh4
+S3oqiIYl6oiax8xJ1GOaPSM7HaEEcLczjby+E3xpdW0ofc5KFuxGsBZmrfkXx5+
uPUX/BC/oob1XP/qtgMuAug2zJYOr9jhZGtESJoJATXRQmALLnuOwMgvTLLEsHLv
a4F1B9orHCoTzDNoxuoUNFnQ7Dq/apvdCNScUyqdY5vR65rRfgOYklQtZ6pGWKE/
zWph4nw+oR81KDrTh94BoesGbQGLR9Vp2zhiMpFKC0fkTiM0X8nwNdKIXVb3h8Hn
5FHxDsZ+1RN4nsRjjHMNurET3A1UXrqjj9iboBssULVSJZm3scQR/50O5cVNbUHt
wp6EJCXYkfyi92U3MKrIDCm5rpmuMlh1AHxbUhVJuKj/fFKnu8i+JuwTzpu6AvyM
PLJl5FgY/LwViRPFqcNiVmbTs6Hglm0ktafSXqq3czKTfmN4Hw+7I+Ym64cQt8YB
i9vnLp+3Q94KVBHVUdZUFaPtnG/+UiwlVwK/2cZaYthalf/dIIoqMPCZP3h5dqQL
KIgVzplBeL9IPOmwkCo7EjaHSG9Vlwr4lzXED/Z87kbBYXeSyF2pGXFgd6pP+kIa
1dKPPo2pVSv9FFJKnXTnIpp+ykoLzBsZlcpmpCfQzl149yrB4A94oL1YGLNxG43x
ISJMCFNfTnGAvdR5W9Q8VB9XjC8isyuoNiJLz1kw3XAQHlhxKZ9Wd9XUyHwlMUja
5VF04qMrr3ucnqU1YDk1szhoayPfKyXDKjLCFFepPER7CYj7dnekWmKHDzb4Uq97
PYeHAmTRKs1EYWU259E9a+jZ0cZtdmOuYQr0kXxjnrF1E+z6Tonypr9LuzOCgAKe
YGv2GxAsmxYXpkkgLHiqY4SMzEzTCa5Es8zEP+z81Jnu/syMF0Cwhhyf+Xnij/LP
xMds4nbSW9a6/sWdD+EhvOs2HBYY9vukuVMZ2QV7oEJpi/UnIkoMGYJSiGw9HqAv
JqFn0N5HcFLVZy0iSGJ1YOdhVulFjSi1UjV5h3Hg5OkxBmPPhy0zvxTTRx0dZ7z6
tQREdq1IjAocw8Y1fu7Q7URUE2UfP0AmGvH/5Chg21hjydX/jR9ZF5WemKik241w
Av9EVueqCSIrwxUMZwKCTu6WY5uHjPAlli9zqJ90VWlH8FGWKrgokD+6o45kEFVS
ahxOTaVNcD0iVkX+aM1MsmSz3qQZxaWuz70M3/zIwmdQrW3BzNUM2gSMI07zmL0Q
Kwco8J8QX+Hd4mT0+ThtIvLwwYZMetoRzkGMujeZvc1/sYSTvxC8tmRiXmxS300S
Cqj+EBxpnQqnBjVzenWKGpdE5bkqi3GlnCQsxVoauq92NNg5TQbBIwwTILAOyouM
mdsF93yVdSS6pe3ZRrCAyVfSadWkkZ86E1AxEV2RMe1o//o0Lx7z4+IMGUXUr8bf
usLWO6YJvYbqvqN+UaapIbbQbDmcs+QnY9pWOhevtlF2Ej37y2rSBa1IsqOfGAFL
RSMY1DWyy9rk/W9a9D3T+MEbpO6x3NM3J9qCRrzSMX97dfgk+MfkHX0+wqgTp/Zf
mxOEayehtT19xu5+5JBfXz770Qkd2SIhGhjK9i6364fpGPKh0HlG2KfP3nVVMmVl
xpxrYPN9LHRK1SkRbv9OEOQ78tGVH1NsUt92Z+2Hg+WtDVb7trT+Y5iYaQpmAefq
nKmvVl0rQHI0IT5/LJlhhL8S23vCwk8nCr6E1M5y61oYD1gZAyOvsrPm4ETmO1bI
+Yu8tc5itU/OzcC4F+SGX5u5i5YhPvQPVLhfXG8318ZAL5yWskhiCSW8hGEyGwHa
eeTZ7kW7YNdcC8OYXiN87/aRK/aQ5fiyPo0wct++eEAcU1eGZaoQ6AzVs2jyfoSx
x38zWXc/QygmcZU8uykUEllU3t1b3DlklRtkjcX3CzWcVBs3U0vPU+sPcO9btjjm
+ZkgP1R5E2NAR4Ary/X5EQXNKjD9XVfOwVdQOr7Ko27UQmfNEFzgxs3zxLI9mal/
ytGnR2BQehkmMJkIE0fuPF1lHX2G3OzWaDd+G+6XtO5Fyytv0RrahOIyRmIfRiUE
CriIN60monGN9NC2a6Q/wM2iN1ZTi7wUXkXgsHGGhoF6dHXvNHekk2P9a8+oZXHA
4dIMNYIZdI6AOPQLiN01m24/5DchLy0cYe+p0vqpaOd1b053RfdMSuQOcANHQoMc
wkeiBAd/HgeRMGQJUj+S9+LKFewxw+/XuXcmvNCXq1t56qlxLBYve4Jw3My8zo3d
UsQL4BMDvov/8zDYQK1slhtqhnbgmC+EFOXeIl9+KSsPnGr1RMmcJGMy6TlRtMno
N4A1t7vm7VnaqLJEBllmpGZB8OXYdba3wZHQaRdS9PlXRLUVtLfjYilDJdTrzPPE
LueSevLB9UjrnDLQvUCGBrOEt2/5YvlmG4cRsy2+RYC0weFg4g4Aof/kBMpWXhF6
0rQVsIo8uhahS0KyvJ0FQ/MGGapLAWYkCEANn9pf3Oq6iJXiguzc334RQNRQvNIC
VFHKiJwpjH8YtJzKtr1paPDUHMUQHfJ59CGtSZ3cpEf+iqE9lNcUGTpaYxQeDyX8
HGAeECTUMDQio266ZJ2P6SMNHK3K6goOkC/RCd5B8zCE0o0PAymULVadLtirVlOW
GDoil1x8CQEKF7JImSqk3Gn11RhPXm+u0mg+K4VRByB0RJUonzc5q12olzXtXBgW
s/fWN7gDpQgzNJTcfLUhgg+wdcEk37HJjFF8lUwLv/t8gxzAPYZVAhAF0jxZw5WD
/0fmTJEU/J1uFLEIafxth7nC48C9FwPVtReE0T3kSUKnhyUQuphZSt3Ng6BaE/uC
bGzGr6UxC7DVj9j9cL/mHdiBtpEW5qabS8aO97qxp85VKUdW0kimhmlrF56AIMZ9
5vDdw1mZu+tk8o02AT3fYF7gcekKwap/T2kgbf8SO+zpIAdxTfsdt83vnpbG0V7a
oIbYNdKD4q9I2m1UQ7xyyeU3RVG3h73RpmKPtcN3tqbioBNKxzlWdWxAVO+9LuT1
7M6q3FXIjcAouQ8kvegQNU5Iu2Mp5R3eGHHopUxQWF/PATXxZGiCdzWazhvoPVvO
VZ2DmDXe1cbgapN8vK56eYmtm/d2IlqbfdckjpG+x1TrHPkJiUukTNqVW8enOs4A
bUUDFuBAZ3LTIdjZm/73Ds9MygfEmMYZc0gvZsBtJ918taItRpmYS9l9Ke5Wn8bg
VWj4/fxdLn1Rb9hOssVyGSxFEYpAbGNK6KhASnVwHsbjQZcTQgkAOtqKsPeeJkR9
iFGJ7q7kuBxMvUJR6fARfMJZ7Wch2GE+TWThrmjEfq62I8ONC5EMT9pcFcZkpX7W
+vBCZE4uiE8+32hPAy8jwD6p97OwQ4GivshFkMzOGCpX5NJD3MPS3rU+RVH3yKXx
tOxwXHrdckp25WJ6c1OcpLZ/73UZosPpf4qxizzcft1yOXgkHQqhIAOxzywiTdKP
eyJXIoluujn6+v2E5di9vwMpJQAPae2HHNUeeDlrP8kaSYIB2Q8515MBQmjrauhd
sv1UyCsuD3v10QmB2066P4S3/7l6vSsIBrrVNtfFhwT0L+Y6QyFz+9P1TeEaqpnj
J+K9ZTuUetZMQM5XAp1EGV+ZLAKBhn0imJrIrqSYYNedkUaXvuwXlD53XxBdriu6
pO78FK98p4kVnQqcRbKn7n9DDMSmIPGZrCTI/ryUrEk+l1gcJPHhMaMzxhmsczEB
W/QZasIXLmPs9/C4dRuiHvCYAlxdswo/6C3BxHqYdGimWDVEOQLNY0lfPRGUwt3U
0CyElOMLQ1XANoIvzWpVsI+bwbDREgRqAEIKbK1fVBjU338nyCErrNcAeCNjuEFC
O2N5XVDh4NAiWfuCku0xCYUmUkMoGAQ3J29f++hAuMz9dRvmaUgkaY4s/gWeDGDf
f6x5Q/UCHhJoAGbpFP6wtV+7YKTAoqLHPagVuTO9jq7FfpAOGofrDLULbtrqx1KQ
q4z1AJQ7bKqOHzqq0QCv3ZeBlZyxAIsa3sGPiw71624s7JmFHGWSONPe8d9iBX40
gUSCcwYLFYJSnDTjwUotqxgesUfP+g8adKQ346oGhgZCHkEH9dlAF+f1J4KJSGRS
bYNIS2BTGZCNTmj1zuinGFl3F3fPLfOpgzW+YimfoquFApYFKcLi3SLck6Y6alYT
++Zub5cPKNX0pWzPlpKR9jjQO3iXzZIpr3gNvyhU0ZvrPEm6OsRj1GbyDC2vudJu
Z0Dbia9tKuDcXqQ996lIgrtDnsn5wb5PWDR14gD6v9aNYsfxLQN7gpLNZOTB868Q
81DGHCGpTYff/YfR1JlulMONC33+vNuw5NkqZKRu+4JMeO2s96W1mQxDC28teQTm
4mX0PkQtiq/KHnt5cj/n9GL8rVP5UJQ4gGyMJtfgFocW5LY1BlQeejtjIIbmdVVV
zWZ19YLZgz7zCfXWkOkKyivx775E4d5ElbKxufMKB16d03BrhU0jQg/C/uHqJ/Zq
O2BeGdK1Qt3sV0Dh42tdSqWaRNg2bi3ZWBDsEBjCYv+4UeghzNOpxYhJpouQslMk
sx1Hize+rJwbMCqNJUI4X1mBQ1Jpa1iXCfrNClgzbNMh+Xqj61/xYXybRuorgQSg
MMDcLzC2NYZbFJ6JK4L5bba0qByhx36AavjNbWrQ7EYPkjWTycPSFW9+gg7mCnDs
RNZsw6DJVQM9Ouqu2yANZaNtpiGWRvqIqw5cJ/mwvQPGi4NHWfLv7FcEsl8kjBCl
1XrhdMl4fAG/Qlr2gO2S0Um6XRyXgYnA/J6BBaTkgKMh/2H3oNGHyh2RV/Zrrz9n
iKabu+ZLeJXyy4lviRQpztangRma0i99Z6/Xc/U72PLtM6U3WgkB9ltA2okIth8s
QdFW98B79TldtgcfgvjRsBySqDTU9nMu16OcCWmwS78o/asM3surfvspoJ4RSp6d
C23l1iT2fIwuvmSo2i/2hyfMb6LxBEcYtxKkgV5/MqN3DVW8wPRuuRoy8hkSFZ+3
54A3P3piEVlXaSYKgvdO0vq1Jon+NOiRy8kfrurkc/CAfCIo73B9+vGaggcR5FbB
Cd7HRcAQwdwbkRBD3T9juMpXYTH7MABIH/8ccflwuDW8GrhX4L6GRimLHgUOEt6P
ZfzV33f8xb71A8U7kqJkwKGfote5d5231I5HTLJz02+7nOunA10Mgdbem2lCZTjF
ZxgCfxydMp+5FAZRrqDk73z3SErSL/tuEsw0bKKrG6cSQHpI1Y1a+b8/24HD1kaD
HSag7IpJidEHDjj9hN3ihV7yom+X8h/zt5TV7MDG8ukYdRC8CTgzSapzbh23mkN3
lQsvdPCVF4Uwx4dUkIBHPK0BouI/EAOFmz/lkw9LXRqi1jLGCUvw1FZEo7IDuAOd
vG1X8VeyD5DyLwV1wIuXRng2/0xhoaCWU+kcPsqypzTuiJ6pjvLrtMv6aEFOf3vs
YStO1FMZ+7ZbbGkYjnIwa49fOwIuOfSC5Uo3EUhI/QAdceaCBQNP6eFWDSpXbeLw
CRjre0bM7c02Z8JwWQit5BXHSqVjyxXqIXhMnGlH5gLFy2vlDumtpf1gfGcGKHPR
8ND4KeMBB5MPAbFkKSipEY1qMvb0mo2oLR8i28QTDtVgxoeOVmLf87C+od1EG3ZN
crxU1ANbBKqMaH4ntW1UzvO1y6mE4i+GlIYB4KJeFbWH69OALzFjnGJeEBziUzNY
zNt5GeHCGsY0PkbRBJQmM7/EIR1rFVSXvUK9svQNumtF+02v8OkcAXP+3ZIdFFpm
MZWuvjCVqjs6lsCjCr+1ygwNJgBSIpxT0YXHAaojrCxrT7THUfHU31tqyFkIbPVH
3Ieww27EqT8LBFK66Ex/ggodneqHqDIcJXkMweNhcPK1NL8t1b04GtEG+Edl2nEI
7T9YjVuLIh0FmYWCkOEneP9h/uimsrcGWzsN3Ho3mmroP69KfOdRQvIgE9mbWubh
CLh/PYHVrH91nqLhCtha6zu27ZnOMk7kgSHW+tR+l0xdG0vTA+pPXcYu78xcWtnU
ebyPljKfjZYzAIWhaam0OJ8GT8rDv8IHFZzRsJw6lNAFWH89syp+h64wFz7FE5iQ
GI1nEzBy/VU8ymvXwFesv43QLLWpzMv07rxYpjx+Lh9RML/uE3/STpds6oKXAukr
F774jjE6qa9cJMzN27FWrIv6fWzt8YhEI+vklJ03wdEwJDjzBqsPqqs7JkpUPxmA
RYJjXmI82dNdLEuxW2fwOyBF2NM4RaLKiGedE3Zyz44mEOj1YAKnfn0uypE3hMop
xAzbkjjdIpcJR4dYkLbADtGyD7sDb2cypMpihHkmGlSXsXzsjxyHlb8F+Ic3Nbit
fal4btbAQ9/rTNkah3sYMzyvfKfbpXeD+WxUZLDL4gJEKt5qfxDtmQ5++1+VKIBy
BlPscyv4boBNsbAitpqXrbmuq7lZ0NqY8Ce0u+iMqtN/ayLyXEQnLVXn+5hmj6XZ
qllQmlwxFNkWV4Gj8pKYwAtyhcK+y3zxIT7g7lJfesEqkQpX/WhLMZBxCMV/L+hY
1AR8WSVU+UOdHP41by07llwxCZOnL20GrvIvDyB6n1tfnKYzJ8O/exrodpLA1W4u
dY7k5++pfJC+yRUS5LbqkrkzW3FHutUsKMUIQ6T1quolPS5YfFWi9qNX22YRhMD4
CZTiyHe2/Nn7qsoQQrSnyHObSoP5wZ3DPdgAU2JaXHg1Om3OGeJIvqMh+wAInGvS
TGYoP7mQik9kxqGaBoJC7QxShGREVOzIQA4jBKYCwumRqPpYjQ8Hmm2nAn23eRzo
dKz8OiojNVnl+nAjlUMxHZmgL5DiXB/YoKJik/9XKZ9UA7fllTie/11lOO217swc
Qo7PzWCYS/dKVyM1bShN46q7YrX8Cn6pFzPbiAEI+RSGKRrhbHGJRZ+q0ZX+ilOk
U7KC8iA08wIY70fPT7iuPYQHS7qZIxuA71pleHRyHienM1Ae4JKWTWLt4wPk3lK0
KsFEhxuTxn8yO0xFbnfIHuApEgk+UsYM6u55nBv3b3DOvL3+avsHwRvg/Hnvc4v+
5mytmrufuPUFUoQEve3iGHndn2wssXAEP/kkaE2huJjayWhSFFpy9F5+zs8yLcSJ
O8S+McKPWBa/GKlzkAOM6B1DaMV6upKG62shjYXJwQS2/w/YfsUXNPtLLmoBfnYP
XNubDSgJORMVCVry8EbNbr7kGAww3MCGcsY+bl3Hy+LdgmHh2yuCEbYOW/98Jbw+
5G/G4yqbNt/IEiN2lrOxlScfMd3nxcKKSXN2eVnxqebJqhm06+pjn7wpsHUfG8+n
Fl4+SMgYytlcalzePf72uaiXE0z+jbiAvU4o2d+kOfOK6GrSYXc6Sw1mZV6ogumG
xN6ERF/no1VzUC1bXVZiIWLDePSkQVx3stfuECOUpimgh/OkdcW82tTT9qnYcKlC
O1MgQraFh4U8Kv3GebZd7W4pJOyO2ovp/1xUpPmYzvFPopmYyy8jQgnHdjwupKjD
Xxu88sVa2WRpsufr9fWHd2aCBHJ4vxe50TrOUp4iNU/mZqkdE8vP0xm5/p5NjpVL
kQCh4w+sm1x2iGQOk0B29mdKzOxyNqL8P+/I9HAwSEYfEUsvJmfK4MvEFRIk1LJ8
pUkX5lZGoc7ZMq9nPa4nIPNY2Tr3DJDXYLZd2oEPoi7REW+FvrgtKIWS17FdRZoc
mS/XSPqBXLCXPeCTIkBJr6B2bpbFeWKnU753YiRjEfmwZ02zDizvNZ3QwFR88q0s
SSirM0aJp3ji10BsyDPlZglqx2TItwgXseAhQRFhQ/pC7pllba/DzR+FyacyH2vo
i583+HY9IRP6SYc7nJ0E5v0TTcPSW0WQyNFOQ3I/biElp2aO4l+madAvlHbKVKDr
jTaFfQ17qiC88YGCv6Gdk4VpnFPO18CaVbPc/9PnbatBiFntjwcESOzvnVfA41NL
yh1s3b+gTz/XZtJH6kxRGyQRVGYTfaDcEdQRgYY+5kmPdzR/AfqUgaUd6te/7GyI
ZSeXZFv8nalsWXOlORtsX3+v2BSpQpZPArZw2GSZfTVc7h2XFkTkEVWS0aeD6qBd
QkHiPScPfUBZtHIgorX4w4ucMmEzdTInLx5KMfxLGRlyI58Z8kvivuZufbOvec3c
+o7UcLeoGTltgJkouLTzcP+AjdbbohicUlC/A3WYRn7IsFHmh3PBqW+WktOWWpBP
KgIhuZUzWSIwcEEF1av4W4num+0V9IySpyshFRbCEBEC6ozmQUfsm76fOSaXomqB
wy4secCuwHbfWhgrjV1DXrmbnFuaht4EXcJDgIbwh0mwa5zB+ENUHUJ7RP0rWvOE
WrBlNO/1+tRZejLi+o2c2DVNz93NCZHRAMtaojiLvljGoTAcI12s5ET8oTEj5EZt
0HS2wZUIP/X7hLj8TPpHQ2if8xzNMzPeFslAY/AKChDLmPv2jeRvQjFW4E6nLuoc
VrVjw8jYQ/TNrrnxCttzdDUyKHVlXY+q8SNtD/iIQezgkN1kTHmIaCPwB3VZkSby
L7cHy1pzhWNY6gZBJz4gk80YXOPWlXk70tJyL6NrfR6HMe61+8/qqzfXWnWeGpHQ
0H6ksah/cvd3/OZOOZIs2sgytPyxDRRTYpHg5wX8qG2vytW3xv1EbYvSjkkRgSao
A4gC7t+Qvk6UdgGjmkNdeAzGDVqDg+i9pj/Ln5EuelAMK6apIRYkhsj0PGnna8Hj
PIcEDhsCHWI4B38BfrjosWs/tKHQQtOLkh/lv6MasKIjjBzbd2lfIPpya85tMzzC
liAut3d9+kBUXY9milaNHrB4YkXqv/O18vPkN0WygqIMFPgrpv3HYsrKhbVoCOMI
Jw81peFWaxh5QIuJP0d3IVHvi+yiq6wY8O5agvPvxQZE2P56yQbW129hr/AW0BgZ
jZudxziHiRgWrYn4TES5UhX7zPxGhEUdSSd5MXbx0zrVLbxv/al4Y/3Y93aK3nEM
2EBBcqKivtlLMlyKS0jIMAcKZYRav5OYW5UzWTeNYFLFNLjcz8glX4oA/+YWrt5L
dwE1cSn/UeqlakBy0nNfoM3IMj8piPMLEJTnSkpqB/KRmLUql/zlnKd3mFzPS8cZ
nG6ns3nG6DMlF4tMh6CjUoagZLN7kHy9W7DyuRAoKXs7Jqx6hd4WMkZVyz4w64Mu
/g9Sx2myd8G4T0IMuGEVx9RdmwdL+6BySFstv59lHZEhMrzCIxrz83rJvSnWzXKq
xiyEaBj8jqWb+yMweGICyyzUolqbbp5fc9eqxXBUnyMWZcvVZImysUtwPucPkEEG
hAiQxffeKZ9IN+50Bh02KWDRWUJ0wHJ4mWz6RB4lxmmkF1xrDIq7p7tIkgg7T1ef
b/p4KHmCYlV2BumvZYdgHYQmFswsO9hpILXmUhaSQnRUhjQo44Ldp50VdvoJbYAS
Ry5e0pWR6VLRCEhh+/HNj7ZDH0TyBPj6/yZeQUCSWrqkkZC5Ncs/pcVDn8wSzISM
KKEAtpkn9qg9B5Uw+PiUl6AWxkSSK93jxI683RwtR4OQP9c730J8eO71InMjDJ06
OgqT6UieSOCi0tl+cmQovKrAidEPhfkPuTpeIgt7SzxLazQXAOW2brhZGNeJFnQI
Awboyy5JCHMMLenh6YpPKKeiDQ0d/+sOMHHxwtx/2GxiWOTg1AECav9sWYJ96b8T
WV/cKLy8ZgVkZaKr3LJsGrKx4E5mOw8mWju5timYa5bAsR3dMYyYpIypcWQwUt59
CAoac+cIkokyWIy3hpbPcS2sNSNXkBRgIrg9ZFBf0mXxpD/tLHPFbNBgJlJWN+vy
rT4r4+SAozVaWnNxcK50pid85trybhqsQh4jTII6Okgyu+g+TNpEDMK8Sl9ZxT/1
KqTwErxITXgNJ0M7PVhj0ifbK2VEIFib3SzLGIxLXwloHSpV4zh4ve8erExWD/Gy
HTSbaVJ/9PJPQRj0KQEeTS/Dbdt7rpug8FikfHg6Cg5SoAE/AkjKRx4GM+gxy4S7
hvFP56qeeesFDOERwjvGIkD90m05CC2dgvs/xzbEMV8OzmoCQzfFvWJMyFYLBwDZ
HJnPThJcTSDTsoSODmZFZPNt4pRKTw9npqqj5DSjueuYcW6Hh7Sa26a6qa5w1O53
ETI6bewnWKm48HAm9dhDMztFludiCiFrkFPmzIllAkgOGw14b01HPMdoI92dfAgs
VzQFk77n2M/HodWoB1nJqahwJUx9LjKahm8UK+wSWn7oHASZTswa+I3g5Mc2syuD
6vettbs/DcyoeKocwXOZpQSBH+knBzvDtARLupV0bOfWMHPcSb0z5mVvB8B987Jl
QboosyYJUbVrIqwO+CHkuvQqrjVG8QeNK8uHzTQEquKS3zD4wUKVJhmum4gfNXYy
Pmmm7VsFTYAKH7p5AYCrCct5QMtd5sU3vO6zjP7qji7yUYObMQ48lnsqW1njENgh
wNoWHn3X4wr9g5YF9GFqK47ciiXcGspHb2/uI6/ZkRAcowdgDEAVPYjDZ6C6MyY8
juGjQ7Wbo0pfZqbTB+Od88hfK8ujv34PX9MFHY8HMKbUxrxWXRog3NtigMp3zxif
Seo/h4Adsczy7v7GZH2/CCkEm0oP/8cyPtnk3w6LJwz6G856rFhM778e8UFSdo/Z
bvdmClGVwoKLII/9KBvFM/juxwCONvjihFdiw0R5jII2Vk70CeE/uf1Bvvuc6daU
KD42W2nn6HZeMg3N3/CnFX62y2uK5SJFG3oQ0ww4jAFlA6q5KnV1SOtDt04fRbNM
7GYMYTAg1rfC5l9FEtqYLEJyx46OtBTNXfzJCYctxgv1A7OXf1SzeNxRGKPffZCd
DC6kMWQTt58ipe4jbdVRGNlF5h3KdQLCshs50zVFmTKpHGlNgF8KzTpDRu8wbc3p
hu5UjpJafapI/1x12fnUqGxE2I3xh07LWq5wyYYoHA0dIlZULTxh05ZQ90WiuRn7
kHYU1Wjskr3nD102/r63n750C5cPSotvQSXrVx8leKGBHWIDpaZtpxhlxknOwZSo
MnWj80lfz4/tiQnzvgD149XJQJavfyNajrRDK3Jk48/3pzZx8P0fsLHMaO0yxRRc
SE0E1UkjJXZkGpP57PuqhAmrD8b1kmG2tQWTG1JZ1ADw3EI2Wvi5AuQ/6LESpm/F
wApD3mt3dzbKyptERPJpUlfD4sdrEhMhaqyrEKCcEu0Pv95tnM3szMaOuILdW0WF
f7kV7Il+4JeyywLI32bA3L4LEdS3T9UEqGLddWtaNjefP8pbi6NUOJGAmDwlwbgg
evX2q6x4U/83RNuFkexZD870W3oRS7En2p7GZfAgzMcZNe9Iz/bJP8sh0gJKVjPl
cFwatvYqIRP7lJ5cXaFpagWmmuQ3OIz9LywGi3M4Gi695jL+twY4/NGGpiMysLyF
j7PfTFRYmvif4hMulnzF5rf0+hK5GQ7ZgIhdMyUcFyiyj2fTn9y5H2/lrqnzvzn/
klZ8ap44FZkga2zntk9nZi0D+Zzj7azUJ5a78/HNGSt5/d77+6FjcnpU9tc6p38Z
/TaSC1yQjTDH9dbn03QE1uiu1iDMm3+eFAfAOAr4TtbIDxkulkgy1TT6eH3VoIHP
d5fep4DOX/pea1FeSg1ZnoL064eM90faO8+GCtpZn3O8ypDT+TxxsfzLqYNIO+k3
7I3kA44GYikzQKYIdJzpZm6aikViqJ/gXnuE9ZFw2TT7oVl4FD4ba5OxoP06dCY3
jSbnq+Q7wPbVsJBn6m1NU6aZRhH5/5lvrLBPXNIKwDYprOeHYzBplwpFGp/ApNHJ
n6o7h9V9nKwYiObOw2rGkMV0rOdSI1e+MB04tmoscEmNLgMNfejNLbErstx2/W+Y
PaZlPpxTB1TVTUv0QBOoZ9/I0CbxP42gwMFyLZriU2PVmoIwnaEi8I4qQyJ4lSNT
O1OXK8RhBawVbzA5NEg01+kCdZxXZNTMd8obpbOltrvbDIITaAtTR3ylNz8h+UNQ
sJx3u/hrwrgJMbwF4FgyiB0LctdP9lGCSQCY5FWI5fgOIIsd9qDWgg/bFb/o9kqE
ixQEV1t1NT8NMgRjg7ajEFj4R0fGrZbZ8wEUItv5eO9SP+UJh5gmoaSSP9/WgmlB
7BRZcHOLrIOYRijeekj47V/7Gfn3cx1r/7tFS+pNklX/Chj9Zs3gPZKwepKRv6LS
HmXm1FMRNkO7WAUiB7gXfcBMboGgh8XuT+x3QzG/ZHbJiF0Yy/D3t4P7mVfvt2uZ
MJzyEw5jzmpll/tFxh7SoNOn/4TVKVujXhDBU7SmnPgguDN70ixZkFrcNRdLVAeb
vv0AQseKm9pkf0cLnyJTQw2VeOynrjmxd+jbxvp5PWdFQe/g/pK/WDjcXYEgXZQ3
Je1yo++PDIFlkOnVCT0gas8XgyEkhx3b+tJh8z+QTnrpHSz/vwPr8docWYGNBqsW
RyCfoFPabnNvEsWL2wxrhUA5vixIVveizHlmppX/CMoGzFIhAbNzDqYgc4hfBQ+b
uA2A0DcroOgG82NrPV1Ly1TQKxocvKo2YrOBdOuEbyr5TkGf8TrMGpJerFl2HAkn
DZvm1KvgdGDC330mSIwa9keid4jFCYcZ8jO+PxzJIg5was99MFHLhP4nNH9/LKJQ
9QTlOOz2fJ9gDRF/qh4pyThQ5AhW+ThDxLqyrzhUvjqzdtAq3iAqS4dOozTMbeIs
cyiSfgUls7c/k5LxFd6GX5CUKhUJFdVn6J21JTOlgo7NQ+Cz58EhW/qYxPJ9ln/P
BfLgka3pgZksw/gStJHl7YCclWyO/E2t1asISC+rfEi5P5ZLzGYnA7y6pEWAYgIY
sDbbViAWpfFXwrCLv0x6NpjXJtroXyOybUARKQ25Dh2732GowaqXNb1BGYc7MSoV
XuAzSDTgFYoI8x6Je0AqUF4IcX/te4P/BSpc48qbvI4QpJTmwg1XGya8QM7E+8TM
s9Mw5Y/I8tim6x9EmQz/B05h+efZfaO30DMcT2bxG7ehUOnNRTamNA9TF8JvHxud
`protect END_PROTECTED
