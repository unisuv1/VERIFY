`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
K8lxmo8jjtbkq+yGitiehB5O9RTfa0LOWVmcrF78xZb3hg1f2x/X4E2l23UPobhg
m7vmqRUg38t9UoiemnSXCGdAHT3QEzDdKhlqM3QBKR4684JIsLi6MP6OwwUZ8+Dj
rPveR1imIzknpnUtzz70x8t3tKIeaZweieHWR8R5qaV44OM8wxih7DoX7VzEl/j7
F01k1WV7jVktHrbLONHYU5+kk+QT60bVKAuema/w8BiilmVyY0dBB98iMldXSAUB
EcQ0cj5ckiZnq5rt73db5dQP0rEqGkENW65Nl1qyKMH4BUwqrF1vKCO5tcQ10Ik6
lVmyYgkjr4nNpoFbnuPROsJj5pa0QDp0GtdSNoC8C3zHVJLUzD9oDR9iT1WiO3cG
2uZyuFhrbWk0bQVJwd7erTO6M7XMsTd0TTozyjZbx+u9Hm+shwI81VV9hLV4Dz8B
1xGhMKrUh+bKCpQe+p18pvXZMaSS0ZN0RiOODa7MUv7bUpie/PB3ygaauClC/aLA
IAl1Aj7wv3xFhbcpYLHsEKdfvEn8LXpIrOEjZuEZuW1b0J3VYDV23VaCL9Q9hj5n
Z2W0M6fbrbwcwL3TbzZhq6itarD1OzxFLwC6xOQ6CcODYxOexXsfjvqYKzxrnPW2
o2ezAZNYLbrQyEd54LrNdye4OE3WdFzunwLMKU3DF+eGMB99JTVlhXvWjFifkXvR
LxI7QRTs9zyZDtKEzlCR6Yq0Ktu+1tz+f5zi5tNXrhilnpYV2jl30g2/ET0sjYpL
r2kW5+XwLBR8oUXfY3/YfMP+hp+Ctlydaoq3LjrpJpI57iIHr4jVuwQgVcmA7iGo
P2c+j9bKWfDcsQXdSSL6ECv93ctiH7GMAdbKvcYgxrCha5iotfYu9XMmURIiaFK4
sOe6dre50gddynZ7PonxGee8X5QAclT/VOwfovOXY1BlcWNSL1nryV4VeYgV6kxp
3haRA7R3zwXQvH36QNQ7n2wQwlqpcJgzdQ9o545j/v1qrMrsuss3HsXYKycm5K9h
d6PPVVqyAI3UoBaLwL+bVPxANZf86jj00g5k+Z8px2ngXVocZL4tVY9JbisDAPEy
xWPeFglstBlyGYT/qOwxO2bgOPff3cUuIIXgePAWV7H9i5Ob5fDBenYpw4VfBUxa
mlyVLXZgqiPDTO6YllDvZ54Y0FZdYQxOBDRYCeiq2ZaZmsRdbJbBq6rOegQQAcxr
Q6+qLhPRAD+QaLbD1VRu774CXB3EwDTJ0sXv7GlhqL5kyabL0IKclKpVXlBlMDse
sZfU6yjaU7fXEFopSG3NPQZ9KTlQFIpWh7iQbXztBqyTtSSjMIlIRE8GbyyUrcvx
9ktCeWCgFApLIjFiZkxbswG7C4eNA0RUIxQGjaG1486hKA/jA/rtd1bxMWhZrhK7
ehnK2d3vLpIi7IUMVqop4950sIWkVN0g38Ap1+Jb5Pn7A9mDqI8x0HUWM0mpkDdw
cjuLtDUa4nomVseFGkp//Xcod4wPWCN/k/sKg7OdnEaySsRntGTT3EHH46k4/AcC
1LetczOOAOAO1X5mXhqULAzbBpj6RGYc3O1f6+1VrGR52BhoMT5TgGOK16kkjNNg
TEun57GCezYPLZyMQ/jBrXZBp+Ny1n8AKMRO/a6ZrlDIY70RRxc42iz6JheAs4XN
eWq2QPMKiyyll9i2LDJ0w2N0udGEJjoU+Km1vcbkxpWCZ8oeRM28s4asYJyQIrPY
LcgGvRhVI692qRgFe9ErFhTozXDtCT5rVGfbuQcHaYkV8ew48XTnzf/Tz5bF3Axa
JvnIgzCvr3qa3gNsAlWFs/WCdxOQPUsHifHnuccT/G22ex5truGrOyXJ+jcAlgCG
6riYdEmVKwO3xKVAksyIXfKCVPi0JZj5XQ7Adi1BUcNRhXT+iPuz1JHGFtlv/nmA
GMxkFgQ0Ph7aSO2v/iyZfHI2cn730MdSEgMYiPHxIkVibLcc6n4qMfbkFzk29gBk
smLzVOL8Jd4WI6dRJLyxmcV04itweRbndA9h9Om4MA+gEi8AHkoYDdaPZuj6qo3l
gi1J9ASBXfowV6K0IJuqgGIoYUcbd4ePx+xBcDvlsMvp72P/UFqAWUFg+WcpFhaZ
CiXcEey9pmA7oTeJY0lO/cy7nuCJhwY12gExnG0KH7enyYRAP0iMrcv04/Fj7/V9
q2SQSj2jnWJGgfUtlwWQXmqy4H7acbEH2ato4yErqXCQiQSKpGqiCaXIgZ4Of2bQ
zUS/x8AZaerHD9QO0b4w+2+CHdv0pTHqUoSd9bKlvMNgSGSP5s15Zdpwj3ox6bjI
fCpsuTLeyMKBUBT6FxPHKavu3fv/Fh2/gG2DFuVi9Ipi7K9oa+eEJ4hrRuJpgHPs
XjtZP9Ksb6gM98ZQwyGk0w3yD7kyon9FExvJu6irEYtxbiHLDh53sX1yhS/gyNUR
lgxloPS7Lr0yvekZyfAJUUDyyvmydBCAanaqdtLnFavmvXS01QAbIP22Ubv6OfCO
uL006GyLUp47Zm+wgpJ7iXR4B7v9RwW1K2Wyz2Rmlb/+0Ti4zbSDHX5lvACQxvbz
IaEgiaqNOeW+b1lII96RmQHy+uZowpm6t7qYgrU/UdWJAUYecgxGyFQ0Iodzmcqr
ZFQB6pxGUoGxaeicq9FI9vFlA8i7OKDr9XcD5uil9+5B8W4tckILysATizm3xVV6
1wbaoRHrsEMqJ/i/JvzaZS/196qjjuHO3XO2YjRh97Ff26QAP34K0dSDKwQqkdGv
RB6x7AR1jazwUri1Ym2kfsIFAyt83Daimws2ZEWSnLVKAVa/7JKZ+EqmFlzALNo6
+Pej2+PPjXU2LtnXIQ8DYyQcc32e1Y56Fh3NWUt92ZQxAwXMTN5yTtYiYQ7EOhmK
sixSER/c+Wq9UmgCeuSYoeqjL0qXUhzTH655B3Cy1id457gt+fiSF6oQJQfT8lXq
1vHxJwe+3Wu4EB9Y8MJ/bVddQ19epHI2j5ZESuaCsQ4syeLfw8bDT3Lz0VzK4PkQ
leofbk3KDgsdy80vZAvpk6wY9GOFh/3sSjliTKGzSi0ON8oWoRO951T7H2wJ6ck1
/KbO+boLcIYrBTf8qKz4Q7EVvU/6pBoecq/WXf4yh7bLr+USy0aUTvSQfY4uFSXW
1jQvWxOurfkENg7JsXzHlpfSdTz5kf7HWWvjGW0ulO8WdtK+x4IkoOiXcnXMzdjf
156TOoyhWBbNH8DDjjOaZRlgS/aFLqoUnBcUr/sQTObTt4mlEXmKVXFBRcletdI4
Wp7axmGs5nAXjqebS2n1ostLJ4iKFUCvuq5eXM6P8oVw3OmsypwrXRZgdc+dxNfT
fTaIFUfaDP60u8WIeBQR0+ow5c5m1xrYNYPruMqS/uqwtMJaGrp3Fm+e/lopmpnu
OGGxOO5wM00dXLYns3J1xJp2O7pqM7PokWaTOazxYxUgDGnf8SCLCYppXwTOAdoq
JpBRCOcSQP0Yl5vQPL3FMUCjesktVqHGqkbFoMGYMsd1eXWV3cUXk5BC+EIkbGdg
VSDU15bTmGNuZy0sHwjN8yxGF1xf/J+bX17CpL72g7U/SGgylj4gi4fP0sQ+C/sV
DJC/jrMI5zQPdVFmLHCSVOjDFLTyq0So703zs3LYqqL8DborNO3OT3FW37FOL41T
y+G4of551RjZrMrAaMT6DfvU3wDTPastDokjglFWOKr9Tw8i+0qOJ9OFvaONpSMM
FJN8+ZMVjpWbU7Bi3s8ZAzLCM9XdV7Cc0YgdlUO0NWo13MNZ0S5cPYd+ztPqjoaa
ES86NNjUkgS1Gwf4KeE8XImX3MbVSHlQ+79LrSWlsZ5h+zcC/4zGMQVt5gGrN563
0U5+vaormGUlhQf1GopbYeVUtWnti8aK+hxRXBDFMtzjeS9axkNYsHaF2oeHzipg
KzNp2MLFmDGE0QdP7zxkdFGPit4cxWwDIRiOAbaXwoRHcn2aNtTiiBqVHaT4r4St
j/k5vgRFZUbq8Z+nSpW0RWwNxgG9WPjOw9xTZJ59UCetyDSrtqDqvX2UmJy2nd6a
+jtz7XQBWuHP1Ld7Yao7iAwdMjJS3cq9SwnbZK3e16Ksoa/Ns0Na0NJITSJtauZ9
JE7D/RtxJj7I+1qxT1ILB1oQ6Xmr6aBkzYdOieQ0JBWp6pEhAetjxLdr25ZxOxIC
otc46aOHZyhtvG3lz5usSh4pjUhgRBso/eiV9NAIVtCTZPBn1/SBy22lO6gS8L7Y
nWdGSqWuiCP9fUxteteSq4E6uSosuhxt+JHxmwH3rxRUuHy24MGzmn83Uuz1Ijah
lwH5NAfU7CcdjOa/JxumeW+dk1T/IvCGGa50oF2zux0j/6nttJbDZvypdE8gEDnT
MGPcT3OLUyS8uI8/Y0Hs1xRYaUsfpuP0sX4OQF13/6TCCI5nusX64DTqLMaD9M5p
6IDdaoUFEu6Tzjn+DKe7xEKJHQvKeVu6Itgptqr62WNEnlrAb3OXvjQGT0KgasQD
3tQoVM+2At2gGf3uDBNv4mdS4Azq1a/9hHGEG5SUpQpy0Ost+bBvG0kElOYY5mht
X956JmDhQlX6lm7TKU27b7MClVO5QF7/bNR2MQnZV+96uoFlBal6dAYF6CxloxPv
uswUaVJRpeuVJYC2OklyEZI8fpo5SKOZVknOwV/vE8P4SXJRzfCBEgiOb244Xa9N
sbPFNtKFaDYrtO8f2dv+WUI6jaNj6uIUl7vN7SMkAWciXtE0QPfsgo4JJLWvvoJA
eN0UPGqhM0K2oJx52eHK/7x7wundgKga+zbmVGJ5kkyC0VYMmGyk1IppePxt89r2
0NK4/UQhikIMS9CkyeA5fcGQfzbSgin2w63SltM8YfTMXQxEAa7U5XcPgcVMaJJu
8WYdYfu6eAGNikcWj32o/TTDrNGVQqQrP8PK7BmkYMfi/hH2mTx1nh3PTVWLD1kc
3A1xUYtszKIO4F5j6RTuoUaN01zQJi7h24REySIFo8sn4JyedFJfm+8xE5ejS3GM
ELXZZ7RXS+2pNWGYiivnsbEGW+8DnQeEVvKx4MX/NdrxGCMFkDjhYOyfJHwRtEe0
9SkSIZ6Ds3sAyr6QneSfYZt513SjjNj2d4f4hWkvYZsomFMahRibf7G0e4fckY8k
eKGqr35r5pKdBhd9MUYwH/mU3xSFfVsi3MzCMwmjDFAi3Dggkj9YSWRRqSkiehMD
RLpIiVjl+x4DBCwObJBk4RX8VWIq4FB4TyoCAA6zXFwmvJNxUqpmZkq34ZCyPoyG
1Xr9hPXogXenpNvJU/7ke1BSmcwYi3YMMP1bokSrNF2pd+LfrFxnk8QRF9PR3OOV
WP9KG8ANgqtCNJWwm1+jTTxQO8PQg2FVA9RPdyDvNdRveHOiAGwshKP8vtK+v+ND
81gB/rDL2t/BN63OMk0lkpDqjz2dwOKx66fi3rcRTQZImaaR+vgbNGf2fE8uiykM
OtJoEkykypNV+ZaILdjiJJQqT5SONoVtktYYsqTr2Sq/0OcGiJlkQ3gIr8OYj4m1
Ec+p+96c1h0D1OI+2NISfzBTe2V3KG+tfpCvuYLpaBvk/kEGFphm7EyaepODAWTl
qq087Ut26AIkDgmEZzAfrsPgmXlnm7R0fRrS1w/jIunzLGlCm3r9W09JaUylNUax
v+xgZwTc8D7RVs/4382LDXruuoTa2s2fSUtefwBtW/UT3qkLwFfi65vrOPdwl4Uf
t957UGK+VKimGHAHNGpLZyuAr422iMZq8FbYz6HKCcxNt2mipF2C9cGy/fLi+O6E
NJpt/Lbb2FfL3oUBVt85V0GhuwFNh/yZqHkX3KJ9cd1ucs33XoHqleZFDjrkZ/Ft
2vEOdhm6FNyBRq6Xz0LqMQWx8gZrBi0u/ir0Hel3VZHe8F+jh3tLg+PbLtkP7KL2
HyN+UbvsnuCy4fMA45zmj4L8nMpF3JJItXpCDFoNhmOy+kV4/djwXfvaulsncmbn
vqGJl6Kf/cDNbe5qfevmceUUmD7DWbnvulpwVEIE3b+gn+jMNQQ5mh4uh1Qw3rIi
22jO2/2yPkBcSqmrnlmjjZTOxOPAC4H+ZFSvkAOmQMyncE02EOwr6pvBtDdJhaGz
1fmJm1Vlj+aDxBEBjg6NtY6o9Hpb58yROB3EAPLLWnPKeZLwfFHzJEp38OYPl6yV
/G97LIdkYKBnMQOUt4coUpI/4IJ/r4SSYxYEwmNZ2/GyCcGBvevDJqJs4WVxlpUr
cCd5ghOezy6UUZlevj6j1Ylha1wIqxkO/7cgeOqSh8BcPUTIuKPUcA32JABj18io
mHuDuFmR1gNEAGpjYnGVVbY0oTvrWXGN83ZuebLL6YPY2O7i+Mkt/pjrLmgbgKNC
V/VEI5FuLFCspf1thfaWwRHdnE8A0CNDPUOuV/SFqzNm6FeubLSs3ai1uo+RbLUC
/tWTxE1FGzZFR/3L6GMwL4rwy4CeJJHv78HgSyZ0jm9JzXmwSzOnRr1UV83dDcR6
PhpRbRB5qwEVs5oa9/IFWNzy1cAlw20Ik1/CIUXe6oIviwFfBVA6v5GVj/QiYNhD
Gd0sbDg1FLWgf7QmMf5Vz9k0RzWpCA2rD6KX8vk/h814UOefDlr983Wey1Hn0Lt+
xx8YUS8tyxD+wSQwikjNIBPHXNJnJMZrJv8eBP1aNVYYIA08u47hJLPu568Yfwgm
2SzsLa40AqhwL51btRF6BkBysllFKH4nqRHizVMDMg7Z5f53okb+gS0et0fabgmG
SURXbO6kQA/FlQg0cdxTs9ejRp83iVBfZDroVwUPBWoZli2Hj6oeuS2KM0hXWCWo
PJiSH5P5QQGBcRCOBsoVpBhpsN9RPgMMxjm/B6+NiRKI0IamYYf+4iWQhGLFfIoq
a36BxiX8W5E81oPcXx2tyOD+wFltOnElDtOIRZnoEEtUG0lU4VTmesk/u7mySjXQ
dIM3y4q3k2+iMhVv8/d0ZuIXtoaf5Q0D4Rl2ruLsNvj/wO+G8TqHlr1UfvpZbLHr
i29FFt61RsO8wDuujng5g1RZZevq1PUO+tK42L+iyYW4Wtl82t9vA/cEtKK1ChLs
Lbv0ZveEeJe9d9RakWyhY4RGNpXKWWke0dpklYYvVmS6QMBglikNE+yICVOmyjv1
dRfKwNEQCIJXwXq1Y8pw50FxLZ7b/GrWWftvVwsseI7xOQ+YlQqh5z5lLx2eJCzZ
toL/h4P3ZRBgV0FCUeyBZ22COEqWbcNYhR33WhOJKmWP70/IbQFtW2wCNlf1WevW
s/huapGPEX0LQVTBOWQRa7bBNKVIZ53ah42pmFXJiMHpJ9lVIIYGnsdwLr3ywf8s
ZfS7qoksU7sF/gzTv4daV9HgumPyzXsBi3BEM05oIQ2k5yanoYlzaTR4Gon9Zauz
3nR5/nqIcOcOHy5VUm7C7I8AVxNVkEWacDX49gnoTQJ7R/BF9AVZzLr2uFHgVNTx
WSRZjpKoG7Fs1CHIgoW+Mgt3EqN7DwhJFHjPGfZxk4aFSSSnypkqGxPjmHeOsvp4
3RZLrTUvOi4VPFpNb4p3gxANFJCE2e67YITDVpOvvLcYCxGMscpwuvt4ZvEHrn72
6QBBtyXtnwgG66y8Yth2kt6hs8HCz5cVdF1KOz0cnd1Aa4R2w3LB2iPVLFzPn4S1
X+7wvpttrLlQITNVMF4IaaMVQYQw6gG+ifqWXRocWEOVFO5Vf1m9JX5C/9TGt8uz
2in4/HBMmxArW9ffUwm233IhrAnCuVhyKKb0QVyuhEzepcIQk3B+B2qq7rhAnRF3
UKl/48xqEkS3rIO0ig9nQguR0+801oQA2lN33pc0oA5/yCNoo3NKdcknWx5MM7zR
qbY/xq5ZQIUrKQgasrFXKyYs/i8gYEROhh5C/iyFmthqEsikEfEY4AV1D6fzs5kz
HlQi7YrUA6vGFY7ZU8nD30qHADGqGs3fgFNMmVcng07PiYY0ZeYKFfS6q30tvzCr
73XE+uVRwSaHELiyYWfJ2hkX5AVQXsf+BPcMG2h+W0KZM+BEQDK8MeGN7/ta8j/p
fgrh2R7KaQueelwc3vCLXmQwOfKgrVL8vBBvb5LuNKLvw/CSQ2T7MYqwrhiy7yR4
jVL9YUXPz0d+NVgoCjamArNmcFCXlGkZ2w0bDzQOGYd5WbdgykAxY6D+ccd7jeeD
ub3wtcXUlIhvrbiyZ0ri+/JPNHAqfLiMkQXiOJ9+VE2+dIam+yYEDJW29unCaI7B
h+gPDPadstAUoYagKL74FdXfkY6T3fLuOOJg15T2yaNPZM11lhBVaZJHVIT6P8z3
5/ElG3EPAASpYOMPCAez7x9v+cnHClCKwYowMKS57JEzTpY4rL9jrmxT/Ps30Duy
RAzvYek3XTXRSm5ASEe2rABkh8J/fNIrJSKwbCI3rnGhidbMzio1jeWEaocTkCfF
/pl/ZA12JOFYrrYXWHMeVXfZ2TExaV2JNRhkVO6leGFwl+fAxTHYus0XwdIIL+KQ
uvTl9YMFFjzpiiEdM+AU+fmVepXrEm7X6Ga+u8aC9kp3MCcoGykDfPqms9rhlNBv
55XrzXswuu8h4wC2W3eiX6IgxF/dbdOyjk33x+sg5cFTDnQTQZcSL3bAtI3jMGNV
WH052HuI8V/K3L3/LHwkcM1HtOEfGoIgi0J/MlIW1jNsnuzD/Nn0NtXKwJ9Iwbig
2f/1F0PkHlBjhkhT33Z6SahbTr2FonvRo7SCz662TBYCVGiBO8Mvn4F3/MXyAHKI
GoqnT/m7qpsPbmQ4dbSsmRhxlCRtMjYVLv6PL09S5vLWVDt0W//eMzZrvwMVKUu6
rIjoQPH0rU3Gngt8reBKU96snbAQTDrM6YYhF8n40sFpJXkGVRxVUq4GIng5jTff
RI2CGziyW8XMkGKfkIuT6TxsX5MA9crBJaiNsOD9ZBozi336epbA9Nkj3N+c17iQ
JDkNUcJuN21gVlSv3sqk9JQXaUdcTpm2N0dCZnqCRiIRGud0OgArq9nRpXilCH6W
4tZ6VqYi+dcLDwb5VQoMgSviQ7r8Uj5//IzWm8M5Xh9ZUPDGaiBMvq4hp4NLzM/+
ovlqeJo6b1bHvjSzEC2vwHrgoaniOZ1Dh1SCN/rL2kTYIFqg3D/GhDXz8DNYiAYR
Pu7MDwJhP4WgFudXYBtWJGxoGRDdKRQuGXs55DriRiJJOlJJK+Fvp9kuPiqjV16d
Qj5FTB8ahp9BIbCP0mz+1omMDKWPFYOO+3LV+gswg06o55AKsOMf0L/y3EUSLikk
kB5wgxFlSH83htmwF1oRY644OoRwJfTIFTp9YEvh0lIRPjNIS8R6/fuejeSp442T
abcyM/Fc8e5TUU3oAS+8xcssi0ZDEJ2O9ttYzjvHzNrBEm/RpwfMoltvdqnGmJ2i
DoInLYdg0yN4OS2kAd7iVeI1aM6c4zjQllqz9SMyAQWNRVdTlVwOAenVx8B4n3pR
KQYriU1RPWvL0snGAS8SGL3XCozUztBn80EVeuzM6SCsv3I5LSwwXlBXAEU3BdPH
8pQUH6QxeoPEPr9WRgstXXmOJsfRR7qbE8tQx8SDaG6g714XX4E/pkdBkrhDPnSg
sWQXq3TKpPOLJD8bDLlen19ygBfY8iEApEyK9UytNKHMkN8Ydv4rijo2WJ/mjyEZ
SHRNNWZUeqxzG3OutDK8qyjiUHQ+jhWFRlyWZovKVKkfNds09K3EmyJZS+tiVzM4
cuoFpg6WpRccyGI+52AbkEIN6kv/ZEP9c2F5f8333mAmSWLKoXTOb5y/IIwhgjAY
HlkAZaRIfFMF+FyQlR0UEG+qy2tlsFtw8Tvm9cL7tFFmS4O3biHAXjo0HFy5iP8K
I0ak7gi1v0BEKpE74WnpC3dwOBl9ug1hHhTqbN7KY0F+cwCSODf8L/VQvAQY3vCr
TZW6MWT43qm0Mi8bQ4V9ajmIVRkbXgrVpKw7LDOC/Gq3xO0NLKzDBw76k6ekV2lR
/4GaXqyueV+MYsE84/0bFRFVNnrzxOoO+qOIA9q28VNMOPBOSmlT9BEbp/TmJ8rO
2cVYJe4mgH6YajMlsgKS6oM68vonV+3lMuP6n9139KQcfsTAwc+TCihXvw0+giMb
9+4NmWB/OuMdbL7zi8IulG1fSTnrpZ2tm+m2Hqrwzv78N7OGd3nJxnQzbtU2vaQ+
W3Sm+0LshcDt/aqLkbWdn693STKD8vqvZbIEViBeUGjx0VBVl6NprP4T9n59Ra3Z
k5OEFkoaySgENFvEdLo/EA32hhYQVMjmXwLpwEE+b9zc9RJc2jbDaSI7Lg1fINb4
C0knTAw3GF8xQVgYCIQuUC2qJn9bwJEHky3wnDcPZ5lU0gonDn+v5tNDvlA6LOoq
1xqBWJzcrx8av5DSNQs78Tt03SxNb+UWz7/wjsADakJWy+BrcsdF7QnmsB+lkyqk
4emtBtLKxNwlQvvLoa2nDtyMQf30X39zTP7VmCRdIZ5Nv9AOg7y+BGYmtwK8fYVM
MhdCoPk1gejYKRLVW04QusYpDoEOZymBBwoWW5156TBXvXq8P4lw9PQTk7OmEF2T
uMD1f+gwl9vziPe4zYXXYwY8GVB5WZ4x59Dq1ldPbDS5bsZqrdUApI2uBRYmL4f/
qxBYtGhw1rEVfxLPJ5T8XNowpNDsK0ZKcVw73azvvo1WFrYlW03Zdnf23CTpGoLs
b/V+SCGQZRZFKOr1z2GyAoZAknclH+Q4htbOTkGPZXqRF+YboqpeUV2l+7qYbAti
8T2CuZgnRf9NL8DIFyS22HICJkMsTHIKPpVLZ8YRIBSPI8OXFr2noo22niofodbC
FUgYaaSGJ5mWb7ChOdExXD9TbStlmWjPhJ09TgDvO8iBaUmh4B/VxGVC9hSBQsKd
VxxTNUvofsAoEvurveHg+JHEOumvis62j0BZ14aUqKxvyRN57mghvtJz3mc2LNG2
F+LS+GDu4SiZrAYHziWyfWFVmsNEZDq6czpQX3W735i8ocSloggPaPOU3F1OlQt9
kb94gzZArPHcMt139AUJ6ZIkcynNWwx2elJuZi/ZOFEESxYHA+imPLJD02ku9llN
ca66ruvBVKuDTUa8p7UOTQQOvcgyChpMEUXbGS0MWxFt52/6KHHizuv2kHHonreM
M/LfFx+PfGMS90C6Wh0qUVr7o9wYGh5eT089Z3ymkxmVdZ6QtFxf6j+aVlq9iWk0
D+JiJgskIdlQ5WaDI8RaUPQOtFZLWqdYKLD68UjQsB/zF/vk1pmG75T5g0TOcHwQ
l+0yUnbWJnOFMtfgKoJvqnIp6KjHjIzb2VAjTgluOxs4HYJgd9Cgq027AThwr46Q
DXLWb5djmBDXPUrMt0E/DUSMVvN5GFApy53JPfQAYIchkc8zlmJyRz6fFRY1wD8q
KPJhwIPzWu94I5juqC07oCWYw4DP4Je6qVbzfWQ2FnkIEwpcWNgWZZPRxSkNDnqU
VbZCTbQI5al2Hrw75oSNuIua0wWTUxeIZAhbUwcGytIoZoxhSvhNbAwcCfqTLYnL
FImXjaicgpcv9WxOyT4W7LNCI2MKsdSes3rFNERgyPVcZ43GN/AOqHAimzAdQz5t
xHa/KXbj79cizC7/DL2gXjUi0ZoPRussHEg53iCPstVkaiJ9xQOrfUmifIDXccCx
zq4jmGuupIFtcPKyo4NrL8oZxX1g7tiBI9mevAUSO5vrwkg8DQkkxQbZVnFVcB3K
mzB85qxBMxuXcN0JV6tmDlQXCgIr6hDXOVLtgIv8qfsdVehVdzrkw1dDVQOe3r78
gyopA1fn8emW24gK0tv7BOQ4yVV++cZkc3gZaGZzLyakVPM6hjjR71orzDgRe8Cz
jz++G4T6cKtztkR33kccRAR2rRS+3DE6eBjEKx4S4twPPGB/HGU22ytdihsNeUcE
lbefp7xufpqIerAtL6SGNOhcIGgWg+bRYcsvAUmyh019gbSAs5qALLHOPIBvaKi1
QvQZvjr75fRjW+aTpv/jQfXe17KiLu4ze31+hN8pWIss8CzFrinXqoF2UTa4xmY2
nDC8tZEMNhx//BeHfWbMSz261QELuJt8SocI0olie2NMjyte5CD5amR1UwYcwoDO
18YrBjqY1/qqZiazrJN8J/nACGslQXrRHrdJ9jiFoOrc16Jyd4trpYkTYvrCFtwh
lUXY1iqf3Xp6YHp0Aa2Grkc0ig+Xpu8yklXcxWcZOuTb0rYic2VYLMefbE8vOBgY
fx3KRFm19j1Y0MpYyj4Y1TRyLo8xBkcm4dysuZ+ruDBV9FGBi5zKc7IKMyRuOBzZ
7/vLgIaN0BlDqvXG4px2kisInLs5YCo/EeZR1NuPaB2mXCWzil0PblK7u+sZKAcB
gwIb/e1bp27PBPrHCDfuKImo4mkPWx2R/rCqw7TEf3ne7PQqf4ORB4Srst1LUDlv
B5q/nTwVyJOOSlW3RiRrE60wiwOfmmiM77hsW29B/1umYgFDiu7447UhUknzqqs6
E5P0Q2I8DUa9xLm0+Iud8m56bkXz6onjp215CT6QUN5iiUTttaIE9R2gLmg/u07q
mdpySQq+PDoBetVi4abOFJCB45Qbk8uT5tt96hcsDoDpfIKpxF2D5c59ZLkI5o8C
AI2Hu6tCmH7zN8mQEP9moBtbcnNaTJg6SElIO5K2k60CXEmj6IypseztaffHvJ0g
HDtbr/DOHcvzKuMkZ9nQ67BrAjaD0vB6fgDc8Lxql7B47g+/J1+47302AqkbB0q2
tYeezJ3oGftfSH9r9JSKjePlwoU1oy9VTgF21/OPyDB9Qrz5M3/rTlt35o4Xkg0p
jrD4HsCc8J1M+SxKVGAIY/F+ZyR32LxRr/cC8dcIgHnLDdXXTGfTf1M1Lyi2Qz2/
IkjeFbvAf/feF+pMim/6Vd1VqfC9d9m8chmtKINNo7u/UDtOIprkKa1s4iVvZdOy
j5kt6GC6WE8PylTLqGc/5kuuim7mzvq/baBZ5R1qS6TX+bDL7CmRKqVeejU9PrBZ
Bk6vZi15XtJaQVwbbuQgLDdP6HmKBLzXm0tSSRavIMfYuoiEzOK3L8r8ff/ec2bT
qvtcIdrmW83aLPW4HYOOgO1qiyAlV9NJ+IwU3NM0Mw4FXjv02GGTns6O2mu1s9ry
VP3FF+glc75+XAoS3P2pRl1EaWDETfuMY7Mzpcu0mgO05wVQRLuXBMmdkX6+/FMz
QnFHZevirXxCb3hOVk5etqZRh9UV7vipFyki8lTFLZV3BKDqSSJtl/QXzYaIPtRD
Bj2FdG9acZVjyH135Sx8u9WBAbqFA3iPiwYST55VtmWdAKlzzvi+4pxKltWicN+4
d0vZAUsmSEREcaJ53LTyRymtUzfRkBjY0CSaAO98j50/16NvS+nzsuRYRkAx5s5L
/6z9/HDuHxvM8Xp4Y3mNOAPtZuhdxq1d/lk+EEB+3TNzDdhnkcz7S1LkJvqDsyfD
Sq4j4Tm21WsfWKLo5/zJDO0bvAj16PkSJ9js13WpgtyBy/Zi+4TkVuQb2Up34nGb
C0o4EEW/ySabcP7KsAF7u6/EWpiT37unxKHM8Zi8W8t6dT4h+FkzwVoxE4jhJH+m
sL/Mn3cdQ+ACu7Ik7ty8TAMjZrBKUv8s/vOwhxgSAgc+kX3uneRDAXW9Oymy7g5o
IkS/4O2N7efqCjDLA48gt0/8tlkHygmPleV/gaDiUOhGLbQzlAZbIkep8f/vOJm7
fTFt85mC7Jct89KJ4I5RIIcZrDeJpH1jDf4LaPBZA1Z1kwC0MIENRJOdjiP97Qm2
UtimbuDtqB6DSYAK7ay1AN175C34Bh/mPattcISonGEckYGF6WkCI2yVZd2pkMb+
TL2Fq81s6dUNpUDWqmqt437G0Oc2G1OZRxTMZAlc0jP6Ju5YgnKLN5ksWHCaS1M0
yBsKDILItG7Rb6kHgkbaJ1kcYA1VWX5nRXaoxh5aFUeDsK6dlS3dG/LNFJzz4mGA
6vix50SfL/nS5wlIBAR6vMseaZFY67Brjsnpg4hyYsqsguMYdROqV6D81sRXumz4
+UAq1rnfRqAXG0rHl79VKCHMsZyvuywdm6YJVagwHo+P308etY4RGThUmTtt2xHW
TYl0yjujGZkQ58v0VSolihVyXGxK6JRm6wosx4Wevf8PX0+z0oDhsI9dyLWDDl8D
gv3VWDQAof1FznqVsxiU5n3W5i7pIHKEy+hR/kvy4FjekTWi0PLQY/NbJ9T0qzpR
LWaJrO3XhQY36sVLFQFa0KAw1qT3zIW0+VzOq16g1kCkr4lAOHGM79eiDO2artbw
9kQzOtZYRZvd4az7LnFATMdpDYadNzHq7bw93siNlVJqLKNrRYNH6MoxH5wZ01/0
8UPH8fC/TgIig0YHvoIytZ5hlTn/0n0QikKKIyJbB3f+tQAUMsY5k3hesuU3VEPj
Z0ieiMnjDe22JiVcUz8h47Y90irzcnP9roxamWw+fsZBhP3YwZaeoJSAYkMaTjy5
08+kqgDBzBoG+6YBp/2FNZYwwipXgQS/Sef7xXMmboVXhIF1sCRWHo+B5U/zPYpc
XqlEugJtgUGvhQ0pAjehek1ZCq0LuGmf8rJikiYhSyTJs/iwZiAsuET8er7cYe/z
LQFN+TfhcroYA3XVAGtJtm2ZbOPOyBqvnv6/2+pjiJKNb+5QtGCqpJwbxSpWdVZC
3um7E92yimmSuJP0S215x5zYjvqmPT/KmXbYtHtXgVm6nsJt2jrmsVnNMLzMv4lD
JS/iIj+vTM4/qrNqqnP1SUYV7J1jrcWWdfucQvFK2Xe/iWCO9HfuFt8uMFoIAuXi
wjQYqI7/7dNAxIHgo71ZX0aoQ3JRUheuWNA0VApL5uaTRqIMs8l1J5swIL/ZxDIc
FcYF32n1HXVxWiSEvuVjy2gVfAGsoU4CXf+0dpIiBiQcqEfo+zAMu0JhLc4EfbWQ
YKHwABrAjPBgdniheIuXn0DWXZ2aNnTIGOjI7ZCl0gPnK5Ye2l9P7tp4bDOOnyNc
9rGPBUGtn2OqENARufvRObZnKgzXe5+UMZzpQYGMBzfj34czCwWwpzrtb3/kC2jx
Vc7Aodz6E9xdzrRqSli6R55j84cP1VytZcE91sNzWkqUZoe3JQN1hoKxD2Tjt75B
u5SquS+5gzKo/KPXGMMs6TPus4Cm3STUYqpQL7rdYJZ2o1URtyDP1ssr44KMYx+e
WlCZa4DOzt1ImWclA9lvAClih2Ud/inVfG2FarcazRj9soeoysI1VubXae61QFWU
/11rG/W4ad9fSgwFUB3dwzUry+RxCO+ARqM0Rq4E1Z5rQOQ6Zm8qQJGkhTcTGfBT
o9svn1/KmAXjXiXNpHWUuGV3d6wLFgqR559EqQoYqhw7dY7tfFX/PWTgkmpcsf+h
kMY2uVntVny0+8fU6rcsoyK5h7U23gszEzBhRL3bTYFerVsthudybeR67VgKIU27
vf4XtoBQTyR/yDwiU37SYZV6rGntTjKy1ZoOwV7KFepft/btYSLpv4Yhv1NyFwNO
GBFM44fQE6I9yjvM16te65X/TeXRbjTauwYBE+GtuBMGZCY5PnYLNku0NxfDd7RK
yS8OI5NE7yJh4j8tof9Q9PlC5P71hOdf6GJJIUJ5/mKJ7TCy/rbs2djX9GBvkj1R
gTAPXaMj7bNEle4jiUjs2jMPwza8LNiMBaHH40lrys+1OPkHwmwC9pinZjOCi9OG
KUVZ/08TcuMaXjw8biFADDFDqTMBFfrt7WPMJclw4dqeXknArQbdBoThcdcQ5mvv
/NWnBiT0PnaS2igykg/mbj6hr5YWFolGibzSX+fUkOIO8j87xATDMdrFjZdWf9T/
fr75z2kwdNBuerjfgIX8plYNhH3oYngaGxS8b0zJSu0rGzUDbc56jQ/dBIiUkNYh
zVX9W9kidBhFfKrGx4YHJGrVAnFIc9koBzvR3HiNNV7ScaPkr9+Hp5hpffUuw5gz
+M2HVBKAJvd+SIiJKz8H5fS7BjDrllEGB580DsGNz5Tfwb5H1XEhj4x1d2uvFom2
IXKlih1Zj0+B2y12LwDx7WqhyfD5/pLZh6cK9P37iTQpqSTYCwiALrHPJ45lpwYY
lsWTyHKOCeT9nIi7rAsuh6snRlfZuzPjJGZF0/g/a6k+923UmIm7uYBd4yA2v/aI
M4suw6AvEW+GTDYeC3RdHrCC9y4BNqfqUGPQAVz/PeT2RrvB0aA3mjGZYdMNgntr
tV8Ohsv4QkY9wr3RrLGbIkXPYEzg/0XZo1M8QZIhbuS4varwDB2aWcItTWVN2/Ar
pjb1rVlQMBjQJiJiPWmZaAZS/H+LEsuS6hxBK2tM9+S72l4Pfw4PtuPdTMFs/cUa
i54UcwDL68i+ONwQ+fK1uMpEaoDPLDENe1TL45zwYNisJekb1pp5lCludXl8Z9sY
40Mdp8RqInz8d8/W3JivV2xczlqSmJI5B1KT6vAvxUaC9lWbmbqFuiFeaCi75M/1
huvnY799UBarU9MtO4Ta2iSorR0MQBctUllOH8jT4mwze50AJNLqkkwWRjJmNm2Y
AciwAVahoxbl4DTg1q4VHC+KnX3ZWHxRFm4fSKu4xVgpkQNHsJqDqklCLqX2XxvC
WLNvMoDF38157pzF7NoyWxcibY5oIUJPdLEp1loZ/a3EsA3MK4cPtpNopsoE4Ee4
LFCDOp3vgjgjDVNFasvyTIF/jZ6G5QrdzyGdcmqGqqkEVOUmt/bJItIBABA52QBT
ZaCOVRFWrs4PfXNQbUS89hIXdj5iObeEk2uvUlg5UTiO2jnj6zxb+A75kQKFhuF0
rwqG0JNjLNur95ZwatRYI2VstTHPJcTfBOfF93H3j+dVhW+5b6b5RiccgTluinZ6
PPUvFJoccOu64mgwm2XlMc/gSe07yOX305MK25eAQ+aOrepKMsO/9+IHLaKQymS0
m2Kv+uu5dFBzSWm+JREVNiDEOH/KFRxxcNzXQXKiqCBsz2YvxnPEP0uDkz2oOP2+
av1Xe5JtG8ieJ6J3eRCmqHVq9pm1MEHRRNSBRrK+vGT6ZyYGNnvQJ2jBBJhD2nv0
WJ0UAOL1J6zFEO+NZNsIowxmebIzllDOtR1xPrWiSULuZUbcufnsI/mg94HifBwu
XNyMZ2LKX4tTayZR+Gt3oSwYCWAXajC63j/z46JwpjZTKEvmGTYAk2VmBrH5h3yA
49GWeoZWO7RTpSxdSXIMBdhfgz0gcM79edoaCTvW6ij1fGQxLEz0hr+2u2p0TyE1
De0AsbtdOMkiPAkxfKfKJYcPVkCFaxN8+L6En4uF9zoHQOyaa2+k4khQpO23kvfq
k7bnVdzc59FZj5FXNmU4ZekiAZwGi3oGrNVcO+8C1dj7QyUjgJBdWDnDNtGiw/+7
hV9mTwqhNdGW+X5kJPYjfN6RoA3GjGtYVQBhEFzsCkRAcsQLVAXzJ5LPsDCY/bfA
Wj1RGYzdpwe4UHUyUlbOSw5Dj7L3kGj+8BxNJ6UgXaAKy99r40d1HcTOKnY7RMjq
xI6rucKviV3nOK8p2fs4tKsnikYQ2Y8y7FB00nCu2lxs6lncqb73x7qZJuWa3OtW
j39SI22nsVMPbyErSNSqiAdQY2yfVmGqbRP6QluqZrxc9vwPrB4yvSwUQmQ26DI4
NL6yYi6ftUuR90PxWfFmWKGCxLYwUnTaEUWYQ94XlnYie69jBzQFWdYKjxirr8RF
bJtwSEM6a7lKtv++3WhQjLd/JjvN562/pOJtXvEtdivwsIMOTMuDuFxY4za9RcIH
cXj1+/hCLeFfUrRr0JvhG2kVPLIB5hdErhXRMn4FhLW6WhR23gqnLfvlyrkf44YN
x77gcPBOrvWWeJD1ip59QCMoSRSgvklAAbOZp+f1LigOShaZJwQpaMdBLV0wW9t3
K4Sd7lH2ywXtprgPHZXyBptgilJZj5ih7Wdc383RtmL9yKd5F0fHXK50sFfF1a8J
MpXoAd5aqv15thGS/lP8uAsiJYSRW3jC9etPiJTfhAikUURCazTGivbdQJ/B9oZq
wNJZ/JcrTBgFgf/zlWwLS+AuZeScXM/jlO9frhIbmSGVZEjr/xQDpjNSZqi7qJ8B
11+G7PRZn3KRTjZGk/ThIfSzpr16b7vE5cYNn4zmepUArMaySD3VtY79zoAW0ZdX
hJwxaT36JfVLYv3z7QxJYDA8rXNzgKokGIKMwuD2ucvlvfC5kfsA3HobJnh8UfAs
fk9qJveXFctZE0iB7VAyv1txlTbOydd6yzbDSkFFUunhL4wc6eOydpFqKtDrMiCi
V7GSI/nIjV7ahzMjGDW2cbOD6w4fl5ENU7mI895Ck9egpPSvapDt9CGZDN8nwWyi
HUQCe6xm+MVCMRncNTLURQmsCjtGZ7phSGNMLrC26iWBjJaeXcvZY0ofy3eagoio
Eui0oz/yEKVMfLSCoZS2z4Dmr4AGEinYDRVMAzOwqvMoBCgdSspCbduDOsRv+wdg
4cSTNFUxSKjAwww9Wrs9J9k+lU5iA3tQ21L1wOdgBKUc40C4TuHmaPPWfpg29+PQ
GJFugj+/vdmY0Mm98Cm7IxrC3Sles32pEiZfXjkSfBBX3kCOSpXYBmFy20ZD+m9d
fEMJ2bvGqh5CLT9BIUOjfTOhL0rcbHGsseGx9iyK9IBBMt6hz3JE1F0gLonFVDNj
cnRRShk8aLL3VZHj8oQQyQI6qjGFYDF7symxwVe7/eieX2viB9eZQal4Y7YCNfHw
CszJw2iG3EvBjHeDoz/ELWbkiaJslA+sEpDMs10gmuihWso1IOTtCzzM2GXroii2
y4shW1FMmizuyuQFzBvORP70QwfkCQv2w7LENfB1Z8ZoZd2XDKVNo36ikmVxR3lv
XsWus1O2CKoSkiG6hrtKZxkcNDJ0WfG4x5WZZpFEBpgOttG7k272HCDX2mlhE+yE
4iJwSjV+HwGgdgxZJMp3waEBGVcTer9g7Zl0BrOUU0e+4r/lSyqlreYddZSo1ced
tQIuz0NiP/h7+JOubEt5tf2iHyHthJeHSNnyE5Zx4Z81n5VXiICrcs5A4wYOgKh+
DggTTITY/rtpltLrFAi0fmxcTZnNx6ji4yE7MUoPUdcVPCK8rMmGxzcruQkvmG4G
KGuJ7D5KoScqJoIPzdaJP0nGvChcxWOsRGcFp3AItAId7Par+KfqpFuQGA7RU2QJ
p2aVyXuDrWnF4hTvmgdKdBVoqDMn8etKbKSc/TklIHvnrOvurdGQZfOcdV5gpFSh
3ECaeMUm32ZDyV+R5IptFPaShNQQMn1lVsUeAf+U0JHwcZ2EQYlvnzp9kP+XXfsc
kgHuR37Z0lNbwpPAG9ar76fumEmBj7pAcoUgEuauCY6FUSIvPH74Ke5rulpZMMXA
1yMRLlpoeJL+vngGThdPo6A6ZTQJFQpd6yfKN/g7lAaMg56fPLAP7YesP+uggU6I
u3i23Ns7V2sCYMlWCFjryNvKl/I7drcZSdOWRM60ZsLVJhLt2irLp8nkNYGVlFh0
TCUqJNqNDz8fHCqOXzSDrUSAxgwWiXhrnicJrsqGqGVI/JzWpmlKDkKdFaqBL1QZ
KEpCgy/b31NOJ8mr0CyOZUuv+Rl+64i68gApC7RAPIRfYXgTAAqxlTggFQNp2dA+
lNlzEiZ/9OkVO9iMrwPmZIlXHWa7cgFxlBwGVmIgp1rbYE/dguynqWuyde1nyWMd
5sR9eSqAIur/0CWNar1KWxy6QuYZn4WWi848icf2I68K1HLzvaB2PeY02vKWwzFL
4d5Hf3/RiqR57qdvLAY8eu5Nc9mg/r7gegWuzes/IRKuql0YTCUC5vRasAkjvaKj
fiPIbC3j1Xq+olq4DLOOeLb/dSDCNBTnCej1ty53X+4KIaUezTUnJThC/jhvtgep
kosgNGFp58T0tULEF16RyFexl0cJqsTNP2sNTwylFMbnntxNUCKFo5JUHDGBtUJP
BlxKm8v4I+KR/0T6+fCcU73+yDZkbkzrn1uEkr7GTQtC47+hVwx8IH9Tqe0cbA6N
viIIZaWNbo5IQUUlu659MFdYROgLRzrjI/9lmHP9e3xcB9H+NErHs6d01tsSbB3H
nzse37ebpFv+DZgnXMTjPcdnV3QkGZSp3ZGIg+r6LtDLwElmvTI6JlBb18GbBdD0
WAJDc/vxc6tQfgch2XNrW7gtZTQa3zZe7LQ/RvHX4mNGUY6nigtoBH3sY0zQUwMr
fTXOoUgWeQqzBwNtSbVVdRem14LlUKJgtYsdXQTVVWPjjqlTJThgzqb6R7U546t3
poUHfjR8yUD+UR5ZefNl9JWsB5PRKfjgqUfBuagKUcGZQ/2EDC61QZideoNmn3hm
vplZE0ZpljZ3oa4jendeVTOWj9t4teJQqJ0QUXvmMCGe6CaViBIhC064lJSh5xmA
YXtzhO9FFLXjdoVLU6KiweYah9+1Wd3hF5tO861BGmqNBdNz7mFfHblTptHL1hi3
dNdchSE8xW2mnJe4o8RdUtqg9391kvqGOOLyxmUl7dmwsrdBMGJ4D/MYsVzVEmDc
S5BrJZvNMBBEPwXRJccs9qKnDZ9GlM6OLfgAtEpCska2SbfWsrgq4eYS20KqLFqK
LklP5SA40EJOfZoWSiYV8mvjUUL0pAuQvpsD1PGxD3N1pOkeN2K9Bwk4n1eVda9A
BLLo8i0ll3BK+5s7EWPU5XJcuC4Cw60xUWRRj/dXgWjaxsmdXdQafnv9Ao8Yl2vY
4O5FNk9s5WXZS1N7703YLbC0R16GvO+jraMwXGeDV4+WrH37cKMdtn6npMHHGoMd
jZh2S017TI7zjDQC3UzRVAIjMGUfbZx5/lN+LwhRdybtXLR1MuTXkE3IxrSWne9V
eV6EEWMMQyJ0Kw50NaQy2SvLMOSwmqjofXBs9E0u+a/glzYMSw+VAnC0M3Pu94SQ
bvtOIVA0h1z+EUHD18YQ8Jy3d/d3LpSikUOPiE326SVctfXkKvJcEL+78vOUcfpX
LnqsHbMjRHcvy7Db3i0MPusOCxMbaewsS0uMD+4hlLG2GSPBROabBgYB2LBKUgEA
BWjbteLUwclnoIPttoTHRVUjWDBDQQcRomSb4gA/QvWJkoUiLtNEUhSUPbd5VMJ9
g9zxaKMce26fO3nDeFRrdgp5T4YBLlOTzwgk9F9jI1cA24B01FEMjZKA/Bya3p6u
v+xkk7Vmd3GogA9ejsQVxLxA4R3o87t8WCakSUFqM4EhBcCWZtyeefwWLyWz4+vA
psljTtreaOkwjWr+7H84IS69JmmEaBokeanPGh5aszTDHuZXFmDPAm37STz88Do2
muvXh/JuJ/+33c3HU9WIhXI4DieuP1Yu9sT7ET4daD8ZzkMtYFOsWLRvYLPNIdHF
z8gT+52q+Sn7nA9P4Z4hO/UYyqchd/yebM4hnVzERPO3mpnpqodBwgMfqqBC/t4j
iLrVwdjKFKq4vio1me4+MYxSTX/yKM6cWNFVyfsG2p73t9hGu0MvodlGY9ThyMgQ
qFwGMyGScyRJmIctrI2mDqsSmfqe1Oj9ozlOPKoWidMx7419x4gVry4KS+n09ObK
9QIDZHSatV7qRkZcsJbIZHbfbb5KeBs78UESqJwP2z4zheiiw0zGc3A2KhiICWIi
R2MJb6FF3EJSpTazBOdZsdghgHRVkL8Rn3PPj1fE1Ua+KFye3ecGP8AqP0d1KWxV
YYUmNssZRZqI5cu/Ei1q1bZjCn/PRqYvSAE98n4/1xR22xQO4U8T9Tz0oyViY25g
/aJ+SQh1uyYSNjp/qWR5tfqmRg5MLuqOlQMSTrV+1xLPOuEI44/pulqCQG41ovNZ
UY+jBtt0iGs38OyZ1iphPudL2BpFGX0pWk3cU5IZNp5SSrOlLSkLC8iH9UfljUs5
Lo3rd65EdwcmpYn6l8sTET9nwtBXMOoS8VaqUpUTg4jLJcZXvi6/v38/vI0ljY36
CHm+/UUIK3/SbdFTP1lg134FXgp3FeAcIsDVddG5AJE63qwuxFSzvAp0ktrqoTKe
XIYMqLjSsVyLikwEl7fxootXjrof5IqBTyEJ7zPtVelI1aOAjxU5q7YPLzzPWF1A
yZFZ3fIjpISWt3nIz3pEc7/yyWBmt4CR966FB4UoixQM72/phtygKdjSpMegCyHa
1aV6Fxvcz4w9emL7JrGr7+t95AxC4T16yl0sisNSRDSAIusqo16ZEERt7Kc2GT1Q
Up3Y9QTm20GX3+gUsXGQvWyBK9jGGnLSu6dG0gC0MQeG73c5TRGfia+ejAs+09+K
n8IJbQJGUE2d5viStofLfgF+D6wqb9X/ohUSLdUNw46a5TINN6Gy05ns6MrlQbh+
Im6WKSvPH8E1KMRlBD5V8rr/FbTzjsbnvrB6p1+PEcO94c6b1j109lebyrDmecnd
D8iq/C224GFGJn6SgNkSwLheuhsBT5IcdIGY6oYuYDgOLYXmvTSQTBZp4oc84PUv
v1hKN09sb/D9/YPmd1AjtqHTykc95ZLxtFw085wXu6YytJRGUy6eC+z2q1rM5m5C
i1kCwHXl0w3FC2qcoR+7dG6opF+OLznoumTN1Jukq8dw+WZ7Ro0TlmepeprRgKIA
pcxcaDRSXcbT6lb3XyJJ5cXQgN39UcoCPexB+F8qv6apNt7x/uSJzb53kcs0Kx9a
ACfhyj253V28cMR9T7PDkeAJf/ZS8v+mawY2LN+dUId0z3RJranqfNhlAWq0Kqs8
2rly5hURN4WSDoTTlaGgCYaysgA1LxYR748v7J4izuWUUeEQwJAaeQhPiMwvk86p
VP+yH0vNngfMWszSuVBVaShehZbO3tpBbhgBmGaDPxMX2PAmnK4Bd9q97QPZuTEK
d8XTbkCVWqnxKcouIswTeeX5tkipPZJZteymwM1ydC6s8fC5dqDM246eLFCx+tEI
4W6Fiwl5rQR2qIZY9esT1QNSmT25jKk8EngG5a7xN4p+PPCd1NF314CwMTAy3LB/
rGSYgWHgMsBGT8d/dg9CHoQDPwSMjNtubEa+MigSevUXqi9yhVSc4wPemrs2/e2s
8RJ2fvp6ZAtZRVTWRpNZEI5me3QnABh8C01LHwIpdd3xlu5CJS+dMgl8ryT+q9v/
ONbf6vO1hP0ifoMGWxbok57CJZSndmA3LkzMYM0Wuz/2HQW/PhNL8rZHbr4gWlbX
Bs7pvfSC+dY+rezKmRdNvbN+8rKsC6ZbzN6TgDGgs64M6Zhz/8ey7Tt7kOPIzNv5
HG3Xwp7FzVp3jm2Rmfl0Buwm9IJtGpiq/J2gsJNO5KdGfPWulg85Qhg6IkAhKh1r
iMs8HcdiAIyOt+kC76ZufrXxoQPUgBuSEKvbAUKFh/fyqAwKdC2FThvaa3jkB6qO
Pr8y4h8ZCXz86WzJEOust/41vKQwctzz5qRyWtCxLhOBD4C6YBX0K4/sXqU7u4pd
BLa1iIW4tHmlCj6hC8gsasRupm/jP0bTuIXvgWcazYrQKetCYEMbD3DNLF8USRJ4
NyprWoALZBjiZfKmVfSos6DnLM3+3EsEL+5NX3p1GpVefnVLXN1jFmLHQv6xbPrD
sIjOa2ZrdEyunVMp/A9/0FyPRVGE+Dkl7cl9jr5r6R2MK4xyS+zcPZKXCo7m53yp
V1ZjCBp9LvnUH//PMCQEvsBpzqeEDLQuJ0/hkjVebrjNWMhuR066+Qr6EHtqoeDG
gTLI9pRrc/rXASGh805aWMu41YRLuS7g1ToU7ZfgdSaEuPBoqdaCT0+y9SJFCyuc
U7B+ozt6NPJgqWaTDK+cK/kzGlFqqKDcruUNBsbeT3F7e6N7AZ0D3pLWtSe8Fuu6
0uNljMQCfv6bas/XCvnt1JxrGiekWk3rHJWCLTCx6Z7YrySegl6dO5OFtAq/mpWx
Mu0/WRzbS7ECR1VajS/N+WB9BV82oUcSmQeETJbfT9L2ibLaz7jxOzIrZk5o9F3s
krUeq4d1+BnsXaE/zSjCGks7zLBHZ/agfwFKvchxuVf5jB7Dz41gDWwRluwIoODb
3BM2QneWYxI/IYVKiiA3fMVFoMx4IbrZXg2ZmDJgXa1uWxGHgypIA4YZ+9jX4Yga
rhOaGPLPJSH3shWPauBOkrGCOUUKXx6FdF9NVD1MlU21wuQ35liKuMmMLY0wHiY3
/uu8x4HFAiEuQezws/nX2xLo62auWhplDJ+bs6wF/q1yQHIgJnOJftDN4y5OIgUd
IgubRwJPrLikqCCWWZiAVWFE2G/kzTY7ormuxbjCxJuPrNmibcva3MeyjNHOxHYr
HEfF8aW0x1zEZQfu6O70Du5+CM9AaxeLA7CTk6wXPZ1pz6Ty87hV4gFksvWC/64a
lzkwxkxFGi4z0Dpjc7CAKFrfp2q2PZxlFKul+BA8PiZAQrKeCn1uKct5RyhU6G+Q
sXJy70dU+7qjfg0XFo/fJK7EwrDlmwgL9GmZjFswAoYW9PFXPW1LB33NLZ8I9UvL
uyOPIw4+fCoX0/na3bZUB4F4vmnTKsx/oaScfcGiB0B9XWG/Me1VWew3XLYl0OAB
MZ/Oqqo7L8W31feJFyw9p2n37oT+OzUutoTC3FID4m0KTlAwgaJco7Br/Cxp0adl
eTh6/lJyaEIOTZBcSv9GYmLXJdy1ek5HDWwKduGQnq0EjuQqkhjvKgKyJmX0ukwT
bPqfZXFL9zN7kRvGI9LB0/W6jCy7dLsnqLBaWgVJTEawnOf3jLnjQAHuTxZNWOV5
Y491AN1G02fcaDa/KGtFaGO7FtKkXKYRkeEl1JK8kgxTRUIrBSes3Id2cqG06K2P
X+93hMRGKc00hqhKwFyeoHrkUYIcEYk2139ASz3sDCxMbPWi0z5xszRj6bTn+Lr1
4Ak4ocyYchVv6dHQ1ZrOKRnW/ITdEo4spnTXlAxEsb5umFkdCutnGqgIIc21XjLJ
0P57+kyxNRzkOIdP+hgz0h5m0yf3k9qiZn9dJ+wdA266AQCkU2ZXXC8KVFaYR0kM
nX2HjsenI5vH1nlJfgL/xX4MebtoYbG4dXiRiheQB78MA/7fLHxkyCo50zJvzBFg
Os2Bld8W4bb0OsICGdZhitHto/QSl9qXvBZv/+ft0fXWQ3ATjRwQG9+YhlxPRXFC
3MQzopZOfMt8B+fcnXWG8rrRuIFJqD+yfnG85rGtl5g0J3gBW/Dekg9owqL6KYxP
ou3cB5We3cn+9+y+RTO8prZv6Fa+LxUYcSyxKOaZLKpfVRYquh3mTQZvnStw+VB5
xs5CM7b4fVAYOFE9Y6qRHVSSjahVJBdbcW62Fr4ihbGjrcddQvUu6I3O4J0xcgSO
vlOX6X1LczquNH2mA/HYtrFgSPa+5DVj62/IV1re8smuy1LmJZq6FcayjTpMSBWx
foojH0bcMBBkbbyctcwFU59l5HBW1bb87HfgGs4DUSNou+HMuRV60BtUaZ1gPrez
ZLaAYgggf4OXI8Sfz5wuPqVtcQLLIah0xMlnxVM1LvJGM70XwPeWSz4yYGNuvpZV
2lg+p3l96TVNZD/mHZ0fTaFo/8B5UMzYa4BrmE4VhZdQVL2/OD0wQ6sZFCq9B5qj
n6kIfRWPG9c+aZk8fmQzvYkPOQn4Tk/myAfvLGcPBXMlzZGM/k9uEjVGfTuHroD1
TQnd9VE19HisEIKojjei6qe1hsMilcl9JkzkaEFsSPsxTOnzbYW1UsGg4qNq8gep
bJQ8nTpFmM+JgcBzy/Yjc+wYf3Jji6OCbr+2g8Yngq24kzCtQdjFHvA8JY2l47V0
mPaMqD+BtFzK/8KgIxCJ1Pbo7vRjFDyCmciW21/1Re0Vvxr1Vxmh8/b2Xztofzl9
1X5JYNfVpQjfgh+kBINZ0i6RrDIYNGH5h8x1vKc6jykQkuYNqfGdn6ERMtT9fuTM
Gj7fW+Q2x8ODegXjEsbdEpiZYzY4xfBrcoVHkOCvrmBRaBN9VoJtKiwnIxHq/drr
h0+qYGG4wX7hdokTbB6Q6yVBjiTct1sy5xIYB57M+G2FLIvoMMZh+irxloZww06k
SwxpvGPbs7lkbyDjWTxpTIUmBA6KJAYL1xWWl778F3OrEQrrptTNpKHfLWKk22Uz
gWXtaX7AWlgp7EckRktYEOWztRH+TXzRhrsZR9E0Xu+XN7MUlt22Xa2ejY1jd7uM
4crFZfCqLdXQ0EdETolLLcj5/NfTA5Wf9JN9jiE7eYA69ZHTHajTO7bQ3RSzSkyW
M9b3mO2a/vPLB/Dzu4Oz8BSjaFiMiBcht6UUfL2p3bZx/zmc49ILRRaERwmuIGhs
oqSOfFvLDhjR/MicuxVqVq6GJbqaC0iPe7w3Z78HUMHu05OUR5KGarw0D7R8Y6Ma
dN4oMLd7VcxlkmkrPhcXnFURRDCRJLPCHlYhQTeX2j88E2U1P9LVX7EKEFPxKlMi
ePrQXqO3rs9cFro3+knNt8eYIY+M9ZHPSL3xBUiDjU4BYQJOEb207ovmX6/D3S62
k6rEgjf3j1OzX4xEQgTx3VdlWJLImup3PF8PcisK1frNgWIupcWb4hXJsymLzQCU
fylpPpS5XgBjPAk2/h+dwQQMeWLcKGq+mpTwD6l5U2/NlzQ6jnKSvffV9Pp2x+O3
DpjfVMjv6BcqsJhp7Is/D8ztJ6ArSAXZB+m/ivqWBS6PyCz46VQhFZMjJ9Gg5prd
8VuCfz270pIn7TufYSHBRN9+TAFkm0DoF9Qul4Aexh1lrsnwKA5vv99qZTCigSZr
MegUmUoXdd6YiCJ4CoIPuXKOd/LvZU0D4JScI/hLHE4X11jpokNQKsw/n+zE+3ip
37k08JhrcUwAZ9iyPFnGN7jDfd0UGnTS2hMOGWWeTBdJAfPtMnz7zekkgCBTNs1V
7Hlf9HtTd2Hf+JRkfRtj8AOFtTJPoIOjPgTU7VYD/eRhojAaFfpL/RYO7kkveJHp
zlVHJfu5lWeZKl7qcdM1lOSM5FEKu1VBxGFBO0xFV25PAI2dG9QRbtQ/dVsgEL78
m1Q34c+rHZjb0CN/sln+Jm4BtE/FY/nV3coDCBFzmn6CnKwpRfTtB2b/atfa7NXe
oFuWR+8TvZgJ4TsEYtodizV7nKOZvjj6mfej+fdD7YvR1RS668vGa/Jdf1JpPuEr
KLDT8pjrkzs9R17accxbDbW56nYfMUrIuSBjIMSywmLaDZxbKBWraYoy13TFeRqN
pF8oRUa0ehnNLYJ6YKbX8w+36BT+Z3QlkE9cAlBiHcGN8JFOzQuB0rx9jAj7wz1H
JSHFcbq1JHna2JIVSJI1MgBxxt7zozpdXSAIU1pCjw379j93+CEAY2+dLJdw8ZQu
uWBUWVj46Bx1vSYuJxnqpT9677PdxP2i1NHG/MXwdY5fPZTWrUl+J7dwHm0sLgKA
Kqe7oJQSnd8RZ2eyIfyLC18MaOqajZNGavIfAL+YS9NKIyq9r5LHqfh8NanggUjp
T5rJtXNm/kJUeweo49qjAjXl0zHb49QeINFkhx0uXMz0EvqCFP5rAWDsHtZk71Ml
k8/pj77SsaqvzpB3Uz6mJJ72NnVEGEiuDj7Khs22+CpZYLJCjNscyYpbdG2aBK1P
VuP9tVtTPNu5Si5Ow7IuaWTjD/WFwSM4cluve4A6IakbpKmeEbxjAvkauthoLRT3
KEK76aw6DC0Yki8wLMVpOFM1oGgctyZAMcC0N8hVSSol2kFSsK1EzzKkUqXdWpCG
+Y9Kdlmx4hEr5nrisUfLJwM2D08VKm6JlxP+9kOrkplZpZrSLWB+Zx6UBLNbWjF7
yEM+wjPnLA4KTjaRbXwzXEicbPOVv3DRilEjipQL1KDKZBIs18lAuQ2yN5irhO+/
l5H0xDdz5SA5S6NmWZbD0ptIySv6MYopdrw9HcfhtlE6k8mhzhPJ65pAjeF1C4Bb
rc8jjZw6Jq7g6DBw903Ns4YljzZnipVpKsAcPF1/+xiRWLPOlOQFOXCWZJbNYasu
Pc5ZNwxHsuwJXXNR5tQSFIQ36Xan33cgd07wuCFrki/b/bQnzaRSfrv/vzxXdkAN
Dr3XDPdQ7zReuUyUjQCasHICY112hTGFrarMquX6cBZ+YzHP9V1tA8tv1oURx642
BzLiCBBv8UR/z800jRH2llsQW0t+iRcVIL1uLSpGCEIJE8xF9rPxBlRjT466oEiH
V1pN9VyiJdJwXPFY442wrJqOfnqENJkoFbDT+YgWKu0gV6MrR81+NCpcOQ4EcVZa
9GZvRX6wsMlwygEEdXotKXEXHZSJasbRkH88grXQ3POhF+W3Am/0YN36X0kQ0qg3
bbvlR9OmeEQGoDKIK8hOzfXzmd3UcG/FHe+6UyizYhGQZJ63mNkXLkRrTLFDqnjV
GHvHCfwFwmG8RMTVQpV3O5brBV9cIfkqHIDaNYT9n3ccn1GxgWa1fVXaDE1VACPh
gNHNwPLn4O61nQ2D9XFIDmEHCG9410f5AYxaisRyamtigQvEq/DqnWiYR1Qteo+K
pykaXP6sHIV8cpAWtiOphXA0ZD9meMRy7Tj8Ort/TolRJZzv/MceIKMqUDguMsQN
hMZvfyLmR8cD4Fmz21OFezGUrEoAywXAzP8N6afKvrsL+iUPBPeSa+EPZVIhoiqX
Ss7eqYyjKS9kAyoW0rnpO+RBV2WirMM/0OCcODEXcdPbOJIMO1nj0pFM2bkHu+b+
SB5t0LqvM/pdeP1hu03j7eOxxoR2nJsliKBkWXwkO+OX0to13IDAynUpVeFJQqOM
mjMjdGqNPML3bTK/OrMlYeqmBpJNpifnDiH8Ee78v0ICYktc6MJHjV2cfBMNwpo+
YLScv+2uN6desIdnfzsq8n3AFjtVV5lLqFkHiepVlnfgWMihBNCS7+TCsLz0rFUH
dhFlCnZ6/3Y8Cnr0HI4zJ1cAPKaag2nbLt0DQJOWHU01QuWHnMhqkihLzfg1lvGz
BHWB6uXlFyX3PIl4WdETh5aTd0J1DJMymMqYycX+VoV7N726bamaf1TJhBJuQaOw
SsP3kapbKfbHExMfD9oRZnpAk9ic0reBZreWq6bziaYesAk6TeGp9zg1LIdEYWXD
RlwaTzYM5cT8gm8UBX/MGvEWFV/HTBvki5BaAgfFH5yEUOPNRpRTcfoTc/xNq6V2
imzCG02hFrSil7Fa8pKqeSn0T/eZP7yf/+tM7M9NU5vmNXZmVd+o5EjXK9h5FFfC
iOsTnkpVQX1k/9st5T03erZtAqueHOGL2iHStWjDu5S7dMhQ3g/r/LgVh2ikc8ay
7Q7Xxm5chMQ4KPZXajA/cvNhjcNKo58HcO+cFJeOhku2F9RBPv4Ldc/QcQzv+1j2
eKYRQdyUsOpicyB2sR+kBVI+X4kdIb9K95v8PHxl9RJx/eP76oREWTroh6yxqqaD
GaBev1ZKnR6vjZ3xgKXHndxk+a2sxOx0rA8CyLa+zSTOSGmQzPRtiKjje5GN20uE
N5LjuA+m/tHKlOX8iFQwDAewumg2uxmMhy1s2G/T5FlWxycCarmNxGSuIUQV9ELA
sHpQe0zV9QAFccZRZfXgfnMUYwnp03XzZxKfFOs+PPvfj1//OW571Zm2pjpYS7DX
kS0nAP6eHn3v+wnYBNNGLoqqUbEs7t9LNwx3rxJYAIPgPV4/6JVvI4XGBiSWlQmS
YJdehUiaPwu8Hoq1gNb+tROK20fHZshSc93TJ5vHFVxPXVw+pakX3UAKWxRadPcy
bu4lCCEx7/Lw7aTnWD9RaHXYyJUWd/RXFc8bRQGgaWeEuEAZlvzJHfVjQM1rh2yC
+mc3AvHHwNropw6oHs/4PfxvvC2u7T9LruqbrhAVs3WnjPXuHIsLSCGEEjJFabH3
NjWyNPys5RRSozwq7bLEw6hNhKWfi1Vk+U5EBBNP0MA7jnv6NnCCphAYheSFfLPX
2bSrNpYwqV8lkYKGLgHZl2SfyjMZyFy9DS/TInvNTLZ1qWwVDNPN/zlUnGM9Ye4u
ZLDcCCbZ6E8WwhisezuDBSrcRQ/xj9ZhlNct5z+MvyUSCnzR1eB+7EXsZomD1eUK
EDnERSupy8AJ/At+szT9BbF/g3uSyjWVA/EXOO1q2u7M3ty97l+6cHqWt0XjWjjB
p2cvHLdOUcgkNxfHWBkMY6+pFkGFonZJkvkxEwCvaXt4zISUjHYXPkECHuDzHQq8
WL61x01FOd7BO/g2XjnBIr7TY11qVGjFDfJMcS3fMWZdMgrTzRzd71NwnrmB+rl1
QaFPKryZGyirZjE5fXGD98mVn6dDg3Km0RHV9TvLG62kYujXFQNn0Zx4PuiXPty/
kuH9Km49Z/ac9PbMGVyigPRMZZ744f2H9hLXscCU4ti6WKPIURFSfSDAmBVeMNn2
pmQ39139mDYMeGlVBok+mP90bbH60IUZhahs+tq5DFNOZeyvfzOUZAk1Rvpcd43O
HDZIIOKW20YDvgepP2VkS+z70JNOKRZHR6rDBO9uEtFhr0GBQnyyyQiOPxTs2bnL
UZ+NY0JUGlwXH0ieVr8Pm/5bSIPKTQO/m+R/zLJWFc2tIvFW967UFRo/fFvo8KHF
InvLzPKy2aJ1w25Nf7J7Bf9d94YrxjJE5fHa4CAUSiE4YrfQ4wRUpKtpHLLEiev5
FQ50Ini4rz25Uv/C/8MtYPZX91t0F7ACbt+P/EwDrXjdhZhf59YSNbfkKdmd/Xeh
FK0qZ9R76algjBKaG+OZo1WGGDPxxPwJeWqx2+qmN6ixXjKBrwq2w7A8D5Wr4k0m
6I280q8932X80H+lGdR25Ct3RBoWGo7y3cfSdrLsOhWJUT47nKNF2d8Qytrvrm7u
0c/Voc/4rmoFSZWfjY9kw6xkX3Z0qMEjUOQQMQ9g75JsV1KDcYHHHsFUVIDbMWD1
1rWTdaYXrMKYAiE0ioRzAYmdmwOMlxXpp4dxUJBKmqtd5jsL1xNpeR+b07sreHpg
29lV3oN1+yt9X7y2bQZjAphFk882zvildHQRm7Wi8U6vQYbL3xbXRLHHHzFZNEqm
YdeIibFqY/RB09fLpklbdOvfYFLEazQ8c0a/UlRm91jPCieOaOJuT+B4+J+vs2uA
yTpBT4bDjfCXWCKrPxwgFfu6bXsBNsCoK2oO13F2Dbj/Ja1p34w4Wb/EYFsPsXXK
zBnIXGEYiObklwuz6YA1+TP0TanG8aIddQjyaNt0UzERwM9hsd2CHYbkdoce/CPX
9HFK9x/rGcWcRF9/8kAbUqytF7n3V1Vy1L0n9vTFAAorDBX10+VMFX+R1Gh74pt9
tFaEH98Mgl0Wz1KnRMn6UoXfPCcYfykQUvsIMUnjXRoH6vDpcRpdbvveOMPWB8NK
/3ccGzT8rlhMA7hUuqHJ/10tnwNBnggvUaXY4RjNkwXCdC8mX1nBrSjj4BBuKzuQ
n2aR8PPKppsjuHG11LNRNAuXwE8WrwZsX5cuRldGmOaau6kiQIh5etiEDQuF8g+D
/iLOnRqRI8FKSg9MxgTbiu5a7nvQxZh6s+2PjNlibxHwsa9TXuoAKPVtCS6gxO48
qOwWf1x6JOugE0Op4Nc44jCxRtif1YXrxqktM6pZIwwOl/yxYtf47Mkqw2yAYsoS
tdl0N6L3KkN96WpdTHwbWMTllyzThRyusey/To2DJ9807nGWDZgpj+s/7mrGgDOQ
GexhKClGU2Bjq984ZSuFrqjxbObUvNIoXwnQCbbmd3doS6yxACtGEph5MprYgiL4
uGODe3qSIajKEllOQ0ec4VfUfSii+aMW8RzvYxRHo/OCy5trMufvgrB4MMJK78LX
o/ErUej7ErwuphEoO97HsML6pPFBziEHhSIFg+C5zkyay2MI52GSSkS/V4ZKDMyk
+cdtBfPYl9MpIwDe0r237USdK2pM3vzICT1ZMUxm6XjUWc2q7NWzJxaTf0c84YAj
X7W9i8NwOz6rj6+Cm5O9OMnVUTr1+lg0Vh0tn17glxTE7cuEH9gW/4RvDSJhzNoy
Tn9XTJa9nkfaKhaceOrd9/3Vx9KDOYSVAOYWmvcjLnjE4UlKFSLfJFBRJeI6M7Sq
xh9MPL/LPzaR1PKJ84D84mefGFZlcon0NB99tOEuLwxK0LTc5NT+/BRtkv9CT8um
3YzkLaSqb3Pep3mh1lam1xdL1y9X1QOnlQJdr4vSq4SpJJGDZ2Mnsj6xW0YFg+0F
vxGvFy+5wSWnbcR4DkloyZgYMpVDhEmivvT1xqp2oXH7ezWEcahbfYgqsx0FJDEy
GHQwdg0nHtvwcL/iu0EKTBHQ0IKrMmS6zk3Yp4v8JAYdyejUDT9xpHmsO6XE3mc7
LbVRJAklY8q2p7tsNzzwvKHhvTOWe3IuFBiDXQcMN4w2zpY1w5dSQjSSvlEbBCQN
UFPtaMSbk12GJcFveg28nObm4dQBUKLsiSUpulPsVoP3jHVzdQazGwemcREyvFs3
u4oTzRbI6vI1Lb9zRj5u8UbS910cGwGS9IdQOa9xi45GxM/IrBaW+DK3qr2uFtwY
0Hdthk+wFSxQ/EazQVWyvWmlUUkmc71OdzTtzUijNmLZD8wnYkBIGfncKQ139oIy
goKy9FGOvcH14tJfo7OpzOKoHjnZFsc1N6HWY8ENDvPrQJtvdw8moWtsjsnMLpfs
WikWt7Zpu0x8sTGFFt6zyZ9TCein3eVPN+PIexXERJiPXNhdujarlGHzXpJaXON3
JsgMI78gXcgaYh3P6wchB350wSTleoFP8gX2Lmm0H6zxL1izXQWymd2OC2JBq14L
AnjTtMbBWDz2NL25m+1r+yyKEF7+OyA4y+55VIfU9z2AZMGISn1HtPnqLaJ76iVh
D96tvqIyT2uh9sJWu1TtwdN5ehMekp+KgGSKgZYQNoqZRxFda6Y5GYJFW5jZmbxz
EonfTkP1AGrlRn+eQs4mna4HpmAMgnl9mjpKFr37FBY+cW3fDvBb8grB2SJjtR2n
o+ThBz3njg6H3H/A0+EUMUYxqverpD6s8ahHZQbQYWWW75vEc1CuLT3oYGTn9M2i
i5es0dTGmT2Izrv2xUNeM1kvxZcloqmItOIHCmaiOpQrILbu/c8M5LlKtVXDTN1l
MgRV4xg9cfPHmfp8UElgzbkmb5KiES9jxjPvtI07IL4X2P+pRuotf5fGxM/oeMbb
6xfXfqkHtOK7wS+XHnsutu02k9Y94Lq8JvdNroMruMpr80csFCa2kodnzULo4W8O
RCaohP9UfVIMoolWgHU3OmEVORWaUwhrwfaGrCehVNay6hVyzZE/hEGVv1jUbi/u
hW2qxOovmaM1mlxIgJiw/fsUyVUV9uUkTcJc8fA4RAWU5+nUCy4zth9ihbaeMAfR
kdN2J0n8xfbwxFAEpsAGwz/AfrLUK4MyMcUUJ4awZGLvMyGeQkSIQaHLICAi1EmR
k+XpeGpj4u2EcAdaCT6Syom29e9hDuSbbw/mB98CqYJmpcEl/74DfMU0B9drznEW
8NaZdE8oMlOtIAqSARXMlAAkFWdPcmhBU11Ke9VfJMxViLtnEAGRcRpo1/K1WxAQ
AIlfVWd5IqB6E8MDzqftqBAHIu9hdxoWnk+xT+SzNw/+2TpsyqfGav2q3vAjNreo
VejDsqSCbHvT88QfdSNAvHEYfbEg6hhsjEs1chswQ2Mxkp+dmDaZH5c0a07jbiXE
IyXiAgWlXrgIAxaFp7S7k+9HR2q7OlUdMRR7IJHbcIPvflIgwpKIEYXe4ON+/FMM
DBBYxvcIjR9WYchMK12f3ljYossOlVJHGliqAX4tUz2ysmv4sob8x+4d4oKtUGxS
ALkSompE8PoyWXpS/pHkbuktoy938O6a7tGPVrwjBOkp3u5CDtKTK94MzjGtmaTZ
A8aOLM4FT664O7TLzq3Ys6tlRkLBZH/lvlegiQWTysc3i0HhKhHP08P0KbO+osHt
kNO90WC1hYOVB4sdmTwjk7wwKFpQGEzHGRl4GHAT6c/TbzV6egawjDPsIlQGdYdM
nzSbFtmj8BTYl41SDYYvT90z7vm4S1m23eUsDvR+TjGJHRxWqBBtM9kIpd3NHdQh
C2jx2nDuXQat7vnLyPnfWAsZmv+1PuuLQ8ItCLQbKiDkfTkXCJlwC5Y6rqLnMbQB
u6zc434pv800xDnvYKLrNRPvpG3KvLr58B397UCUz2ErjCfamzYLSyN9jkNnrCD6
B/8dCb0ahEQGF1lpvw2a0tQfC33WMvrgGD0GV4NfyHqnrUE2miewe8i9QnOGf/Qu
paM05NvANTpTlfeaQk9dpgFBgk10ebeof/EeNXMirM0qOJAhCPJhN14W9U4TiXoM
7onN3eZBkkQhNYpgkScyIlWPZsgES2ILEL36qj5QFnZbxgUHMl6xWNSyvinqSGBD
535orXpf4zMYh9aTKtEiCrBYoKONA3o2fOXFXh5vDYgYBgiDFp5tPLl5w0m04jHN
Q2s2VA+Kqg6i7Ke0xMolHcYBT2fXTBjpedhRIbODpLMqzG5jv/KZm1NQxXNG3zQC
wZ0d56xKUUW2PSWmdn+8ncHVKicjFjoT/9oXF200jv4G/fdgT2nK4CwTYLU2tO2u
qcmdib5XPqeD91t8aMVsBZkknNTUPr9D60YuPL2WRUf92/FX04KsFqNi3pu+R1CC
A+rGoHxVH92+HtJQVLw9P6PI0u11oRlSP/XNvOOyCiXS+UBFfYDEX03zNSm5GsQp
0OmAUI7hak9+YTz89O9igW8MoMVgYNjZ9rUfnzwILIkILw8WoCqbQclkvWfqh9JL
gLpWyGJC0hU8V1rYebvp5I3cWmzJap9qKGhaJtzbjEclUNLg59YZ94ltVmmK+KBY
9IeVNBmM+UUlqpain/gYyk7TsymaZ9lJVJBLAQv/+Us4OSDCNNjh/SvvD5QALlJN
zK/zrM7v7UWpLmJkKDu/1OcarG6vF+GBf7wrsMCYOaFpxe0BZBnnhIXckFDhw6I1
MAwwIhTtjKHw5Es7DcjejmFGdE0l/RxEqgJXBxCZ5NYMQEb9Jj5o4jAnjzgXCIg9
GV/R8g6RYN/nDXleIGzu/CXYr8gt34z2zZwrS6IOo7fdfEwV6jEPG9Qqj5oLvey7
kT8zTIoEFhZZkT6jdYtaZztmP5aiye6Z6Ptq2TnbloaDzhxrlqrfoUF1c2DD2eT4
eIcXYRytphYbceaU+iNjYzLfaPRYCL2VoVKtQdfGsLSM6vvO2ExBMmBcKd2SgMon
1GuyDA4gn2zgaNYYE62FI7/8yeGjeWWSDPK8w8Gs15Y6BTwy00P1PH4K0pKbjl9+
vKWipbkPmgt3ja+ZKJkYenO10M+aNjFYoe+MGtnKLYKa7UsS/eNhtSx8jBV28V9Q
fHQ2pgPPC9Gxyp/y3fT+zWas/GVTZcXSFQVfUZS2PBHwKFh+FQcMeGBKG/1fPXo9
vHDr+tJSHl9js/nzS2Dn9LAnby3x2UXrU/oS56QD2H+UCeVXuVUv3P3r0HQar3vU
huuBUS547rX9c4JvsDh2ile7KZ8AyRVYku1Em7kQBUrd1b+XGDHugxnOmj2h6usE
VamkOmthrm+pIYLTAKsQBFPIsWzPm+xKKg9UK4aOVk/11SxjxI/NiSg2XHSF50nf
VJSXg5tczavEwZhGc8+n2EhR1vZDNebOFRVvF8ifRCWPnRcEpj/sQk4MbJFuqgSP
Rypxng+PxPj7OmVDFm70Px5vloFu1IYZnWxtLqPBcrsNVQ0GwNYfcwweH1C2I8MD
h016SXcjbH1j87544v2S+skeS5Waw8WOIhpmywFbRy8A8AbfkQWXe55KyCau1sen
28h4LBPbUvvwUZftN2O+0kP1c1nu622XanshNkO1HEaJo/2beIuP5wYF9q9DfFLG
dOIsXM47kDnct+Tm4A6lIMbXJ82V5yoxAd739k1fqJQeI0wG53t1c72XyF5h9okw
BhNWlZ1uNLWjFqICVFbBhgzsPCX+BAeiBIz8JPrfuJOV49u06pBAnYRLfBBlE1ua
1UHYL0QkDUZ8hL/t4ME21/tSfGszyI/fabPOHs1KhEba8SVD2c914sBukDB4/QWY
dhz3UpoIq5ukSWXDKNoJQimr4xJCyzE1nnzVL/aFOP0as0ZJlSK8blmwtG60LnCC
90suHvDMG9AXeFlBdm5aTdigfVHBZbRJPw1JaBZTA82Q20kI4Sbtty5iusj46s4C
FGpSeXVfEh1i3wNLKaNn1PIyJ+ZlKz5AByeiESub+Z09Tw6kZW/nSTB55FUt7Diq
WGNThn4bAwlSiBexeu67BmRWxsmvYNsBJpSlV5QWChpHHvfhxm3jbdQDEAQ7odbU
wo3IRnjrkExv/UBAEInLaN8gFtbfmpJ5MWBFWNZBy3y6mKNzNr2THREjRShPnVyt
k9y94J4nLo2t/k1Ui6VAv7Nm2V+5Kr5uctkHpnNciqb6QjFANCG1GSAqgtNQrVDe
EkD6jmR3LRL/WdvhTx1r7t+QAJcLqi6Ix9KIputm8EBBapER4FI/2qD+uwKaP6vf
/qu4foqsaXsF/4hGuQSTlMBBlCHyw2tCOaEvP7HivgVduZtkJ/V48MP+J3qrlubp
EEoia94+Gj7TMvEMNxLoIl0sfcXQZwDhqLa8advuB9f3xwYT6YFNNddSIvPa4zCb
/bRtuDnd3KkXiNb7KZzSjScgvYuh9D+6Z2cwt4CBVc4WhOGsu++P172rmYdjr4bR
r3iLEmjaNf5Y3l2qGelNCt87QcQ7HTZuGtBhMhcF7WlzTCMixtyZYbxpXA5LEOSW
uyikevnj6roHrj5gMiMXflf7i/tgS36P50rrDIFmzpq2TRQTSjdJxeFpKVlr1Txr
AgCPoiHTNBJ/8/srSE8kYgEnKHlGHqvw17QaW12ss6xFO73fez5hAtxiJe6Kk3HN
KkOvh59LYsA4j3Imr+UbE8tIULJ6d+aJrZEgkhqrezKTHKlUgBSVpfvLWK0HC+Vr
uOGbZIQ7iIny3hfyw2q4R+2wVYgtE/YEuynTPHpUa1EIP49Bo2M1GWCLaugFSrqX
XLyIDlWqrtb8FubykUMSW6mu20b6jqZhDzYEbD2LJIhU+GUvi9csS9Bz4qi3alPr
Ghy4x0Z34cFtkpRCAorBY4XCESW2FU48nIQY/ADsciogpmLpnETvE5m3JWEJVNtr
ZwTy9O5u4dOAeJLhLduuSG+kuyBezLZifm5fM9yj5TeELuju1SyxYx5P7/IVanii
1Y1Nn9y9q91nTpIlvHnw65qNjQdZrrog7sQrsog2HxJLfaJt3cpYkx5LFlj/6cs3
6ddKlC07PP5T4pGZWu5kkT/OjDp95fLvENCMvEq1KpwnBxNIaTZKNKs6HqXFzqRL
HdCYFY3vH2C6bG+vwiC4FegCalrs0PV47E0B3qA7eH9uVudiIHRpDyZqNmOnYFey
DrpB4DNGLMJleic9q9VR9isUAnN8Ex+IkFXOD+O1mQp0V1k7G1omx/y2zTa8e+Wd
QQ4jjHaRu8gHmkaeeyBMvaBIavDCAavCHjQZ7W1R4Y6LjlXFfwMmnyhj+5PYuYig
xRurApTie1eCa3peeAEJTZAG33PI5YesidepaubDZtfums0A6QJvctVGuX9rQMRu
+HIrd2Qak1JmYQTQ7qOjbNq+ZLtQ0n9B8wZE9NsCe/vYOYgR1Ck2AU0yOBtdSfaf
HhV9oHUhaWBC+l5qd4aVWpKey/gHQIEpyx8Cdw2ypMiw22f/zG1u/vL5e9m0TB7Z
+wg9sqL0HkNo9H1WyqR5NZ1BiDuCjMLeBg6JqC0qD23cyVFlM/4fPbxL2ZLRvMRF
Of8jkheD1/miylX5A+Y5uGcYvrEEb7MX/VztMEiN3DuOFPjhOuRhaxPy1nADpM+6
O956AWmnvq/Wsux27N3cxJV6AxceCCVE6mJamua2LdxkyP7N5sjzvQjMn3khNU64
c7wl3oDfS4xUVwe/Q63PRdb79Mnob6O23e6Bl+F5Ae8N74IOhBlD9CtuN5wvc+da
T9WKovFkNGUT+DaSQ3W6Ck37GfH0GZt5df84djGRBZnZUX3tHfTU9gMj4BR415Fj
YGJOo7en2Yq4vckLMHQF5L2IO0wBwNjDqpKNfm+gGhrepVnJWoAlmV8Wf921zdtR
VJp3bqfGJf2iMrU/NQ0PYCmLkH4+pmfK8zOosPsJFyRN1QM+9uPmEdkliVtdQS3+
9oftlJ+MOQ/x3Y3AOC9HU9cCmsaB7TgIfXPmnuQ5zjnAQOrI5+iJuKmJWk4wEZwF
+tIGc7bQAJc8KFA1VmLul6o6C7yVNpFcjaZwS645kjguCcKj6HSBmn3sAloUmx0R
26ykFkrnsrom8TnVMwFMr3yn5jXSGuPCfhmp3W0Ly+7ySOOyCOZqBPOChWhcAuA2
nKLVdMZAldgUAy2YYZlURPi/jqGhsdJ8uDQwXPG9ueK/NkTuRLmdnjtNsvCroFXr
90Ha4q2Cwy/vfh+DBl+g8uDpPdALre+A1tN6L6tff31+HoiSLjETpJocEYKodd/Q
71Bzd1Nw/tbBQZM/MD7A8YYLRCjut5fw/F11xUoBqj/6ecjJk3dq6BjzOHttiCZu
FPI6sBWwy4bxhGedKiI11XWLxzb+IPzdcJNpctRjLMe1uLLpVeQ+6o48s3UtOG/y
JJ2dI1ER45rYUuZpSdX66S7UAgLXqqfjMl6MQ8g6XsrnsEGV01s1disyL6sl/ic6
ZNf9eAVbp8jzB+O6YN13AbtWECRpp5rYMx0lI9FqE/WYO+jvRehc4pfWvircDDaZ
K7EXN6NqhH1ak4JKG8sXz3V32vFjo4/i5G34lyJs07TnGY6QVN1sYJPXduzGO9Je
JUappXHb5Dng5R8ClkFyZthnBT2HttsXCT+bRFykwutJsfKwQO8Pbx4ywS4YIPOs
6kwXQb20fV//Fq7nraPkRczp+jjoIjk18KpVY2+/dfC6Ne/hZhZHV/CAKZoNwkAZ
pf9duwotVIJAr1EyZmZjqFPGRlo4YRT+4fbjKBR2uqo03m4B5/+Ad8bfec6XVRcs
4rl3TwtkkV2HBSrHGuzp7pth0uhI2ZBa/4xgSK1bkb61BKIdtW6206Xbv3Os2E1p
Wouw+bWAiGx3iwH8iCVUTQpd7Q4kiaJOFjU4hf8gD+sh9a83U9WR/6qYsejbd0HM
sCdBSYbqFJgj0Abu9esFg7OKEb0fpsFkoR9ar49PBfWApV55z2OcdYNZj5fnekno
Y6LKZeH1ml3p4VAXNCHxobYk8MCYNP42j90MLcRoImiT7bIMsB4o2gMOXPbWhQRO
2vWwnOHLpTByoKRQwNSiSmqfL/DbeTTBIy+CIqsyjxoch28RdOTXphCcRqHBK2+J
S7E/HZ2pn03ds+k/x1YjGcmrWWnHSMc4ewauhtcHzytq0372rJNn80jljRxXmvRi
yDnnOWOk+3zV9ZJBIgbeTyN2mq3yPsxPLNSbl13Qj9ynHdWolQ9g2dNH2GDZZsNr
xBC8wJzh27Wz0DWTJvcBOqjytNheGIeDHL2pM0uFXccxyeNGDxrYPNLQutNnXtMq
5+UoVkxqg3uWfFIhTdUNAdVt504J44NnA+nfCRRNITNnK7GL+nrlQg/us1fqtrHz
Pbe2aENYQxF7B9ln7H0HIBkbi+t93gPCJMKo/DnERoQA1ZOxzlQFREfDaYvUmkTh
M+QXU2oXLt0cHWS/Rh+GDyZwTUwV+ik9QMKQ2Qc8GNEISNjN40IMEncbkZ6xAQrH
mOwd2MG4UY8u9xshh0EJd390M3l+qIIdnzx+y5cVOOUxrlqpMzAMFtfjAiA8wkdK
3G95XMcxSMXJn539CiDnYGtyMKl/VPqOdKy0r38pii6VNYGTsgAD2kfffsSvl0ur
cAk/2wVo4v/R6PBtysB/KtUaxjOtqjnfXvrkhz+KsBKOCpJRLwIT7QBhNtK4R8Ul
GOv6JLod3EtBZx1N9RRDVrV1uDllBZhYaJZIJtK19B9TIyvmqpzPssatvmNZznGs
p6W6y5goYakpiMn6bKBjtXPvWg4TAirOKtIiMLvPyeV8VSa2HSx/Oltd5shmCjQx
EBYfmWVVBdG4maTKHJ4vYduuJGDFwO1Ps7HH9N8NQ4a1m50hepmyVbu5dnaXmoj7
tei1R4MOY3r89pvKbOpPeWdwXw85t6RgxSQsYmUdKRBnkQqbISx42o78ymMaC9Sj
ozIMsPOFRv8S9Yi8+2VyvF/sTX44eRgyTOty6k9BTHbQKLqe1XNa0pwqZ6TUFkoT
wi9ayGSA9gNNY1f8P0hTocfJqjjKNQ6Wb5ZIiVt7VLYeigFEsrj4QSXH1r+NfhM0
gSBlAutgXFubUg5HwKCiAjrzfuxgT5J563rlcOWPHhsf1zTXgqXMWTJVjHok8jtK
OLWkGSPZ75pj6CagN27K76ibi5wN70ILkASM056UN3U/K8/hEPrj9+JcfmJnfnS6
WcPwzPPeoNJfJspff9OW43l09XcwtZMLcTZ5br4dWfk6xnUjCNj9Yshgj0D72FWS
sXuZSMBa2PP1rNafbdPC+f3yBa1Yq0NqOe8qDrKmQFXBKf8Aj5ivzeVPyb7gclht
lHz70ZRYHmnKnV2BFwjH0nmit8Ft6Ac7+bKYVNwy2DUWnD7pkAeyEWL8swYsRq6L
i8oUwjxiuBeFX1oiLrIeTn+oFqpnIBlcckHdDnjZfwRrRBLDrg1Ok3vZ1wZGxAGD
KKv2JxxHhIveYlRVkbZKX+MAJ/HM4kuDQ2HiWaqyycY7aMhK5pBqjmAwY7QDOjMF
j4zeJ6wyXpk0EFMNqyXwvZslS2GkzCwvT0FWTwJdqb5z3rFe2LQGTPHC+qu+mC9c
H5Gkoq4qmrsSEB4mheHE7L4NBxk7M3ZprS6PwXTls1qRHLX+ffaErEwFP4K8t0Bz
m8jn8TI6GJJr0ax971redOyRrzGagq0KhanfWyJFEBsDwH75Z6ckNtA8V5/jAo4p
0UK1Ecx7vQB9bFsbolQCRxUuCRiPP/Ej8NVrYwRzqvtD8EGXnFOSXPW5uegnSe4N
bxiLX5BOvPhXs4UUfp1zN2rZjQSqtjbH3alT9wnuzG/xtnZpv4FX/Raxa50Kicbd
ckBtwra7S74870VEIATnYNzlbwdoKJsKCF4HmquUL4ZSxyocnQ7Kzj3dkRKTXV+A
W3f7krqgS8u7/kzrahZx3NqE4rAbYSKq1Lf5HwDOzs1pZXvoKCynGsIzZOMHD9BT
hZNvipjF9cYKxUSErZvQOb+KbcZEDUVLMugoX1cWBhhOzxtp0ufgPc7IPsKtiz60
GnMrg5mMJ0Y6E1GheAtApR4kBlL/TbrpDnkQ0velILBRG8IBqDFV+zhEt0syWxc4
IUw6TWKXCL6Exmgu24U4nDmDXicgTaKCAlUMg58XJzcVZ3CRCxEX9zF9Sakyw6gH
BNrVzE3/SO7ZA0kuonhsGiNyBZYo96OioaiP6EK5QL9VHnfVp+1wLAYHbO6C3VvW
C+3ro9npQjIHZwscJRNLJIu6aiPFrTPzm7oi/HFhjqL1gLaPsUB1/mjHjM9lOF9H
QCQSY2QPP8MlZsQYJCuJXkku0V8M52/zf9B4pDz0FVzOGhuB9oS4PW9HNSmcriYE
kC9yxo0UDcnfQsALrbPmhFVuTEt2kIqPPpOQoWsz0IVHaP+7ZHAqT8p4BRec+ZMx
UNveON74COOD9oa8zvOfUk1753waPahKyLBs/OPVF12dxCiIR/rU6W43c/WyBizD
hdf7oRVK0byBN6l8i+Je6OuIZd/W+tlkICIXWyV2smWpz4EFRRRLIAwyNnpFboUS
anaPw3QkuK9P39V4fwdmz2eLVWHcSfv2RBSY24ryXM7qNkYSnMFYIeDlbw6NB7aB
hUgkDqX5hfw7oU8VPqMVrsPe+Ry9UuiPgDdyLjFgZnnblT3ysWReEfWwLFvUcRIs
2q662pwExvrJYeZ1NzDop7D9+ZKqCOaFvbIeCQqe0ecbqjwW+os21v8TxQPbTVPG
jqbklaHKHJGZ1HKtDIhBmgXnlbTlhHc1d9xRQHSYGP6qG7pQQVi0DHnDx7ArnaKR
JkMwc+V4tkq6Lp8xcOf6QnsCZqDS5CySlzJWUM0+1nlFEYeIT/tfyFBtA+E8f8QS
JqmtJvZkVCqIc9aoRtFq5vjBmZKn/AUK7pl4VQSXsobl7X8P8tKlkeicmDuSs1Hv
2vFFQw4S9s+I7F5uyVIXRADHunLhyUWVsYBsx4E5ScN/lqCJpZQcZIuc2wk75OWk
jRw1hMBn5bsomogCD/h+GJtw3K2vo4DkxPvotSrSaUm7s1sw2WPz/9Owm3mt17nt
Tzo02ubqeJwvskFO5Xaaiqvya61irHLaJuonMNJgyIQ2b1QzamVmDh9bHmEXCoES
eVAXLHZI3tZOx/pkZqbm/eVf3wxye4lzvycCTm+Mdq59PP6O53K4I2b5tBn9FsdB
pNw6u0T86D35YNZkPEVUK9wgPJ18p5nX7LYv9pO3zLcZHRGbw6iEuTi1eWv0eBjA
Lk5ZUW6fXqsGVpcUP+SmE68TPsPM2p0yh/kp9Usbi/bLJSb2RH6V+J3LuXXsI6Ja
eAB6Ewp1WBJW6jCPAbepYgjYrqXFltc9LbeCxSzQ+NuZRDlpMn2XWcqJQGdbwtn9
49pPrOjb7en6qm8e04R52JqmTogozfKGlbln+EqcQ1fmB3wjekb9U46PqS2mtmLM
cT11g4vI0M69Pg9AW4dG0EBS7jLjdqOwuzd1nZDWq5aXmpPtQ/mR81jV91OvFWIR
TdHTCwxJY8DI2de7avrJrx4/V+ZKUXPIkRcjXlpc3SPdwzzA83sJvyh7DIzxmoZ6
UuFJxvGDy5HOuuzP+tfCKp7sYQXmbpBY1Y79RlWYFki2bawsJUcwiOuU1yy/cqDo
RD5tLs94qSlcFFzET7wmaM0t93pRUPT3KtsPakogipimJIAcgeLZhs2hDX5DbX7N
1eRIUytBjuSfmspd9gzueIMYG30sL3bkHZd39qmHbHLMu6bMmxQKrLbBKlzhfXdI
1VVdOqAIjjw6E+4ZIOT9QEJN1NOOZipQzu6Sx3bUt3uuEKw6hoYI4O9QP5riyzFu
ix88rP2tbHfgw0sPj5HVwq+G8DIf7ewtXlF9LgoN4CaHf4fhsq+HT2CXZxzkocHY
oZdBHu0xlUy3Sgby18V5knCdy52y/L2ZDgwqGembiRLpo8rOVxn839b+ygFzcATD
D6svOQ1bGb0KLZ+EidFo1xS8HJk6IQVXX5UZpRtOGMnbTA7oniqCvsehFoIx+AUb
o17YzXD9XMpcwaI5V8T16b0SlHUN79ISdR8rVgXY284Bgvw+8yNNxazYSvGJpxuy
6zLoThnKRl15nSUTxlCFLq6kshFFnCWf/NnVGUOFWZN987YIcVkC6KP2GOz9iGHT
yP5fQIKkHgVB4Ny7jJ5cT1VtcmBBng33R1hFYecCjIHRKuBObdGBeF98wd3tKnzG
sygS3CqARkk5wckSHf2w+6Zz7bn1qoGUqSXQey0pA4IeIze8aPdVZRCwxJeVJa78
7qIIE3plkyVzmPuW9n4AtXlHAkywibIvoCuefyOXQKhw0ReXD94lqrbNTyjb/ocZ
PjTuVrhgh49HCODyyfYDrbU5Zav5uUq0wmOaqo55Y8TtF+USwyB+Aim9ET9xadaw
KJK49RBqnnMo7m5+utM72KIOONk57KvL7zpVLT1/SLKbFi7dtTiLQv+bfwd8EYGR
XygwzbFxp0VKBmYYvzVrXrbfvofnu8rjcg39IjOao2/AdFEyG8IsDkaXq4aAiNoe
kz+h2SHf7GAjELcBcklWkVNcK9OyDmJ11fZmqPpgRSie2roC0gC7IdfvluRYWicL
OJ19hNe5jKarEtyU8OiV0fFQDIurDtca0gYQLgieI1eyOhGZMuTYPgf7nddXUQMB
Ko7BnccLax0UYX7OJ2pkZOreZMYfxHOS3Dw76OY4Czmq5i2WkUq12T6kStatkuOV
o9i4ZmZjUEX+A2gZqMzsza+Xcfu7U8nJvjkhGgc+PLNP64wFhD4paT3d6h/CoJhO
2ISf6C9Opkut2vKxAL6IQWQPawrNuDP46gdGXU5o6+SQMbmQn092Wyi/pnr0o3Lq
CwJI7E6uhandjg+D3r88FBXwiCypD28AFV4lRrmQeXjRDh89CuUragoqx01QwFuv
N0G7NCmKHXgH+IotCJljXQqy3ZhwS3Gk4VodNo1gsOvIvdVUiwg9ZBSVGxc7tVfB
aY5mjliFSApl1w9HxoJV5s7/G7alsn6iNZMC5t/l6d22mFMeo/0LJnaolav60ggo
+0axvUgP4qDuHLhrVBPTcSQqzDy8Ti/ojSE6VTe3yeqptuYjQZvcJuv4uW63VrXn
xm+f8CEEGLcV03d69hLJ3L4x9YCIJyuyQhbgMBbm1U2xamc01xrPHRzW39XYq1Fj
JSZTd8s9nD6kgxPm+gPlXg/Wz+UMc5b4GLwbJTUmyeBfHp0cS5O5TTVbk3eHN8oF
1WjTjuF+GZ2tMG12owEHY3vN5Hqck6iBWgpBvs5j1oZEIFq7+pVtEzoRXi1r35/U
fBhCbOxJT7NQ53wj9A/Jz7Tc8Ec0tnXGYaUji/9ip8VTOH8jV7OCrGq2wMnMvsVL
Gvn0pYXBGU1xauCidvnXUpAzEpzIzjwDqGYY57vNd76iSQr51y/NbG0TDEv7e1Fc
2su2qgGUoJ8bNNQhTo0zhvZ5dwphMEuEOTzY7QCYneWikkweGKsq7WQWJrpsW2JU
s84i6IaLgs5fDk6BIHPEvMIoLaTgcNWFCX6Z+dHLitjS7wQF/9sohFt8yuFch3ic
OTPlu8vTzi7t1AE2jVjL/zXy16r+FzqtEQdH8Ku8HmI6dc0/aWyUUUQh1aok8WC3
/cDtUOvU7dKJx1OjTc0r8xsqvueOA0qJ01QcC0UbItCDgnvBxJyb6J1BPhl/24Ne
EyLvkIgKNzOcSg1eb1e2sbrXXYVzYzUqNXLYhZcUZQf8pqGcbPUVzMkCfFOahyHc
INr6CUAMYFonRUbOnBR0HQ==
`protect END_PROTECTED
