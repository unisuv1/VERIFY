`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fuR/6kh5C6ItBDpl5Oy1suXcVnIdOvq3JS3kPZKxq1ul4TubAbC7wDdk0xJq1woK
DE1N6KRvryKfqc6U0P4yCRKgVHWp9Yd8plyrvP5KAckBP1ba49RRgeJJPxoE9vAs
Sc/9egsKVdiNDUQmYY1b4yJuRVTGzB58UklFbmO2khXTqxuBPt1GK2jg+g+5eykr
/dn2IIjF0aFeIReHgHADwi4FBIu5KOJqOsrOeTcgnyTrQd6PHWqmUDzbyTn7iBft
REpxcwPeLGlwhGHPhp11C9Pe1BZVvGu3Nz+xd8xo1uGCax5BGctu0kwhU/GY/C0H
YRvwLM+T/xoucM0HvpvU+i3Y9QNqb2isWLerv80YqpVL7dIYhwxNi1meq1LC58Oo
A8LWsoJERj5yskjwHcWp39ORpp1T9iuv+ZDSmzH5qlterIDCTFTbcieRQHcD3j9C
emlAcYT6s7VOoZ7w23urBFmSeWe0kSnX+1f3TWZZZoLpOykfbpzixQw97Qtcwgg2
Jv26p/AZdEVp6uR8dnVBTUgBOL+5luAeMuRNHBNEPOeH3bLfX8F65uxiMjQjxu/m
KtGZlmpHDkRp+5EJqX1ccgP8li85uepDtE2Nf1h6sYPdyyzvoelGFkPQGxtp0SmI
rfwPX8n/PuW9zKtfw7AzaqMAmWlVoSvZ/nUMsELTpAgMlsEbgKljWyatmrrPO/Rb
c34UeqfHsfnoiyR7Sq6cPsaizH1B5qVkdLQgWHs3bNgL3s1LJTnUsAx1/a4NY+mQ
ZS2663iBZ71NMlJiJ0ieHtKDaF/ISZawbHvZ/z75cumYqfWAq8MEHq61V6ze1NrR
PP9dyA9RsLqGRDjckHWGfpst/TYsSRZlKoDij1kOkbxlEHWXn0rud/toY7NtZOB+
LhWQ4/m2Y1s89AItRPtid/paXbqwhoi/YZEeq3y4qcJs5KY9xtOTcWc5cOirbYnS
OTLlYaWVJY1nEuVHpWgFlxJd870zd2lD2XhjbvL+pCT8N/KsADhtE+J+JrfgPgYz
ywQZgL2LQABDA5Vdv32ap0JOYg6qXdXGi+fvkoqVsjc+TktOxhZWj+Ro8bq9eO9t
MN1XvGIBL0QFLccwFM3CkpsR26ldZBqGy3ldv6ZcPOCodYUEYIcuQRVG+FVZ0YRZ
ue7ba4Ppi97B712WxUS3XI4Vx6W9QzUJ01otMd60k8QmEEQagiLI3Z8Ufp6ajWCF
mVoTi9gHSqZ7VvaSQpca+mS5l1tQPhyPPt/RtQdHrPng/ihD6Nd1BpipWZ3zJMPX
uXBrkXQjkOooQd0oH8CppOlgJdOAnME4GH51hJaEXuADX6nzxHN9LLoQYyXgIoOo
BKhp7pmBoRYLtPnaJiFoa2m/D/RPp4jLMCbO35jVozxAB1PN8JvSHQw4mIe5rhm7
Zdkd6+b062W4Z2KyCnz5O1dtcAPGEqGnucK4Fk0/BoeuvjQf8+MYYaWF9TdPkn3G
`protect END_PROTECTED
