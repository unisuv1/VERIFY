`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8qDQJQFrViqTzafPNOFmcUGj85tAtS7x2fkAwcuK6r8vhMC00VQ53CrEYLeebmjS
wqUDlA8anUdKOzjKHggts9MGaTCYnCdxxezkcOxXVbENQK2nUO65AgjZkTM9UVnC
5NjmP8VxzMrZNzxig5pd13HLyPNiBI25QRLTKCToLhUG1uzPBoAv9a8CWq50Fh6P
U3DHvGdwANuQvpJGJblFqSO1usVhdPPE2lNfJ2+RqGzp0DJbKG8BpeRIzGQuYqD+
7SaAyyy1nCU/xCj1wGccboZ0Q/TWr8VGnVZKmMPm2GsGAp66GQedSfE00VJb4w2c
1fsmjOIE1Nl8uYuxwXoCyANrHw6oFwrpc6laF0XBEOwIOeKFF9SuPayHJuYSx3Sz
fceJ/aTIPYLJn/qJSAUGFbvE2pbKrpEgnq9SwlgKW6yBG5pyOUSG01T2vrNvOBcU
QjHH/oSkimUoKJCQVVaN3XGseGwEozG1srLBmOg6iYFaqGnmVPSxOk/ufZZsQ3W1
pOid8x4vc0wXIy58mGcaPVCJ7g9fqvs2O/YPcFPqput9Zp06J/IXmC/maGY1XD04
IrPY6pLf/peHp7JuJIh0Pc1l2pj7wUT1lQ7kp/IuZWGIgCi2sEalQiJ6+ogUoEp4
eeCixRhk7mEueqSl14u0/a4/5PTV6XD6yZWe7V4f6+WZh30zHwpdz8+sdmMfftK3
KL7+eOzBN97ADentrd2NTIFQLPFbbtha3OsnT+pUV0wpDIhRvTv3UoxpX6pohJxH
PNVfPiEIzN88eHTs1Afpr8sTEtTXdFdI75sc5x2DaY8+15OjQD1+XSxVx01MROPj
1A5HNtLoN8fTR6TnVyEXnV4GNrusCRC1IQ9xLmeFWj6TEAptjiSqazA7mraImqEr
jDy03gWROlHQeDwTUMPvzHw1dzhqL6aKYazN9fqVoTQvWMVqceoirjOJycxB8io+
WmEArwkoMLeJ+5uJqgZw5cdMUNvT1K+5ekn8nPVYEFK3b9PhBy7xSOU33JqZMoQf
els75tRu1OnQCBsr9WCP/8hiMIKakVdGWt+P4vONGMu50lTFASFHsqHIKRRbZRGO
v024QpFl6WinfchvdiDJ+xCxMvYTH32Ax2ghZkAoXqI2BwQf0r+3O1U4nRiftyTT
IicWfaQ31m3HyEhww9QGScdLGxl6NMnxylzqZdvi9Nafnn/554vhVjuAxyNFYsxi
8/mrD0S164rwyWSCSZQ1tjtaiaJmTjCF4XR/RcLnfuZfaVgS9Eub5BXvG4Mnb0HD
yqHMDDm7g5s7X7nfgGB5YKMnLOa3IYk96/cVWSg8XsN6XIaq70S+lCgDM/u0+AWI
KtYcBjXxc4lt1ehm3t9zCUfGE4Ou3H+WOsPDwKcyUJHvPpjpti2yOAYRrJSmclJI
9gEbKwdBb1ruPDkW1NWNoaV6Zi9f46GceQ2tpZXgednRdhTb4Cas+SG+aDxRmOqu
kZ170ab2gRC+wQhUtl6l1fROPnDyL2s/DN8QdXDXv6XqUQzum5YvDUmIFhp2o6qP
Zoociw7jsqRHm1OQ4xdciqkAGq4iZdQq1hmLXBplYtZoyMk6SnHirkR1StYQn9T6
TNVOHpsLiZ5w/6+v2MhEnbeROiWk99MuYOkV0Qb2NOfyNbz7s6NFSG8JoktdF/5E
YMNjwfuSMtPOdS3n51fTyUO/1bf1I41sNYkomCaYAwj9xAgstskroFfteZEjSAtJ
9/qtp6UBA6B7Zpemy844Ul8O/8fvErXzJPZcEg26MtYl6/kjI4ydbP4e4fwk1o9F
XUr4DnZDlSFQalBKgHwO6Ywn+8W4AYxwsMNTm0XMWZJhzZkCj5LcODDfeeh7rqPZ
1lrE5Z049thulCnrSqsqEJ/ASR/+rjWgq9EmKa0kM4kOfyWNadmYHERQ0LeT7V0C
X0lpGEGnsi3AaVorh3/AEqC3c/ep5WwT4wby4Vr+5bAtoyzAE1NFIDAovkaPRxZT
JFV2lMYNlqs+XlsfGbgNqj2S4K4HPZU1aq/O+SGuNOpSxUSANfEbArzn0GuLV6Q3
muPd5eJ8KyHTUR8uPOYqSXnL7Q9G/KlarLlO+fas0Zgfu6BHusd2t/U1sqmCXB80
lyll0ozhikeWm4bvI2N9zQnDgo2LKrxXnLqtTLOfPCiJvKI5obNhKNxrGGO2pIeS
AKw+7rbBjg17o19dIlmDTmTSE2NZaCZS/2R2+dhaOBc=
`protect END_PROTECTED
