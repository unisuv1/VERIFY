`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D1FPKHAqzLfw42+u9qwf/oKlElOaBA+ONDpXOuSldxcFpC4rhKYmLjnu9wSp7+ks
BGc895l2peUq1zGYaM9uw7G1X3qocDiohNDeOE2ihVMWKsKTt2qUCvJZN585JtBi
Ft+ktcrpIwandHahtVGTc9U0KWN1G8P2O0JBFZMiVP5kl0AY5HUmgYxXgQoFwSgY
I4VhElY5aP63/hJLP+AcGsc29Fus/131aZNTkqulKWL+rP9zZBvlQU7Mke8qIv8V
GbF2nH7cv2Z5CtGahmPjfI1+99+Ibg7P6lbdAnEGKoJKdLka1Nqjrv2u/gFx9onW
TqeXYKoLKpRk9DD9xB4vPiJ7MaS9PG1NfD/z/rK07S64uJF/arWw2b+7akp7E302
jyIzPLY6A7RIz7SpQZbidvl/YO42JM5s90AznOncqcBS0jFxzlr8Fnkc5UYzMrBU
tVQtJb3QlXNONDSdm0rI0JPOEs8xzztAZBuKvUeJloL1HLKSIt8vY1/QKiCiTgpG
oXrxLdIxCp0fkwzdcY5kldUQWavUGSPkM2facwplrSlcIDDaypnn4jYU4aQHov17
2/vN5TxKQZVOIaKrn5nGlS4K7l5aDKMXvv0cfYbq3b7ViY7IupJ2Ay31uZblKGtK
1rVTYHj9dxndp4eyz43DxkWiEfA/p47LIGbfIdXeQllEfJGFZB5QwNcblzhQuUxa
nWIYT8OYOXFGlZBZwMChCQVTrigNshVA3ouWiiG4qweIc5K3Jp47Pewg/Ojo+wgr
puvWfKz4dMs5rL9djeP4s92mFdF3V3pflBHKB9BvdVhvdrv2JAnpFYUerCPIl34Q
IhGVsha09cVwMRyPjX4dxTNP2piSKENFm+8E6fCgWnK3P9AvsPPGM0/bUuhzHBaI
awPXxwi5uSolcj4aUWay0Q6Q8z5J5bEZgWLwIJcWxTpqgDkifNtl3Zu7Mlij9oPt
6LZGCRO2cFTAdIBXCje3DfozheEYp0aoZlGt6zYk5Cqvl0E+kj2zRwbUF4/3y+Qx
GtjbRclHsnxV/nFiQNjATRtZpzvZdT2IIi/HV1r2C+z9Wk4BrgQriqkq/rcxdmd5
`protect END_PROTECTED
