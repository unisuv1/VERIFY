`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lfJswn5zYLn5/k/Vg3f5X9z6HQoq08KC+L814zcI9p88E+h6W5EWpzJMSblNfP0M
aQTtYbPkyPTQR/9XKNmeh7Al0G54PIR+Rp6uHFNLLiDr40YpSW4cSTqrkcOjzrIK
1a+rfceue7HnetQORB8YG/lA+SAF+jtSu2AKcgN8B8/BsAtcaEYFOio3Qb2yoPEg
gdEQvjefVu/R+ozxoOO8hdXtaohGtOPMESUj2VNIZ2CMc09CN5w7LxsWvJ6f+AkT
aEw3CtAmXqVuTyMgfSpV5jwngOKy7HwvdwPC7voeTYFOPw5q8DgI6bjEQ69i3WB5
EhlDDK+wJxdD5oqvuAavwCA9yk9i2g1TzXgXmWL9QtFym6acoLdMs8VYNiQw3ESE
4nmwB8yXyAaMlQSGgZVCmHfnCq2rMfAGf+CVq62VoA5nJnE/jTTs+yuRHT+fpTYJ
4IDhAlNMqHfZgB2lsZHxfU9175Zp6+ppJQPM2Ix8C9WsKoeMACZuVRXsmmE4/a/+
ExAOBgpMDsCqswoaa8ERF4mdB2O623pQCrnPbknnzRutDgs2GuGGFF+tj689miPK
K+rTux0+X7FpZldg4LxpxzBFqAtVYdSNjjae/sfru1jsXVm/iquYNuf9XRQfCAlE
y7jddlBy/AlwiJkWi86PGA3y6vtar5QVohNBPJ8lZwKkRxRn+6LXEMfGdbNd2jsy
lVU4kERAiNeR0FKwonaMWe85P5z7bUAzTr6u/QWa1KHcriVZC5DUZSREVLRI+wec
GTs73R8FWsTbSApH4YyDRtAXwcfU49UEnfxS95HkmVEWVEHjxYKRCOMY0mn31wiC
hppY8XvlQ+gQQJ0Xm9+cHXIx14iD750tZxN6Ggx0myKRX+61gw/3U3XY4yZKdbnu
Sd6uH0KW7tsxepkR9SRm89iF6eVV4oYeVEwDIJSqPD+TDcb8ZLfnD1Eue8RyVEH9
gTUP9XooL5QYuveejM0aInxuWcuHmfQ//ZU5Kb1UHGc3SrfmTfRNEWybrvao4oJy
ZykGqAd/9ArxspHei2R0x0IzPnonrl3ar5ySEXlk1kGNv7V5ttXof4FAkr99DH+2
/w62VKW9QYIeD5hKN1mVbzOvUzVMARLPLbm48UDi/urx4SUeFYZnyUd541b1lDuw
2YMMwPnaS1lTVW2LqWGGBkDvB93jOaOHpA0jXM5Tb/0CekuIjFwH4tiDqJmIVhv5
VfiAY7xurxjiDqXf4WpncvvOhARgIJUrejngogfMhefwfCXWAo5c1u4ZB9GnGbAl
Q/igP9gFHQgbxrtVFJtCIt0II0H9wnOS2Msld46WVWwrQE041Zde1vdXPo2ZcwN6
fll1gjEtPAJf4vEkSFlTtOZu0FCjpoDxPjT7+yqQeEyut6AEkjBCHKl2T901XdhB
R91QdEMQ5rwCSAoEzFMP3v2G2lLY7FD/CQvjfbx7Pkfn6MHaMJnOOPuZZa4ieRfE
Flc9QRkivW97aqL1g6hEA/JkFzMDukNjl34Kc1vT+bffqHJVCuBcjMfZle5vXOGG
F2sLh4R8ziz5fr0W5lNht9ZA6pndU6k3dzA7DTdVDCg=
`protect END_PROTECTED
