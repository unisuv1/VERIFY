`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
c2AQkmvsRsl5OL8QI6Q+80sQzAKmmRshApi9LQETZi+P2YEdYCd0YB06k3GJAREy
f2OZ8UcnQQ45vhwXUSvlv/Kr+SJ8JxJSDnwVY+bryXxEBJBrKSbbipGDQDWsYxuI
blDR770m1T7JRmSsPWLEnDfgp9BeGqB57JbTxTEOghJN33Cb0/c2NV6RUoZ777hv
xCACF9RmNL/k5yF0DBpC7c4gPtt+kXYq83KDJVTsyS0OUbxTcIhRHDbJMigDp4Zq
EV9/+/mFQtnhsLFL2nDOzNGxVf0U4FFdYHydb7lpeZk6iw4mnfRtEr0u2iAfK+h6
Hxfz4u3PScgKFDI62RZFZhqXCGBBmIoKCLzg6bmSPBMj3DD1Z/RqAxAZKRZ4hCCz
quo3SqJ72+zVzai/K4i0kISuYfpReqVl9ZPDb+rmZZaSOYgbx9QYZnutsNlleAKA
cSYfALpXtdrECfSmIZRbWGTfbAk0aim4NAyCQIme2TAN5abESZdnERiSoYmg43rg
B82zTDub/JFW8JqwGYG5Rl75twzPDkXHJUGYOHYrl8vXzmwmLLdxRtRRai9sL3F3
6ktOLuJFVil6FJTP6re3jNbuEYXVK1bLil7j5pJeW7xlWRtLtHftH2UyqFXS+YHh
QFTAoGbmD0DVDq0rs1uAwNaqdTCyeDK75s7cqz7kGvIi9kv9q2LdCA/smKycn/vA
3xnLxS07U7VbUWzliqWP3k5ZmLRKGB8QD6UrTbmXMaQR1hnyCSddrLpqjbFbDMlk
7QUQcFuaB8TjX/uNOn2EoBkX3SBuye/ZA2TerYXtBIhML7c5rWg5+HGh9FY92am9
MJWza27D5WuniyZKXSPRad+Z5ERJrCOXYJgT86ejgyu1MJkgiJ4+9lhYIRc7H+eA
AVzGz613Tc4VRSf4NvrLxf2PeTywHniR8RphvMWR1p7kUwFzDCmbnAhtJ/72eTe7
MB7eciUi0SNKX1kkBqf6hXoYnL0+0v2NaOUh3KUUzKuJ1etwhe3ygpFB4NWAKzZ/
kLMNZYXZ5AoGJmfUdWjv3V84b1Dwh9EH88bHY6X77DT8a8qP3lqVZ1DyUXK8bswi
OhDQXv2CJJmMuMkgNASUWq3/81iHPxK+JVRVhYDxZNi6Ln7YvnMrruH7G5zDP7w8
y8IC/U9B3prwDGIBzB1DGsM6NXEfURR045mAmM4PdNqtM+8IhOqHFFPDEKdhyCwo
/0MMeIablJRUQJYfsRXp3Fd6r6OKwL2gjT4Z9GXo9N6n3aHr0AjPECsl3yIroxvW
lzdoLbLXVwGrzYtRfEEBz+pBxdqV223AOWplC0Y9Q/Flynt+JsqjCnvrC19V55Kn
hiJDPJranscb7rXxNretPUMciYSnzIac4xxKaRZgnQtyE7u+zd+Z2uj/PHI5VISn
LuwG0nH5gugsHYp+P0ReJoPGn48PBXPtJLhJKC99jslAZYLpayfUPnmbBcykgmQT
8bRW+HP0qq0hHs/otJz3qlaWTCTEwUghbNcStzq2vv/7tFjdpWZj+RkoisjCH3Hy
Hdy51YSj1UVR+/PPGVu7gwZhE0rxzBK/mH8MmNrSZ4eKeYVn00PPHKSZPr9hvp7e
Cgmc3LGPL7LwKgS3bMjlMNLrqvEQlfm7A4BYQoUFaBMuC/ogJGVqjL8qjLM0coqt
ium7864iGtW4Zqp1sYMdRv1YNOCmmvmc02Gyjyk5p9CAvej/kmwy/p/QHq/AcH0h
usTlfjB3ka9SMZXTxA9wixldXj8mZi/SSKImrA8uurffmPHW4wvUh0cGNXgk78x1
6tziQYWZ2QZLc7wvxyEFPdaynCgxpAxedfoP3NzPmIbAzqIWPUg0Fu42cClfehkq
kBtuaG5ayBXL+yma6IU4Ray8hLOv/n2CbBSAY6PfTgpgNb0+k04DfSv7+N3Uzq+w
RH1AEbYwiQ72noWjcJKWZiNncIuRgaAMhGuve1F22udqZXeEZGeqTvf6nFE21/IR
VM9+9A8DUR6JsMhqQxTg9qqDJa7eDwuZE9DJZTLE7OjYs9YL7YSP8ijJl4Sbk/xE
L9EJB2gvVFP9uxPYZEegaN3KgUXUK7zhPT1xo3qT9e+SIfismCN5EKByLzyysDkR
cnzE/l09Vyq8ZcwwWssAZS9r7Pzir7qcHH+J2vIen48uyfLpIz/8YHxtzof0ZSMp
ZILPmvsmth+kFqZH8hiplAQ8L6naDRKaAmupyUWT19I+JQGmKpeLlH0EU06aqmER
DSK62eyXWN8EYKJaZQuFxHq4i51SwCRqItSdikOsuDITNjrqT0PkR6uqs4u+EqEW
eC19qSAW9aapicrE8y8UnqJ45wa15MIaWwHCacJB8b952h0jSfRc04HO/mXOc552
b4hCyHdp1MigRymO6NGx6X36yuhKSZQ59E8Jb+jdPjdwTUynmGpbY7vGC9Gq5yAs
tGyl6PEllpQBKuDsUWeupKLVzfGYGCiAiniYKhJINdwwOFMiz0xYByMQE4SOPPK7
KJMhP6UFOdmjR1M5YR2Ew3ftGlNn3ZFzRWeeRmGUTH1SesxEJ1R+eDJHDHnYtqG7
haLx4jmYsKXHlMDudtE8lO50/aU7iT9bxMazNT0Yoa17R1GiGFlpgBFjHgUkkUA8
oC1moInJb0wLCBY7dTMJ4zaSw9iuCYzIVMBVj2Whu312a9gR/JekhgNRk6zqSFPQ
fDuDDc0swRAXxe8srlLQeXKGZQqDTRu5KmhHUKYV94rc/X9JCd0y9Qi2kmb/QeMW
wbVUQ2GLV2csgf0nRZ2WZGEXykXWexjW5uCNGi+9W6fZ95D8gIQg1sSYAxt6cjj0
qKPMGj9820gXjkN8Gj/p77OqdM94qMxNeuIQO+h8vSzTKkJCzJOfQyWTvqgDRR7e
D7lMWZH8yE3TmHNqG11/XYX3xAXrjOSZ2emoKB4AO0qFKYKlAMEEBnEh1SrOzrbk
fNzFL88O8030LfvnP/Vlq8DZQNxaw4P/k0gHLdXwtJ2CJIFgLh9M0JQSCqLp4LD/
x6ni9hd8XILByLifgHEvF7V3eJO2xnlNVeRNe8m4XTelZEwSDwp4b1VyBBUQsKKz
svSrD9BuqezokLPJ622ZnfslZJz3bhNSo6k8g9uHp6xej0BYMxYzHceXrxi5NE1w
JOcDFz7PlhWHyJFNevIP141oEnpPTwiC7ZRht4U8o1ZFVwYdlq7YjIHlaFD+dMz2
iiEQkwW3yxI3omtSNyCKo12SzPV0iSxzXGmt34z16S8ZmAE0i0nWFCHhwqpqndjB
6YVWdw7XXrRLBPN8KIpGpwk7oe7gB0PmyYeqdPf0e9bR7LeQI+d4EhWrRDyt4a0j
Vh1eM7pcwH9qDfXEJ9wqVFxlDYK5kf/wOD0dnLWI0jOzN3pmvFUsNHgr8FecKTUD
GmkRj0gh39HkOUZzsURRcmcHaaojvWK0RRWO7Rv/q6+O0+Pds2ueTE6NfJHaWyam
8y5eKXyDZ3gIok0gqJ1BZNeacyuIWs+CUKl+doKQaEte1XBC79tviAn9fSfvv4LJ
IAwsoh6RaYr899sEDTlPWSjLMYQJkvEdJW0wBFTP3eTzctLSgjBKUIbU1JrhaDLD
PBIb4wkUj9CgiApLSVfez5c/0KvvupjpYuCKbRRqB5wN2LX3UGbu914ypEw6teIt
XYfja6GkIHP1R0WBeouMnGqXbxBF+URJWK5mJwm6dPEFLeKpXTExknj1OvNtSHPj
UdazMGhg4dA9HhFPZXqwgeFv8nsKWy8V9JdhY2yykmefbTFz7A9sMkykOPR5raHP
mZcNKT4YpbBmT58RpgxP1/s3GCiJ0usFZUMIZmCdQFyUFu5NxZSmu0KcaacDUiXB
tdtKFgEjF3IqSiDY1gxtt8KFOP8mFgM8jfu48PGC0l41EiByAij7ekj27M8pe24E
2rHuzZWNpVq6au6wz9i4P7HtLUETvvdw1rh34GcMc6tjjFPFjj6MEir3KJAmb9dn
shui35k4xaJThjH2zJKIm9AZQ7I2g6CoQobk5KMGS49MVB4CmDqoq3T8VRcQ8Ni6
tSg/QvJpCdGDJxb3qgVpw7GBSVdrO9Epz+nQoweq7rzEBV/MbU5vpuwJLSV62Dv4
FLgYR2/IsKESvSRoOtfoQlNf4YYzgbkQkzssoexhd5uZV6RvgSsmNEoJKNFYvWWH
p29hCBbYSyz24YhTvDFquxkLZkzL547AahOToAX3Nq6J9Euqw+2gtuVsqN+d2Pkv
WcOe1UoHuP1tFb9WWwvc9f9iGJi3Ts9PbJo928ubQ6mMim87DRIIM9VIYCHsdwlg
naakb54Lb+iwST8f6piXerba1flezYAhmjLpdhL/cSO8YO3kPXg4dCQLr1mgFvkE
JEPkBqoYj8QtBPyMJBuxRbPmABWASq60k/YtammiYFzOyfXHtG+E4j7EyBFhTvfY
mhXXBT2+iuhs01JTS9iTBndg5Gwxdp6tj90hR0Mg+JxfCpRUU+QuCJMb0EJQR7kB
QBM8lDNwokPdpNIduY74k+ROPEVJ5uwLOvabn5ud1LGk4Wu1Wd7/v/b7/vfn+aN1
AG0k1qoxghp9GvNTS6/WSrMQXzy9e8aSQfpGc5rITsWINQKgGC3GoJ3c1s8hRwp1
Z7Ibiwx4/+Nn4dZb1svoVYF9vXTG+VaNz7tdZDnWvn1bclhImXP/uVRX7G6GzaA6
EP5g7i4PpG4vrqDct3N6kvtBJN3QrKRm9MKGGoumDZ/bib6VTxewXif9IJtyLVet
Hsz4AUUY1tgduPYFCtw8VQewWHHDR5R1KtyqCsj1bpBTAKbxhgYGYsnPXeV8jzc/
csrkVorPmnuQS5/pjiwEW+zwMOZNb391n8l4Ee3vbxh4Ip6bRl/SOvrH8d8mExIX
fKu/811Dg/DR8KA5ZW7NwCB0GHax/vb/fzovjAMXZXTKWQ5xZXp6Obux84zQYi1A
BWQBvr0DmUfCp0y97/FYkXs+fm2mqi69iyqH1rZlsRmhHHSmwWVz+n0QoRH5oJvJ
V/lG+9X3cVpOE2jZ2eFX7Q6gjhESr6TlN91QTRtoRv4M8tNdIHweb1a1hqRz6u2B
6K6Hc3UNcUncglw9LBweNkQpWzjbsDKBvOxEESPgl9aeCS5MqakutmWUh4XIG4pN
VtnW2ML6gnqQdJt2rbGBxJqXQOsNYbD+BzBS42ixBIk9k6kEl9HSU+3dw9ipatTY
Ng8gs2FCMwLWmYXdrf5CIoj7JPNYN/0+detgTx0jKVbSbCtOqSjn+1Yz7fqpAe5I
OETSy91qRYN8r/uDiC+4n0mvpKffNkMY7Tnp4gx6xmVgxCl+TqViaS0LN80DporQ
F+3Fexv0yAm8S7yM0MgF/SXqgLtaTL1p423HvJ4zcsguG0n4FonpaNjNuVWQqCAA
RnRFMXrZqQxlD9qMz6BawMjK397Sk0Kdnhf1rBC6MbWdxLnPpEbzjmVVi13GxsOX
12bBQigT9cZO2IcW9NYbr1rExUEmOMO6Jir2eMCh0uEMWTEV5o0vsK8fTRlZlrOB
+CpObqH8oLuoynEM4eu1cpNXcyvlo36IR+QxIQe4NY7uu0tnk3Tg50HkhDWlp/xs
q3yEeoGnbD3fY+SioqVok0NrbXRBlE0v5mXNMtq0vXkkGPf0LVshKyYBcm6WxEd+
GYX4/jkh80xDpO4bD8TCveh9uwQSkEv3kv2O5UdkQrtUcPeYbE8dfvcCelcNW46v
WaafpJPD+Mzmyh/kd855daXV4WnBJVewDf9vbpipUCFA8B1Uws7JMqGsxXp7L1Gz
U6ytLyBJt8hkLCeYxp4y7h36/69rU2XmDgZynmvYXGSz2q5ANqU5TsZ/xMdJcFaQ
A87K3/2LLo4x4sPaE3HqTjDvMV4/MdLNTkl54yyHl5RJk4qHbd7E0+fDXQjh6xCA
k6DuL7JVQ96TxZTxMCjui9ZLi9RtLkc/zU/JB9hDPN5B2i/7umDJikmUxeF+hkzR
Atzoq6fwpT4+Svz8fe2RsEoeSfc56dFVR+6f8DTnvLlNPpXsTX+LmDN4Jm/wB5Yu
4alMzxUvCTpa9EOfWagdeC4oARNhdh5CZEx07OROouRd9vu5LELql4OBoy70zSe5
zNcXh7w/as4MMcqXq/YADfZn3Kc0ul/WfmXNN06BybSljiO0ExveukgLCO94FrDi
yVOj2QLLjLYtVo1ccWbM4At/FTRCP/FY0AaGXoCcWVwOkda4oiv3O+rhG7cDWIOx
PKPdy7+EQS+4yIa3YDGm/TaBu8Ykn4qwu3I+m9mpSQZj/3u8DWOj04UKoZEgrFZO
SSlohf9tTMQ1jpKi29Kf73/V09o1XpzyvviWDGEYESIDjDr7bdscYvJngZI9kL2y
mUNWDVMpKe1QPXxMRX7vVC5l4ezUu5JHDUsIEsRjgNFSkf/AwhAU3oTkR3kBen7a
KN7t+Ijs3BvplnUA+zQyhZV759Vgz3IPnu1HgmXHINjVciAgWmqpcyajtRGrFs5U
jRS4VoGZpRMfh6XWM0Dy7s6IT6vGXAvx2eQ15qYEedqffCU5ss3jezulk6Wxbmoz
AzFlIRxsVKxbPC2Q420aBmIRmDIs/oyvJQf7m8YJ9Wsi45usT7ZXpCf4cXXVZphf
J6NAFjSNlqTSZ8qZwpsSRkvDtN8kBB6Fz4hpqJub6wcYL9tLWsTNLsOgQQI8EP48
qtOxwUDnLaUPVSFOhtu/NF61zNyEqx7AMJttGmPr4vlDoAPZ58evTBmVGJU8fVPF
kQilCRhva2GpnQvn29vyCn7koCIs7meXxC3zoneuEArqrDOpzM5RQQ+9rNUNrs6t
Fw3lrZzv1wEXvM80h6kywURXO3L4+abgzVsFY6RSL5gtJ0advx+iBdStCfw6xhun
GZVP92mQGMta/H33/2d+n/MLn+3prfPvky4Jb0kRo/u3Rk9AawTxmF0Q7gV/cR+w
Ok9G/kAZpUOMftJ+rxcq5OcVYtdBm98gb4BL7vNFH49FZeWi/MzN/ZB0eNM6UkWj
I29RjdcsHjueREN4bv82WmjYIw4Ga5CI6z0CWD2iZvJXCyMqcKPAmmcQbwoNdasc
LiQbqrkqJI5kWLilt7xL6TYcGuA+E2ajHlw8kfNKYjTC7bsiIgJ7uRtvea9y3IiJ
4fVhe0SE8jBInW99GDgygGelsZ7bXX9Y0ZBcqhu96efxEga9vHWlj/7nQmeYIH4I
Pk2qlHDWZtV/hAUGEQP6PLmDnYwW+kYOmdag2LUDPfmX4jd6WAM6sinN7im8NsEP
2NY75GBZ6HkGrtwOgWFh2dgt8ZLN9LzBUpQB6WKpzD9ELhvRopgDaxUDAstybdCQ
KdS02OzcpkxAZTGYsVx00AFRn1tYKotRWwqptIurdsDcN0mCZRElTdzLrF4HiuEG
zOOEyEWomdRMm4Q3CMmPB0ZIRr/mbXaW90IPlEtNuAR6H26Baht3tXL2ADr6+sBy
yArKpLUt/txJ46rfzm3IFuso8wMmkXIp5GvB3t7bxy96IGP2OAbQqq8+RWitDtpx
WrPZR39JQ2ZoIzqhEzXvBiYKJ4ujvsS66g9OQ2XsmhAtW0cjetJWaRYguXHoLTBl
4FTROJQhMiWIKb5iWJ+bR6CbXCbFHJpe9sIn3mLxOZyZZlZDYOIBtK42O/Mz8fDE
Uu81aCMGciCb2lp67pUKOQlt0+gCy9OaGkZybQpy6P4YhdORjfMrhBTx3rbBnWwS
qC+aik6C8dZb0a4TsYZEEJlYGQkkU71s3iIafTyFEuR6RfWVO4B9dVZXuYAcHprL
1V+wsB+5mW3qKRaObi3muMpQFG17V7xByoN5Duf1MQIeBbfBAktqT6+YkN6FXO/5
iWYY2Bm1uI/VApNXawArOdGIaTxG9H1qaYuTdfqfV8eGin3VelO+RU4VBydGKVfC
SACysopR/9kygzsE2nUIfmA06hkxaGrKzeP9WgP4NOfdAi7W+QexujwdqXU9YlG0
EU7HN61xToeyJTc6Cho5SyQKf9BQMcwNzpTpSsLFru9IedY0v5PBgpctyjSPPnfU
Ud1KspJ8Xr4jv1pDa8hfFtwhfLlHDdbX9vnksu2T4PqQa5QHoHa41DLJ+2gTUWWh
lOg7iX9LU3xtllPhS/U3ttzhZHChvwkTrJNB7m8RnFvphcRODLttU7Fm/Sx6V8EL
bB8Zwz2kkEAhg8aceKv8nQFFb7LH2tiX+9anaQskLsgUbIwbg2y8rZ3Nm7y1NvOr
8tl9Cg0rjEOJqqrxUK66Xc2AJJD1R7v3rG1+WysqyB4DM7NCIucLM77coeejYSBk
tUGxDUz2nXNB6cBDmoFGryFVUZMAVndI+G/zZXlpdIAwjjta8bYt5Tm+gHATK8zC
MNdffDatNFk1vH7Kvgi7AfhlZIR9P4zuWRber6fiv78oX9O76fhnlfHfB82Zfbcg
lUhLhg114yKF8ZSf7fJr7MHiMHdyu3Ova6+d+XoMZbMrA6weaSTZ4JDT/cgcDRBi
ak9idzbLaLfd8fZeG+ywerC3+2ZZRE4VjnZA4LgPXtjQVhVs4FbfW5Bpc3ERmd+r
//4Tiu1AAW7jOHiS0iTsKDBoNmiEvaiM2+fUXQa18sxwnEtlu0O8E0MEiv1J1Det
qm56LuXW+V3vJkFRYDihy4ALKryU6/0SRlE/SfGfwxUEBT4IDedjjWa6U3vVVo9N
LZAOFtT8irQCZGteX+02UgLRm6ca04z58Bl1NwHkCcrUr9Zq8QRvSi44MGCSQFIA
1SsvIrBa1y/jCT48/TyD0soQ5BOaIiz+j3rE3JhNA6MDmjxVpoo/MD+Ii/j1Gcpu
tVas4wFW5T5P+h09fV1mOeexn/Fnp0XBefRnYQ9HrwCV9/A3VB6xuio3mz3Z3f+f
QabAXJYDOCpk8vNZ60THhnRhFApsBPH5h4Sd3vAybAiOQs5dF5RqFy366ff1RIjG
/13mMkH30MimC/Djsus9xeq8/JkVPeqAI9iIi5PEaTycI7+whkkDh8nP8hvRyaXM
JdJaAmhH6hurDu+PanBXm+1aP9O53GKGc1sPSrSoUaXd3BkGAOppYHZMo8ZtqcJ9
28eNUGshBaAM0qg/zAHQ+hDzYI7tOay2vS1UFDkUre741OwxHrXaD+UXuW3U4a4N
Ub2AEOvRn1kKok2mFH93HjgwzSS2vIXyqQmTzj94nuJW4dTSzx7bPTkF1EZs3NRl
7ocsAeLpOMd4VJRnE6dxvcPB2YLMXmx9KLynDDnXwJMsf9uLW7fBrQf+lCRxmzzz
JcCYflx56HtypP+uAwTOl0AAnCknEjOX3Xe8ZkDKOc57ZT8HJzdqnFH93ifpnrcE
Gd231UinQMhn3CuLBPHrzKyNP+GFNf+i0nOhM0f9jpABCguXdaEBzpOmm1DT077a
JQ4dZULOy1O3vLBeEgnmXoW5uvDrNOJG1fUhfGRTUr/dYZEdhcxsN4ifecyAW/Kk
2PX3aF4bzGVr6fy0BvpqTL4WKcphjKlVF05BIj6ZjdqGAM4vGKapG9vfi/ZwysQ6
wdvZsYtlrqC6MjX6PyXAn+DBZ/G0/F/YZMx7TuNCMAE0XS9ZAZmkJ+e2yXwfMqFk
Nws/EDAGor6I6Jc57lmKBG73L1bjXsCSvBCenycjGCCkBVDVDrl+j0FSkjXzOkY5
LtsaXybPh4kwgrFF3ANMBAbvokXvPOkUjip5JI2ypJJpzCTCryevM+zLKKvGhHoK
Agafn01a3NQlop2ClwVveiE023wpByoTKn68gW57DGKfWsDphqAmG926JZ0AtrsS
5N+Bpz8vhOINlKwYoEwZ+C9F0gcvp9axmTPmVoIqYCfDbVvDKAlYvJy6eioGMPWr
3KtK53el0K7c6oLQ/m/fNUSkqxH3a7awVkYhlALg/SYlu+nFcr0ewwRf1mPYZgE1
U0foaG+GahiFMsamYVNHAAWJQc1HTJmomBI5/S0sz2Yhptjfiu7Ni1kaRdznTr+C
5o0Bltn7yk8r6M0jZrGWApOFoF1phzgXMXSklgMmZc6b5cH48FuHhkKUV3M6dAWC
XVDKX5sxZ+B3VJG4UGwX3L3Aud77udjVgk6wysm0qW/64YaRdDId/8XMiP+mLG+y
hTmytMRn0jTj92z8w/C1hS16rv2tePuKrN7lpgyx3DodYA6UV4tRBLhQ/I1xfFMP
pmVrmYfnZd+biVV58JpKK3R/r812I1Tuj23UvOpFXPg4GTWK/auTVm58ToOp/5dz
BhEsd1Omdk6xqxisDhWR5QKCLDXHT8q6WOOcxtE6cho77vVE1LVDusYqUozXIOL9
CY8RNnoqCE1wqBjYTMKD/AVUBvTYRmLKVb9uBKFM65DxCi+eTqHIQgXx5HIuAqU1
/dLoxWjZKW18fzu+ch5zWcRyPvvqTFSd7DW4+gNlDuiA0GO4IiaYUTg7LH5F7p7U
ldmh83xw+Bqnp/ZqAeIxKPY0+By8nxhd37WlFKoS2uSP5FSS2wmT+oNVE4rxwRTT
ikznVBzZdBOD3gvyatT2NthZJD/p9aNc957vaOI2WXUiKHncocSnLcAdTULSrDRP
cMNiKgaCAvENKw1OGkM1mEOORJK+zoboJVk9g4C4noOsJQ1QuTHt2CVIojLjT6c4
UEcx++tck2hn1yk11OFQx6gY2dXVfrwcC/FEypZgXQ5epAPtLZK6jAxoLVNn15xB
bg4rHFDsVw+FkdeAQw7SHIw4+G65zvGhI/QkUW9wIKjQESxcUeMx5z5t9tHomncy
TtsgQ6T/4Z9mhPDGktmJFIZmPAK7cwjs/5Pj0BakvjFltW3MCX0Ih/iR1aljd9fc
kZCOxNs0QM8i7Q071Dm6p9r3im7QcGxGz0W8d4OYwEJR9LQ0KP+i0tgoxq9L+2WS
olug5q663vbogCQw53c4gUObhxX7KycySZUMbAQnGNNvqM4aPqXVxNX3FbqhhCsF
AtLNck+JXqOtSv0BpjsER+IQuzjmB3UczmU7ZP4v5tzMYh+WjGOwOfmmnCwfgAiB
Bwljk5m3N/4ZKpwoXNXOyZOJD329jUsFEQ7U3oX5krOLw3P01gHcnhu2rT3x8VP9
WNR8v3rynr1WKm0J3OU8BZyA+vw1vMfR/L4ar/KcFZxtyejDsgkGunQJ8s4tcIL+
tMte7zZL6kwOygUZgIMilJudzBThPzQHy+5KsNSMwjDRKHkriqFdlMhxu/v/BOUc
`protect END_PROTECTED
