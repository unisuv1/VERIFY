`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
pT1BdV9zj75jd6fBySipA/BI2D5G4wMP5N0nbPKnNstmreg5Yha+h3nOIO5FtFrx
uTL7Wki6uCaStammpp1K4+XfvGoW6Ec9gwf/bjDNECviEMnuBzVLIOxZ8X2meQ+A
gWGsepzpYiPErM6ULY5S7DJjX8fjJy20wMzWjxJs7v69Y534mNcbao5i2V/+z67K
U1NQMAfdtWbEpe6pfaKlSfrGZH9t9tlG1zp2ryrFHpsoKIlshoO6+usCRg16Ako+
Bt7wQF6pYNhpGeyFfd3NLVf/FXJ2daovfaLvvXFcNcjmq3ZIBMOSHE21XqzKFWPp
o5rmRwsf0Yz7EXi40+4hdxc3fhFIeFdJKx7bcrL16L+oK/1HS9IU/Cy/C234HgnD
atGrRIUItwEVApvtzGVBIIFIehHYSj94bnDB4l0zvUXdnC9pkDXCs19oindXh7/2
dVocATmh143YBWMbvIpgBJemZxG416tqvNoTcaSkuCba2G5d4B9S+2nRg2L+ajHK
xqqY+aBsoWEuyoRvWM+CZD0o3r/28DShJWyYIoWM8MLDp/PSP4zCR2l6dIh3hCZ0
M+xoUiomPHoLr3vpF95mSJK4HquhEQxfFNP7dEOGgJdZvGKNE9lIfxFduNhAnIWj
K62YWEE7Mn/2/Wfh1CWSE9MjOwgF807eNArMbXkdo23XTwmb2aLKO4r3/TjcjXPV
8fULXRMIU656jzhgDMro+izSLhmOJ+0I2K0IHbxVidMGs4ksmPOm5bpbAExsgT9B
Vand39MNvKoFU1lWf8vFAPpfZYDwGMbJnhc43Zg1QMjntRIYxmNZLpFN+70KrZx5
ia4O+Mj3RkKOGPqsApChAzGiWZmmDrwf+/l64lnVxW+YIYH48iKxYzjwmh6gHqOG
96hCYzX6Og6ZWHHknBw2xqll/do8+U8VVwwbHTKK0nezc5gab2UtBDufecIUFHWK
RtSXvAPBqpLvh2yhdmZrXmPc7aOIxeZx0CmLomLMTovVoP4fNaeR/wBlhBDl0/pl
CY9lNunDwCVvxS0ZMVCifuUJXxH9GAZM0luSINgzDZrGw7iSf87nGkqdB2hgv6YX
7nzEde/FNbScTo1Y2vevQhwrS6M9jDuLn9iuNH6RTatRRJzmi4rIAk2UWuIDWYsR
2WTcwt16HZIotn1/L9ZQX2TI9lu681BVMoZ6cr4GzbHDOiFqGMJ8lEZFJvk/KmDf
TF1AjkEeOaFip/Q+LriLRU+6C2KaUnxkv/cc19IdWqB8yD0HitVGtdQ2cwDjR0aW
3RGHX+8tbELqR4MdsLhAN3AyDsS/5kGkusp1HfBwvTvN35NrLpR/x+mirZq9l85A
6mTkbKBhSu9/u+cCSaB4Lu4JIuBNqJzJKCGLMhWHmJhEKJqew2rUVz3ONTQ4J5+S
gjMYtP2MC474OjgvtTjES/eNHOjDVkwYqWV9Ky0T822O9hOwwZMjmFO3u2TvCehU
QKrCDHAdbuE3qlOo/p61Uc9sU48zQo+ywcxAAiVwAL3942sayDj5HdAO3jPpabuG
w5ZN7BXiVZHITAdkhjvpVTWsM5ATJzZTP7NCb3mzw3UUbYex6l380lku4hjKDuJz
lnnpR+DWOJAWaevdfnXd7xfquM8hvDNS518GKSgE6R0zdxYIrRS8KwuuAfqd8jhl
rZ6NvjRMXKjsrYM4oM3RNA7Hd45JeMcx2jCAU0y66IhWNP8lW+8rDe8U+gkLXxs9
S6PmFjF1x/JjIFf/Ra0Oy2l7AjVAlE22y0CZlkMRgaS4LIhqhaw94JyYBgLpZGBW
+OGOSSQih2hK3qq63MZtZZlSTcqEIYmCVLrHihi0RMUPee7ciq+uOH4VY/UIjfNp
8R51K5VTGlB/shUr6h0q1FX+jG9wrOCK94ft7dhu+rIV6x3gWqPpI3GlDpozJ+I2
pPK43ZVnEtZ3KY7JoWuZVMFzc1KzbnbLBELCpCoCXnKrDxGWdF8FPflbUPCseKD9
ZWV91Ju7sFtn3XjBqLVmdXmyoxzS3iDMIKG4O7liQ15eQQOffcUG171WQn1tQyBw
kUBM88nhyXSEom/86wngor5mASVv+6zE64F65whkkzwD/9HB31mNZYPOoHKDHAzw
LkmzSx0GTi40YULoW6TxjIA9NUVaffeIlByF5NXi+Hv1Taa/IX7DdYiA3C7UjXpr
OwsrXzzTiP27d1N4PTQIAH1+HgtHOFo0JPwbW3NPqIUo7/qORAZlYfbNZ5Iqh5/m
7+wcRcySqv5ZMYGBNZfqgIGIJ6eZTcUz+X3m2UpuT5Er6okpxnzfhvCOTrRyezF1
NDH3VwaAl0hnmHP3f2sfgUMMAntuarYt4xkWw/bde1Zso5SF5qr69hftIGDOftjb
OP2jFcgrhySulcan8AWWbhPksORaQMvgP45iub1FAkBXnSKS01zIcosz6HFm0xOe
dIf5zj46dds9vbYWkuqer+5tb9AdxexEWzE2H6vu6JZOd7TsT7+XafwDMb/BdgGJ
0LN0vDGgJlgxXq7uSw9sUuvQAPRzuP3qrUTXcqGohgUiz3aUIoaKPNvA9zGF04BN
MnAKajrrC64FRAAb0KAfdOQbFLlyI6aj+ad8AIIC2vCsud7WveW6HMDqXMSY5HiR
Zrf1mpB6hBhwdbEUPDFFkiDWsLL6MhiRlayrKC8Sqs8S/i27T3dV+v9TRfJ8Kc7E
bZUeKpnqD3vmIFOiahecm1LvrUQgL9JDZFflB14HrQWZYR1Q4JccqSzmwqqvMmtb
DF//lnF8wPSlN+ktgK+JW9xNMm23etbZlLNSXex8rxyiJO50VqMabKTkAPRtdlr8
1Nuwfl51FJ8KfFzyESCZ4OLaMzN7oP7sBngeLS+JsVAamoQVvD+i7C+hiLVGlzxt
H2yzjEqlLZBtaHDjXugI8fY0sLKuj/XSogay37nAOjHnyWFurqvVHvfUzpTYkOHf
pWyMe00AlGz9xuqfH8yaXVZvBuXLSoCASV7T/B0AGELinfftIzAZX4RKx2smffKx
OxhGKifTgaK1rLN232KC1uqgLQ1VLzsEGmpe6yX5iMV0zDk2ysSMS9RiZHw7eAaH
A8LtAFl0eJIoE66Sj0hSzfGB2yME+x+tPPh/ZjJ/I0mf3Glu++Xvtlx3LMdy6Z9n
nrga/5PJcHXBu0gE7RkOL3TTxM5rbNFwp/3sUQ6oN8c3FJIHzNqAtvjTaN8hInM7
4z+P9GIwwGwj0rzPbGWKG26PVzgntNLdA7Kqiav0204uuL8MnrQO3UBW1UZ7JK6Q
e7T4fMEkvt+dfO1Bq0aV+Q9Il1ybvS45RujEgJT8eLk+1TN7xy8C1g+WROKMdx81
VGgYtNIqu+/H30DdaeX1GZuUQDfENock0p5zxqprhDFxzAh9cillwjr37/Oomo1G
lT5sPZs+eCTfWOMrdzToBEplIC4+zyyXH3zmzHbR7qYo1FtkFuoPAucY7Ogs6t0s
vLz/BV/JETuyoCsQf81f6k5St6+kZcE+4MmcF0r3eHXwFVMXW2RFyJXdqnBXSly6
aXp/BhZpR3u8ATWJmiy9b+b6PwlrUA9mNZ16+ItZsQOATFdI4Ia/mA+mBkorin8v
SicVDT+DgcMYRgYTW2R6FH6FgVrFGHJ+4ZKNjsp8Mb8K1QKRJagXLb41DyKQp+W3
iCTvF1tnBcGUktJmPcM3e4eWEjRwVRICpcp3pTQgdKctIkiS/vcCxmlh+axW5i8H
CMapWpWWljLP2A8STjncyA==
`protect END_PROTECTED
