`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Io44alIgd+hKeTIY++orP/mU6zax+vS8LFop4AF/dy4d6s6XtaHASu9tcmt019Ga
OvRwTIYui6HH7BPWd8NvQU5gkitZUKPQdJVPFXcZWCqrRsRnR2wlaplsk+4mDIAF
d17IWqGHcRwYmfrECZoSqYdpIly4NiTIWtwNF9fAYkK/eicZWtmSW+v6QIz60yY3
F4NVi7NCAu+Bzz2KXEfv/ID5KBhqs8robZRxDjzqbFL6QqixFdaxU59mstWr4tB3
N2+NMK5U9L0njwbzxp8Vz69kiNLP4Q1Idu9XOrYvZ6rMomFV/sfTpamiY9n7M4uS
zID4XasD2aH7nm8kPxm46BskCnIhPWQoh6qMoDFQwn7JUiFQy7GakzhbigghggLV
OaIwai/yP2NG6eYJJJGwHtQWJRiGIEoyofCs/b3TO07Ltlb1JqXq3I13+ugLhWA5
aTBW48Ubx3Kh1JwaqU/8UyJe7Zv1mteP+49KXzyT4e3sMbCRIVAPw0NwZFzXDe6F
W2kfROdZABFdCDy8miAlAGgO5IZSizrzbHs5Q1o70bqgup5rn8DnpNa2Wn80k8kX
xtS1/Wr/wa6JCf+YRcHWV/AQCgAFektfWrNZlqP1m4HpwJwD8GUj/iQ41STw9QDG
mtUynV533vj9o8ZDgAaosIRn6+ImXNZGAvOFU/G0VvkGS+JDXBLNnhBmeXyxr0Fd
kcYG/CvLpdisj1PvQ0/RcQrAWELCTx5Bj1jCGbgfVm3/XO/tHx3bc3vOTqSnbZAR
aGm+0ZOjKPFHFFsWFvLLUnmg3ZEQIbJR7gwGKjfrgSGs/OtSvtrqVTuObLpM0Dmq
Gvpu7V+/nsbsgBScG759T0SKlSvayooHBwe527A9Og0z88K+h57rXNdL5uXh8QP9
2Czc7KRId7of2N4GloxcygF8EY+dk4FQpYlBPbpU/aQSnEBdZZLQYiBunL1gofgi
LZ8NrxlIu84ubNv8SiGRI5RRR1jG5nfewDaqsDG6g5r+wmuD48sZWZ42ODG49ovc
GovQ3BsBL/0pU6UNVurGyyPahPIRDCeBtac6IisHDzDjExcPCFQfIuTCxlBkKzyw
BYyqA72+WPyxroTu9JHdrX84JoIHPlvTTt+5fg2WfBZU+/R140/NTqruWq0Rq7ow
IfBiMxEkYn2rWqd1n1ZPgSpms9OycomGABv3+8UIz5L57+Ybns+vkVxDFC7978t1
uDwuBCm/ixOrboBzdNekotVIlG6avZo9S0Y9UKSLKubLJjO5i0fWluTGYUquFIA2
Q2vOKEQUxY+pjq243fH9UwotGlGt7jI8rKtlB7H7d1Xx+RQ9xFf6xOp1Xd60LirI
sGwRzR1CUccPUm3w59RUsrY5LEMxz5aQtYQp/4ZaLSaJ86vozzbd/yr++doR7qFT
VBsOU6amCxXZmhsx6eEkiY0TSoj4/0LbTt18RT902GTrViVPsjE81rlZXAvdiWEA
ueGM9hqP5SVyNGeVqTUDR9NH92/pOfEYQG2L+gxTfV0PKpVxURrSw1Ksou207dua
591RmgjjHu+BU38JkCVnHt2K2Wn2It+Nx1NRp8G8YLnZ+nVR/HjA4q0PRb4AU6+y
lFQaRvdLXGmOEHfdggw3+5XfsHIF8M8paCWswL+iRB+l6KS4LoxM14QRr7Dk8QvC
IPP7puFfgyXWAZUpx0F1aLbexnH8Xj9VR8weWHcZnUZeyA2i3/bAujZMV/fODnuv
4exr7mDeSP08ngW1HakHDDSsRuJzEqoQiXhNXluhqO0WpXLBSP1U4d50/f8xti6a
kNxZ/ArZZAUKb1ApgIV9OcmArVNh36wdonudy76uw0OkWvVwGd2N8DhxoRWA7bs8
pfEHIt8YOT8kYaqOA0gfSAVCVlpnFRkjjVRDk0yQIMxkheImRmgUC7ZaInD7k3U8
q1bUwy4pdMpWsvBz61hs+E/16hlCSr5Y8KY7xzWR/zAqTJdjhIkRjZ7uDpItFMbg
v1z5BgdEJzOjB0rabEPqfsS7hWSwIV4JLEiZOHw4WN+b6x5cRgeNAOtXxR6v462c
YM7NFfwRt5fYfklBRDpE/JI0lSMBSlH3ZNpgRN3sI2NLj5Cw+FF6vJyn7aB9PbNY
DdXuGG8SY1HQP3UEtSvm0O0ERUCxDiVSi86FGhY+kVzcLpcgQhP4yvJo0y0N2Xjh
zAJN3/RiHnKZVFofJyXcGLt08YlX8XX19Zivb6obcZB850scSt4jnIT1Rcnnc9C5
ov3ddB1CpFZ+sVqb8oeEbBBnp+TvoJwhnxvqVur5wwUI49N4Mq3o2fSqaqQU5kD6
dc/mIvQ2WIt3UvJdr7xzsIXXLA8HXbrwTLzsa9Y2c8RWvksAkr6ZX8civjttF8UW
BI8MwJhkisjvqdKmyUwuPePJAEh4+EQyfuAPY1lMpXpOeEb3UgwXkuegsL7KiUZV
fD0h+AAH/8TwytTd6qmRF3leoCvK5/44CnnRdsj26JHgBjmHR7/bxj4G5vVDaTJI
GrZo+5pbAdGNV6oolBfv3DgMqetd+OYu5DXe20UrLlRLLu+Q9rp90GR1Qoqj8YEc
uFHMI+FTCC0ULAkhmegycDY1yGDXiMJnZF4R7Q0DqLezTfdPx4rr/Wd3h9EiTEX+
kRNFnyiqClGDaZ7Rop8aWcDtutVbZDp+jAujA7mSJmnzV9vS41TRthAx3EU1ib4+
0l/aDmbZRBscu0ACfrbWrQRd+2oh1F0mzRW3PGQLSlvUNr7dAUipwNDL9p5kk9Mv
hXqlN4iqvo7HbvzTutJyTaTV91mWTCF69EtNncuG2cJxffefy6ZAmSPO442BRegy
nKeDC0To7gw3K5zSPaqY4EEpUn49drdauRxaV4pdD0wDjaZ4uOA++TPh9uWluurZ
xRkuLDc8+KndmKujxsLPWrE0b+7RuxZoK/PiRBrRTlPNsDO3VWT8FVPGNiCLGQd2
/X68l3AfITKDzBeruuZce7KC5RRMPg77kGMXdqtfFE1QbUsPDl4HasqyRYk6HFDI
kK8QQ4aoBKkxrJgC82wjeB7qJGlKewyR/VO21GI1ZIbCvRmVDXHfi47C6gskeI3N
84Bu7fUoAtR9sqi0+yv3uOJL7IcERf7Tmwrf7jZzczYJvQLPzsjI/ARKhzDqZ8TQ
BNTBOdIhOz/dgfpGIL8Wrk+gOmPv2YoYjGy42p5zN3M8skdmJjf0S/BhTiwOJNWu
evNvzkAbI/rqtmh1oQLDe7xYW0UJ3saWV1hzg51onEofdzFNAuyQnAsa0EwiMFzz
aUPVm86CYAEyyQwQDVNGMKFFfoBL/HiXwlMS8Wp11SBu06QiAptk9Tn1s4tywhHQ
Uefkeueq9WIRP11LzUcRqJYih7+rQdSEV17iPepH3zwWzSiBjLE1mZIBJ9R3xI2U
2q1ACeIxraUfTbCmUwPB7fAPnwr6kV8HYN2LKjlWXxgysACdmCtVRLYsRapwkE2M
CTtnkt+Sine72SMlkIJV+knj2Dmsnm0V7KtHlTyNSzgYpnx2efWWb1G2fsPFLdBJ
BjJBUTzPmW+12voK+F4mnXJy/+8chFbZJyy6zcWG/uFJC0zQESY1ZcBOCb64V3Ap
qLN7zBg0kixFLKD4Gxt+eXLcZpKZdKV5QdUDJmwFlTJxxT+/HH3fe9gqpxZgb341
c1Svftfg+GkuVFeyTGZP49sj72IIO1WHqtLF0qhqaulC6qnFubod3Bx6A0yp8ZZ/
7qMjLVIrSfGIAJGUuNhrkjKP5yHEIIM4VK6cbFDfZSt6RhZahe1yHjW4tRkj5k+x
Qsd3cUuk76dtimMq9U+GsBzpBGjP2rZfJQm0RMQNwyXr8jTodXWwP3/HMJl/uGzs
oiuWtZy+R3JQWMJjdiWwybrJw3pblwj9WQpCFgJngoSHZK5J4gBOYOLfORfCvFg4
scf1oOmLGihOmIQtOVU2KnU22uECRnXe6GpYztmIzSJiRglWi7cxXOlRKsYPjqvI
AnJqJ/OKKdTKeXyqIGqb7E11Emn9CL6q/5F3Em6Esht3o0Fv76CLrZ7vu3EimiK+
dRWZtt34m/sR1muLXkjmsQfAmjspdexL5E0j3l9VmeB+jTg3QtftCL7yqemuRBOP
c/9+dXsa2o8DV1m6c6DCN+P6C6LgkhaW0bFnOo0QhkdWF0cjWRavjtquSYVS2X+q
TFuvUqw7bbGcqFH7EKmFTH2pYzAEXSlukTfaS/jUr2ZNTbB7fl2EA7ERzWKogvdP
iZ+rB+VH9SDhkkPMpwbeRH0pMT/lj7B4Sz+z2omprhz6Y2qHIFhZeWUiHRY9DahS
/yBU2uG90tJfj68sseb8GOnpsmW+13nhHz0Jlt2Qbau//9LW2Mfchc31FEIRHySd
zmT2Hx7NuSnuDkD7RQ6c5wmRHqwmuYx1ODANAgB8EY2cdWxtw57E5hgtwBnG2Kcj
w1ZqKdu1gMHRccPDg0ZEidiCj/r7EljdkPTe3UzK8hXUVlPRa1iIDh2I37P4qxDb
7QdzBsm1Bd+l0uPNuV5k+YseNg8OGZEVEVbUP1QbIwYzePDl5cNOCjpanR0iFPqS
pUl4Dr/QGUgiFcJmwNtoUkRElhg3D4J8ZNX2u8/IfqBRaagU7+xPPgrQiqCQQ5Nc
m6L3XQRR7QUgZA+EM8nyZjohm8Jmz6f+YTh8azuY079WdHo7H23BVzOma5HddFTU
mT6xR2jkgEt4WNSAKpmqtvlBxlqEgciv2xtWtpZHhV6m2e0fMkG++ZFbvRm5LBkC
HDTi1eN7GOLcEYiWXOyc3iJ+VWIukXn5EfohyBU4IbmtembZub76kNyn/nEhcTD3
PSzIpizPlqaAzW6Lzbvpr1Dy1rlRq17k/98/lX3ooy7hBKpqOYk33flCnfjgIyE1
wYKOsGEMq+Wtm7LBY3Ms2aRHpZKs7c46ZH7XH4VhpNUv8YiIJmOKadgfOBe3T8bg
5cqokw1sguLmIPs2D0jPlg==
`protect END_PROTECTED
