`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
uvKKvYY/Y8Y+3VpFsMbCjgbgrjw4B5hIDpGScDSiasbVcc1Q8y6mOTNfomUcHFf+
3VevyHnKOIXVvuzSTNcN8JTN/GfSStc4hcRpX+HvY33bsa7n8G6gVe8m/4rTcfBs
E7nGitF8iQT5dwGF8F/Ww+5YOhroCkgPIw/v3sTEp1pVgC+vbHuWa2VPPekYyLq8
oQxCf4yeSUD44LCGatafdHq6culCSWlEQCdTtnk8muGhCwhzok7yKZvMmH0mBcYE
e78+ROKRIUCEjW++T3jcs6SUyWn06SyccymneAzyC0pbby8kxvDmDWRgy6H9H5QG
0T22j5UiGD3+CrVrXs99hMKsYIWRJsShqPb1kxEuSB4HvAK7qNe2Qf0PjgC3X9C2
0+vJ5S892vgntrE5e0NrY3LajNHRGrae5d/jjJTnEto=
`protect END_PROTECTED
