`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ibnMERg5jLgp6tbZUubue2QQ3DNFcJe7ENqUBirulyjmPnVR2lqvy+2lmmyfe55E
OHPR+JI4XwNvNQPa4QbgzX/qq5dnFrSA+tcdDo1v6dmmqkHG5MihtLh7vY+NOR6I
E8SByn88E79j0nPt3XozfMeAR07tw/WKgf170WfzTgHDbrgBMJRfj2McN3C4QDEb
xgkVElyTWc66+lZmaWTm6ErMxFI78DoaUKyqo2pF4ENSthzIqCCRB+twIYXcTwpB
QIHaDoUaoAH2pLTKIwOO72hPnV1tpjhtZOjjvSCoLx9sQEhK8pH12Igbvko0By5Y
WJxmYyn+96heqDD+BFLeqEVO93hIxfLmqS+P3R5NypjpO7G7bsLYWgjfkU68yQdH
UfJToJHUNkKnxMy+jQafEMqhzwaTGcnH4n04+dSSk5e0epDu1Iftvmcs/HIJB5lw
7qlAAP7dQ1vVjTXif5mr+Ky3QF6qEL73v6rj5uZTagIgrw2uB36xMYq3oWG/pmpN
a33fXOIU+atsHv7CcoPqNEA4f/HPPZ8GZMOSuwzQvc9HchjTXMu3Jo2AgIHzsyIE
N8houiZf65sog2ss1+yMEnu+MKidcNLfphxJ2PKbkczmX4E+2o/6yeTkVY1Z8i9o
PGhKY9QcRdYELSoVNAHDJCUgZAYDONro3pz3/O11Rd78OkKN/u8OPJCfb79bfZ3c
krztL0iWAZxttR8lPd7OmxwBkFpTGrWF4hy6wUswNxVWFa4TGTr11fJAa4WnhExF
pplViFvseFIF7wT3LWPybbiOqaZbgL8iAXPIiCwc915N+4R8X53cpJ0W57L+nC1n
xJBR3sRZkz13BqGR9zU0xnwjR/EYZMVq3sAicGq45qj97cXaK37jjuCdtcSZ2irC
da63/OgiuWghn86CDGPzAxd/V46WJjT1iXBvD4tq+rMYlGDzb/4vN/G8nmCS2GuB
fYcOhjVoUH+eWB1ZQtmiQjOVN2U+54IfmKmx5+fA8gga+kHcv+j/eDHkWhMm9yNm
g3SQaJhmKyjKkiZLu27c/HdvCJneSn7BzqdErEZTtiA/BR5NAyXT+2FVmxGrLIeu
eTJAfpaQrLwCMSucs+RWGcgmUT6yx2+cinbpNj8NGxPlVOltE0I/F6oRBAG68Mcs
chLcUnzJ8Syp0XHoRkJrd7m1f64GiHXQM4E2O9bBWpQ9GAjLyMpd80wB/yaB9jAA
I65WgSd6iCJel2rfVS/i5L3SQj8hSJKeW6LrcDnxq52vpgxdbaS78o8Hr7Fyv281
OLrynR2FI4CPhO2ITM/Vb35/L2TZX7pZZgFsqlX/fxCgfM8/1s2s3Zdl2luMo3Sq
FEfacpR5GTMwp+yLElEX9EWvx4rXoAOTDC0pJHL/NNrP4LxgjEVZBVWMAu2L3wof
BcgyRIm9VCPSYvgve8pYsHI4761GH5iyVguQGxaD9UBZTB66/E0v0Z1n8c1VKQlA
rtM9wkiWdciDWWsFSJyk8lrKMUvbW4EmCLzmGs54fetl3uZEySEA+IvcZk5NKiTZ
SXE1nReTZgyvyE6igonZXA==
`protect END_PROTECTED
