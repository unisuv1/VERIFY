`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ga9DFuDbRV7yHTq0dl5F69NUtAzGvN0530ofKoiveysBPtVJepYpwC5uUsKhcGaN
uPnHOAM0mwFV5veCgoszWq9QELh7GZJ7lXVZAyC9JMkvMHwyqXNYRoXX0LorVZkg
56bh/ECxlcz3+nBDcaFseT5WHWKuXtNWUiR0cTPrIU+4g8jsxp4QjkJtDEpSejKs
pEdZtab8CeFmY0PTG8KhNdkIVo/8u7K71CLhcjJBHqm306SQHPU7l95I0xP+Rsmh
wBACguRsOuPA3k7ypGKlmPkr1JentkdsVcQuZ3Fmt+xJx2bzNignRTaVEDdWD7Ig
qNh578a6xv0tYURLqaBl5qXIFIstV4TdZVdetVqICA9s5oLzE+VGNz7aUFqmapVQ
h804CaHe1FM+0NMgngECquLgW2/hsGXvqPED4lKJhMkGVPGjlCXoMJw34sYUh1vt
Hh52PX5hJ9rX521eoYnfieaajnl4jUC3ni8C76KXrkoqa7vjsTd9XoEhHlKUmqi9
GQ4AArozmBSAcp9QE3VGq6sWoFTxm2qDb8etBYh7Q9A86wmGARmge058670X8ddi
B38D9gYhtSF4frOGzWqOIiHA9BSElvb84fD/DnXSfqo22TLuhKDeOC8eQpr5BSNJ
sGpwszg2wh4sPJqP5R1Z3FwSTdCa7P3QHNAfGbc0TGWwaqKZ5rmzouJDPtLDBabf
6UxchRav/zcwL4oBh+7NjroGOcNVRJIBt11NZHsYbuI=
`protect END_PROTECTED
