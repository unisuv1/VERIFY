`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
kgtzEhmchv+YgNCJRpEVAjpM2olJ3mrKtxUkhWjb3ogEcEbvVKcF69YBPiPbFpFh
HU16DassgGS/UrSzvE8h7ChztC7cyGK5FsOZF1bopnTM5lxO/LlXZTt0b4wZCzUa
zHmWSN+q1N+W1MmkRo/rF3LFgyUJYJc10cpV2c/JR4J3iKrGBLWZisNP3rrou9nN
7UqY1mo7nZivp0lgY6u36deDDqGB0K4mSO7whFXy7C7husyuW1i2E3RmiuNTLUez
dB25ESheIfXSQd1xlwPpWKbi327Q8y8cQlQ/DztQM9vbJCiBRpUaMf7e6Rw8a2aN
LRj8jj7mXVS0Ux2HZOgVvIw/RZ+G3E+Z7uBoeo6fxmLK3q1LIFDvnGAht4nDJetw
cNHSjRXrxZaO6lZTCfZnzMZsrfRV7GSp8BcXi/R/Q3HQKs2DKYZGvQ5BfP2O+in5
4LifHUjjuo65CD+I/HspoG+LHCXTJhE9hy48275OM6N88mD5J6CLUXT+shQF8X8h
3XIQ9l91aB8hqRjx8vJjTbc5L1f9Z3YdITbcvPMi/Tn3r58bXJs/QLK6UNOJCGmv
AtL+GYgFvzfL9ThJAX1XW10mpKk6xhfLNzyiwXqbYTGNvo17SGYu6vXlTUP3En0G
I1EG763XdO4Snrd6NT357dwLsu18tnf1b+AlBPHLNnIzgOlqgKm7eSccoN4jAluW
Y1Q0RlPXEprYOrxy+gnfswVCFIGRAwzUa6b8fwSZmSEaQ1fSKFWSq8IRM4HUseWI
kTQfTTseHxZiQOEWcvTU7Tf+XjjE7xcnRAYuPCKZ1kTvba4v1Npghm2jamMKBTh9
Jq3THqQ2eUI+VgdeX9iwrAWQEVe6DCOhOx01jQW+nEY4ILYtSZyLu4lQtz1YaTnE
RKAF/uxQp5a71gW3/qGW3Ut9G8H0WmC4+c0S05UHHFfgb4PdsMnsqmXS61h5bpT7
c5vp2F4Knv40J6SZMlAy4uiAPXR7BNSnIq5dUTaFtmObnnqsdmVEYHsey6ho2O0J
f4UAnHmGzOtkFklRrw6Pl0YFOHJF+mSKZwCBKZ6MjLlVQ41bZc1xAOaTmkfncDmU
pPFqPxghzBdHIzKgAmR9DyMj6ZIGJPlQsaHjslKAhKT8XqxaAAYiOuleu4CIk+LF
tLKeQTWvif48FXQ6Cc106Dlw94/S+YnCPkXzLJGZKEyV2KXgkncZNtTUuDFri06H
qYHGqreRmYMsB29ai9JoJzgfBDfR1GPOIGASdTWJL72+aRd3vhIKwMgs1apjnHyM
p3iDtFUf9PEDzEV9l/gPA7Y+keDGUS1dhd85joBM5BuF66vliMiQaK2UVYUiOg1W
Kbq121y/ig6dKkhaRFOTmbS5hl31k6FytB6X2/xnGZADB0LSKglGsVQphd8/up5v
59xize7CSBnJYUU3UQir2kU02r5YyknfpUwwnsO7T2WdEtzjVEbsWGJJF1gWtJph
z80/cQKVGaG9Rj7xuN/xE2iW+MiUMBbil/uteRBV0BOWjjbP5UG74UysnOBErTWe
a/LQfdL+5cnqRcAxuzGmBHpJxDuQ7QP5P8QlmG3Dt9AJE/XWai/mdBGDXPNb40lc
P4iPiSwgfoSc9ttcG/QOn7tChcZH0+wnBBHbfBWJRo2kYUG3MKLj7Jqv+kXnRwJx
XTLGZZILJBLtdBsnwYfII1QIgQrFjdiNLAsZjDOuNxc3AX5RFBCqgM2eNKGBpViG
B+7+djBp4x9lb19DZriI0qSDXz5hZ2qXe8fNqU+6IwzpAitLhTHGUAFgzm3Cso47
mpEBIZXyItYV7jaQOKT26pvn1H/5l/ir9a3Y4AbRuksnUSt2gT1Ve3Q+mUkJYj6p
/tnoIsuysuAOrAxo7luGF98YtLRFgPwCYzALcXjELWMcD7BiWMLL+cdfBALCQXpU
WCPdDnqbfW18F3BIlUTYGMuTa5vpjKXJVD93+eZHXBR7LYIGadtgltjhiva9+JyD
YdoUjqKNh+q6lhEC4/a6ccnX+r5rxEvZ8RJI2mYCaVy7heu5Ag6+OauLssH5vwJt
wqXlTVoj9H1tS1q2dxdLWrnIHbcRZ0cDTMJfJPMoAMB8kOa8t5wQC1/AcmruQZVp
5CEIOPRP1bfxpJsTZdHLE5XBbhBBSaKEsqIJgAs5UuQSS0tBw6SqKdJjUthFDCyX
9AcQmBKLBAiWMTGm0FWJV8S3t7joNeZ31LasXr6kynHFJF6q+s6WO+9L3zNzScnZ
lp6OKlyAyuzdykiALmXgr30m/ebaJ30LKqpaSKGmPfPzfUe+A8VnNHGEUeobaWW4
KXxZk6x30nwaZqE/KqzvJ6nWev3KSdCITg2x5bYNFOieb+0hde/IX7/PqIuElhgX
cO7g0UnVpNGoU8QAk462wL4WeL+8VgAQvnjmbCTjckh81w128pst26zr7eyk4W6D
0rIs0HRhe3pQjWYxkOBCmCajJlNL+XBOF4mFuSItYBxOqR3iUzbAYtexh3sfAVY4
mSEXLmqSvvHgqPJ90Fh5B7ltIHPMedu1Y3+znmXaRptW9lB1CNXeAGU7RwCmnliM
1Iz1AuC14S9gxWaDveNH9CAxYDO2yYzuheAyooJWrMEIMVfrH5qFDOi5f3VXg6V4
XB4DXsV8mC1NphhENj5LCwVV9temMXpZgw+7Eu9b3n/OLfyqtStebdacrCbfFs0i
bRy8/OYEsoA5RyD19QSl5KQ0wK+9jkUZv7rhfSbhZi1g2jCtCQ0OQvo9YnwczWNO
y+uXCYt8GU3K9wycwUXLtCE7Ds/PppKUqonm1aGKGqoe4/M/iOW8N3v+zInlMPfw
JuKbjzDxJkMP9359STt9BnZWBgzhnhV+LBW1S6k6ta6mFBAVg4pamFWgkJ4/6ay6
J31cbaHKYqxScuaigK5yVQ2lB1MEcbR0bWtf+SE+/wj5XG2gbZuPvD14sTlAAHuh
UEj5ThG720XynHOfPbc1ilh6WrE5t3PcswRwkJU/XNxPkLkBokPbRBC/vIyCEtfx
4JpO8vbRaoPs4HaPLfMwUwZHrqhfYkcedfO2dEkk4Cw6o9jei7LS0xJjwhxtQM4U
YRBfRnwfnwIRRE7QNBKjgr835h46JWQWgnT+PFiUNCD5LVjC+QKuq8YyovVZUtuB
CqpeIfoHh67YTQelqYnjOfBsaf7UaWSe6VFgTV7mfSCTayfVukJuNTgEOqoUbnl1
3xPG7ogX7CNMpWTnDLG9PYIDYLOalMlUs+0+9sdV6fi+lBbTDGSha2YjqrlpBPkX
VgrL627CAuzoxv2671bEFTvCEdiUr3CdCmKUtlejagDpO5LQg6BsmbqF/cRnx6q2
huNFCMdPJhgijVNE8GVnNWK/CAVPUqFZ7OCB9AshHHvg3R9s/LBa9wNd6OB4QxTd
ZplMzAb4gQ+7kGxYCcglz02D+EFje/PuY8bVoO6rx0hYreCHf8j/ilqeUiMj5ryd
1aYrsNnXYoHCaU5rAGfjdil3dpZTQxwcUZNeA1mCdCGD/C5hP+0cmz9GZFpxhr6G
eD6kHzQHIAHumq/xwFVVBEl89NRjMgbncrhcbsHVjpH0sjN7doEiHoAm/FAeJJyy
ZCWcGBs36XBJttVplMgr14ARh5MPqo5+kwPdZut5J4IWLtAFs+ZHyC95SygEPtTA
lJL4nKltccyaT1Jg0/BJYgzdKV/aTfuU1f4mDkoY8wQ2bq0SBfNx0bVySbR/Ztf6
qKOw3UmjKJbaChBul5j0h1hrdATcwlJRwMLq8KkmN4NyoFYFE2+2yf1d3Tb/aNyw
gjh6xiusZiFcGLxjfaVLW3gIgFES8XMAf+yG3WHGtn7/r0C+O6j9iDpW1OhwIONg
PuvG/EZoeRBR5B6CNAbO3A5Fe28cynrWVd5lVYLmnfsiKHYEbXnqaeO1QTH5VyXg
nQpOvL8M6qTtlCFqjnqlvpaBB/hCVemXZjBQJNB7WvnUkiEd1VgBoeg43bepSlXh
UexkBJuXZ4CPzIyw7GRyCbff48NDrYxh9kV/+MNuUqtU/Bp/lctjMWuiLVadJGUc
AFm6+1Kw3gwoBwqWn2MjPUVtaXFp1UZN+eddaGQh69IEpB9flCJOfJoZajuM87v/
MThcA9bB7xjeJIrTewDAGTdR4fCvGtJOgEwmt6caMUbG13gsmZR2Xb6p4JjpKz47
JgZINanA+mbHFmsNIWmzYeGnzqDP/7vyhxKkxPtYaZ0h+c6SqVcJ6sl5vAlBHN8k
UhCBqrxXFY1XiQSs+hpyhzdgNQGFRJdPyQbK8stR0U2NS9IUOFC0iwLZ2FxEiMZI
bIPEKu1fba47Il5qlUCfif5sVpXqKZqe572kK15EH6laOUIlZv9OqhptrpesEXV1
kWa4iaLk6XDudkjhmNI0m5lS4zd/UpS0Mxv/iyhCRrddI1vkSHIKEBNsZJfAA/ND
ZvGvLuVlPaRrdNuU/R4AUUDybyzWY4IuSMRhpuHYtaii/B0Y9Hdoj+N7Hvxq6iis
bOucO+V8cupNU/RIOMlfd0soloqXdSnuv829j4HbgV+DL4ApGk2u2eNRoETuhtPJ
+TJkp3/fi275eYfT9lM93eY4aF/0vY2zNYmS8zjlANkP0pXjDCel8hccQIskZRIU
khZ1UsQYCA5oZ8H0SjhcRaBGbZObzi42KXzbDJZbHYNivA3xFRqjEFA4ETa6j7b7
I6sThkvXH+sD34PDahDSD2Yqx6A0aPH1YDm0qpGD5zrLrGenJaEt9GJJ0TCc+sO4
Ya7b+DIKfpFsDg74qsr0pznwN6Dw+cD8tawCYU1C5mTh8/k2p0ZcZW5M/j4e+EZ8
IXzWLg+mZbcz07MMiFCM2kkzKyyz1sJSLy9xhFjk0Vx3y3eFt4SazY8VfrN1hZm5
IPxhTMgw+0/GHrDs0vGPSHK+Mo/YKAoFIFeHSmzvJfw2HSDPHiMLHCBwfglPEEVo
qxoQxWeOdJ7XLr+HLVW2mgLM0aP65PNauQVYxymZmkFiqAjOEd39Ul3MzwGcY2+I
QXD5MA5Thlel7xKe6p/0ftq7sBEbQJASZIyvNsJzpQ/isLGU1NATii1D7C/8PMLC
nXJdP+av1iz1j0RI4Sd8q2xDYW+Iw6j4MS+8K70tFs3IFpgqp3iY8om/ItONIQpt
SGdZb1Ja6AgEkEXYSGYbG6bi6orYJ4/ZW79PIk3fsKfQQtigG1nFm3y2MLHBDDKr
3OZpUpBelVDXDbLYKwF3nme17C42mwXBhj7LfYm43eeNVX6YTc0ASswnZHsfaXie
kDT5pHXx171LCw87VvN9NwRgNVGPElvkaOfSy+jA0oMzq2AT2C/XSe42Q2DqZ9yj
5ZFHx4vn7K5s6ht/FmsnFhsHdoCYsQ32V5wG1qJAutBX4ntRGXvLxKvXCsX5Pqiv
/fcFxrBh+3wAetZ/9Zp2Rq4h3KHqo64gbZvAi0k/+YIroNM38ZGdMXOCtlygK3q+
k+j9F/PypjsgCa+HhkO8dTKTgVubZHcLctaTGL8RyY2Rw3LpKdA07jfonOn4adqN
PHw6yw6u6npdq8izHZnifi6FVcFZI/T53sZa/UOfPYwGYOU7pqyjU9P8hmSq61AU
kalPaLDNzHf7J+9OELpEoxrJ1EDSP8xnssO5OWEi+mIpR5a6nrnF/tU/jYQloQmG
jAQ9wDzi9dOGcW+mHV0fP5q1T9lT8A3Y7CIEac2cpUyE3G/6s4b1JluwUTKaS9kE
qgtY6+LhoeVxpU2W3JnhwccIWECg0nIlC1pMFSOYvIfFNpUTRlikK+BUjH5qPyqv
CUKWJ69y3cwBBrN/E1xYDXKP39E6vs7Nv051mH7OhEo8yryThfKp7RLtDyKUZulx
ChZy9pGGySrI+CRdPdLGnenmpscZTfQJDFUrgsCkDPD7uV+wurchLxcanLKzwgXp
God+JJP0u7KflSE8/WBPrYr+bjxzXcdoHXKNopMPyinodNuqqCb9TxZXkMMatsqo
6sXuTyW/rOy21LC3xosYNwaxPaScIdoCAx5IQxfbDmozfXqHu1KlYqMdz500M1Qs
aBnRVmbY2M0gKIkB8a+bb8eVdxW6seMv6YRbjNOo9Deh5ZyxJc0dFfuX4F2FtSJw
1sZhQpKm+3fxqaTKz7Wq9Zu89pqB5OdRTNSPQ80tNuYuZg/oQD0fFG6JEn+LhcA4
dyE6ScGAWAHM9wXHhlfhou4MiFgCGuw4U8nLk9AcAutModFX4bT/Jryq+HF0iOvR
HP1fBs8AkclnYuJz+qtIHXrj2Bq6g1+me8vqghq7f5a+/Wy1klRcHrUJOl5Emxen
FurtOjxYyg4dcat1rj+9aoSsRsdE5JtaM3YmPKm/bMngmDxJn+CW7FZJaRHpjs7C
R1w6KhQxiyO9iPzPw/h9HwiClpQMjtwLzbyw4uhcmC6BGan4TA8X4uS7kQVg+oeS
3fyWNQj+0N4Iec5ikyEXYkU8YQ8rs1J8mUmyaVVchGbghm/dkE/lN3JCcLHJZUXf
c2gF3st7iiJTarZUWKeWYJCofwUh9XWfRClDAgPKo5rnxJuJYYJLFzJtngwikfwM
cJLftwUcEXQmHeq04a8hq1DcbzslxWRIA0YIF6zZ5Ymc5uvGXqNvxc6M9TGgL4m6
S4Pu7SQJz6IYYSmolFITPnW6K3kj6Ea5kHYnPYHPBvGQqXcxw6v4J5VE9LtKbZTk
4/0OULYGVTq5rfwVacBQsX1mEGp0B7YhhEcQ9nBfdX1yuIhv+MmAKJJrZd4rnjyU
G8tQA9gBItiLV1vjWC7U0shanQdl37FuSRjLBw120CiPHsinhOZC0R8Oi9OZYDV9
i5i74sGcx8w5fiNTCQ5/pW1dahHViMED3hSRZ0l95MZSGIrWoDtP1eo5waFHjk8j
cYxuUN2E9yEGEK0sUKbASazr1OKrj2A5vSl6gweD23D2hml2s2/5mnhgjsjecrnU
3HAu8PvNKWfqo3JGq/0OeWZ49kTu6DWJqGJMmXvV7f2bHY0TD3VcCzIxLC9eblRh
hAtmdCCZpzP5Av2uSzaUUVdZN0XwTPk3OLB3yr05NM5uPwlDu4PRph5dJBQescvx
R5F+slClOgFO7YtsHgbK4Adxc91GurloWInfrmtelyFvgcfkB9IADmwibzz0zm/5
ZKAQvQsK5eiShjS4dvUffYSfp6md3pYXxl7e+QzbNCWOIr1ys2O04tAyMotfDLon
hxex2nJ0Dku1c8qqfyIRlKkvgaE4RK2GwAA/QRq8cv6PwFKHz/i82Esl7i2KH6/M
T3IfOkJRkCdK94ws2sFiM3wOgZ88i1St0ldNz9iH/CrjBRpL75UzObX9olUN5YC1
DmksgsTz0RRVDAdSkny/bl65IImymwVCKzodWkH3rvoNWwO5kZAM1XkE+UEYnRyd
l4eZv8SY/gCRym+8W4IaVAafObnDuS6tGTWk7KLvnQ32nxZuHImxvkYSNdjRtHTg
2gmcoyCTVqxO8z07i40C6/TNsur2wnHt/of9t1d6cDF0SQkaAhooGgpJtUBrelVv
WippzbGBZPOt0TzSirgCZEvIAGnBpzZeXryneJ/o/J4eIp3AgWjICiel3kuMXr/J
BCxrQxsDQlqcCUW6xuHeb5AHGn3nSGfZBj+nDApWt/Mmm/SdE2lBxhySlupBfYO4
rlMrCzEfXreD3jHU1Qz8YCei1PuBngnHGwLZdiLffOsIh9xMXhzO3vWC/K/wjLwk
Q1kwmgXBz8g9gmWV1J8qPdvoeC57yK6xBu31zB4vHoxTq/7Hch6osyJO3T/17yu/
X5qmMwoN3cbRzsqcJLHRbYtSQp9pkN3Qf8qKnqsxvN8NF9d0T9MNgZ4/oue12+xc
KnJAYhuj07nrtRpuHldQeoUVqu5YczSCJrbR3KnMaMdh/fM92b1Vgc78duRvEoEC
ervkZp1i/hG0bPzKNgh4YEQgWfPmTxsQr24IkNWH+2/KEy5CcAyA0hiNSkqyyW6a
fQfC17Pc5ZX4DzUR894oPbHqyKuRT08wKYYzifgta7f4lD2STR3Wrwf4JdjI/LER
XYZRdnMgCJKkXaT7Mnrcuf6xofCOv6UblIi6dAxGmhrP0vbxF9+dDknWBJJmLXKI
yFDxlYtJcAd0qbax8PWSs0o+TRpV1LgOuZwlohal+lo3zFzqzlccxgRr3a8tLQFE
wZYprexicZ9pDjnvPKfussyqPSS7+PjohcYCLMerd1T3ZEHVkcOgByssLLvg0Cmf
dZ/NsC+NsYlxKwXdJhkEPocf5yTKH1OyIE29BadWncbzSltBWbCUsN5wTdBzYs0K
rztWQU10sDQsEPod2FYkUqrKmGavrRKdHRtoBAqiE3FPdNMOgPlQ7eT9B9l0/Pum
sLkXXMhhe5zQngNqTxcKcC5oHWR+vfzqr/Q028d/Nj/YRp7kK3g2ghKzIvia4y+H
iNdbVHv0JkyV9dcRKgwuP+ajGXAS9pjBjwjZKrhG1aeuRLIDGtPfH7XFFcPfCBj/
bX5B6PzkBGbn+Q5CUcKOShq5whw5/RN/DF+bE1mNiVtarcVpFvHrPu/eJrvp0YNQ
jasTRPOHv5b8YTtCwpoR1/2zzCEHXzjseZFEC744vmRF1WiBad+JgQPeoBGO9ciA
UVNCy5H+Fj6RvGPqekL1CQ8R+a9J5BpxnK9QE7T8s1C44jyBxuASdfdzKkeLxPa1
Zjlv++oAuqCBwqG24YGUqHySzkNiJJHLTXxR7eZ8ko26H2yx5pDqjO1cnwdgL3rw
K8UgTnhUGUHIZSo/8wGOYOfMmcUClsvifCC20+5DicG05YY0v51kTy4DZceJR3hn
eGg+JWNTxy1mdYI+4d+kZtGXvj72bZ8/kKPvRRkHkv3oNS1bX7MV4u44ikLCdINR
KQMjltzSSywq4qXYsC2J5DFSikpTV+fsGuXko3J2Fdofc+/1AG35bcFeL5A420H4
0dCHcEJWZF8xPmThp4fsZ8vgdkT8AIoBrjV/btQn8UuoyCSdBiZjmHONZW2Wwk2J
oPhsfKx1lMlGBFDavlBi4fxZzUiIMmMDU+MfW6+k8ChRtpu5fblVE3fY+ZXZbG8+
LHlcBY6bEinMbqZRBIYMJK3R4b+jhihVBrVB8XGzuF4FSapPIWfP1dChvtOV68qH
5zIibIeq4huTD+Te3Xcj/lo9z5mEbwFPKxvkq8PxE48dxbgXAj9v5ZeTRDjLQ21c
k83CQUSJ0a98K8cbAepAd3WtS+NLrTxVeIn8Lk6RRbFCf0jwzuXWqVJQsScudCF5
bFxZNe13wOfjSuxJckOu0O1VM5q8dXH5ftobZLj/EB+n8HBpQLs6hDV6OzP87GYx
vfoLRRMFe+8XvRkK7gpJBUbfuGLUahQ4gz06GZGH3A99IEjEFfqctMyRm0e4yzrl
dSuxuqCXiyTRjeEWCZ9RPDf9/qV79cbl1y13ceq5Fq0UT7/dEPcTTXythXbGvE15
s7+R/4MtyUb4y/XAPpxjaYfFMNJ0K4TX/CItTdj1zdM1+CxRykbJjiKpctuZRmD+
tct78jdc83BHblJBy1wsKQshwkm0G07xOnMv1jcf9JAvEEoPuqmfA7vmq7NlU8VP
wsoOH02aIvLgO0RjgROItemHXkisPmRP+1P9JqmB3yF7Nbydcxs1zoNlaljH6qFZ
efwsDW+wUrMUDZQq2npxkOeCvobUN5vS0boGS97CyKE891nsVdXa9YC9ugrd4zCW
Q18QkDH8xgr8ApObvJrIt/cq1wtXlaAj5lYwV8XXfxQb5YoLEqzQTWhw4uNn6wPy
wY6hW2wrzN9sckXSoRsuT2zCeq6oRshKSxTy1ofYEpHSRc38Cyf7DFGmvjMYt9nu
w6L8M2wIkwzVGm9ZrV8ePSRFODq/sQZFRVtJgJ5CID1h7EcpZh7CiplFLz9R22nZ
N/dTRUUeNvNgIRMILhSfCkjb+FI4iBBOklZkPAykvVIUDqafhzs8pL8eirsekJDZ
zkdo5Z6tLev/nH43AQarzjH66BJLh3qlQRXGyoFTxBZCGyWNMIAB06Dy3+cV5eSG
QlrR1Q6tip3L//LUoe9m60hVff2q4XYS+psdcyA/+ZnJG28TqNJ8fMAqTmEGT+VX
ZuRnTzejUzU+39dIMHHa2OSGRDiijNErVleMFIZipCXJELqemYsa3MsJPP7Xeh+F
UibCIOEN3b4+rGpvbV9sNDAzCiyjMo6itcAUauHkDW3GAu7kbNnbhstDAOy23k+U
eZqOytjIJqy90LMETd3clx+K42AxL9x3r56NHJfH5OEtNJQjd2veZBbvEM4d6i5O
t9uthVF4dmtuyPuAsFKZlZ/kJit1hJLMq8qIQIxcyXrtaQZOGdzEX9C39urHF0r8
ekOUEZKImg0HrSM4ICzGQ8qY3m96A0mD9+VBCQsrFw5FMRYoPz28nTXjmAhM1xNX
nbiJBqg9qzLgu0hJC80mMNH3Z6OjPKxpl0OEGoT1d8lhtvS3mADnZ8ctg3iZhHAW
UeSzuz3r4nnre0AuLP2Wp00lrvFLJ4RkJmRtCOejQJEbjZlCwDKGDODK8zWqXakc
zbHKEN7fNIBvixZHTAnSEFjm8B1xxrA8h0sLIbEA21DQbfI648MXCFvn5bo7QFHu
mzQdLFTmJgHQIT6z55ZPuZfTNuULwMGDQF5z02pjLDf4Wz/Zwqeb7+tW0z1KKZJx
7DLUqfAdpWgODERiyiOdvHrcaKB3MG56QWS0FGFrqffYRqJR6odIq8aa+rTesnFz
EqqT4sxM08RdEAGH54erZnpGBdxBolASDgiCagBNgVgmFx8YNkSLKayGdCybkhIn
VH47Og1x427mjCioCGgllCyStBh24t6n6vYkZT36X6Bxz3ZqabqiaSnSMI6rFkVg
ce7I9FMpnwhlMX4jC1Stk+RRct1XjO0tYPqOXT6Yu8l+4Xkesg8qjfqwFDX57iy+
2f8kEMyBlccHjCpEcfrNoFzN2Mm75QPcg8Sc8xwTdFe0zShf/kuOKTMvql1ShXHH
jIzcGebC2QjMYefTJGpEIiuZ3h9Pu/JmJF3o0thWLINUv6BLlOyB3cNS4eDjF00t
CHuAKhxbsGpHYYWS3OOqP7lfLRPlx7Wht6+WxEQqFXwQKZeLRUYNJqAIf52JSA7q
X9zHT7+4IsSYMNCUPDrHDc0zZRMXmoHMb6ijCq5/8SrAd1lPGVJfQKWcnfFRfL2D
y/qfnflH+a0ZzmWzUJXyLrjVKW+3PHZpcTMjW88rXgO0gA6TAt8AeJHLxaTBUGMa
S7HZEHvSw1x92QGkbplof6VK9qeYL9yeJVrMXMWA3qw9aMbek2ZFoS0nw9Rxu2PH
jFg0XwKd3pekF37wgG1dk+O/DY7/cffP21yExcmOlE3Ej0JxzTqDRdzDJEiIt26n
nh8yE2mSXpJtO8pbt42mgXERUQ8g03pwxJ+dTVcAF8c1zn1+SDRvi3RYHLDJspoO
jM04t0D5/Y3rb7NkjP4xEcjHnAxh19M7j9eMdOTFdC7N2kWKD9Cat05A7sdZ68SF
887F6aot5+L7o/kj6KysNLRMZrO9e2tZEjRtBA276vZpAcQjjMvRqa0CcIokL6QX
R0hrneiqBqNe5QRaWPYkD0U0jrxZ7ePNbcmay0Ta153vgrJmHqepL9I8PMKe3eQx
xC3e3oBeRiILZS21VvtOLUf7Krq8KTzzmzAnDIp6iEXjKd6ijLatMzcfw1NOhAp5
o/8DIjfTZI6Ua5f/06LvGT52krJQnaLjYe5dUPrtBa4Nl5IRw1s/USWJsKOrgeSE
5nCkDNQJxegvL1S6VYdXo9dZIhIa2/obyB0oyw7LDd7r4HzZMpXYORS5LtVUtuhP
DVwaZhXzwpRTMDkHHB7wglGTn03xGctp0bmIW5ovJFahLSQEpDCnLFTNmRd4TQcc
uD6ksGI3gMSv035EH/7D8Oai8S4lZMEu/zo9DVk/3a+qqB4ltNt87A9m02dc2eCg
VSjd4BLCj+pZzs5T/AUmWOjB1AtXby+nBRfquoB4WW5qc7OeTji99VCQpM8abiEl
BmJA5xtsQ9Guia1MHTaPHA/6jDmCTa7Bj0DezRx6N3DlPZKYxXfp/nxlt1JYPqMb
5W95Ce1k6SkPmqbFf9DIG4l8OHbJGcbDlEVHoJbufYZpard9wAorJoHu4GCaQwri
qgOlR7wdhbBa9qgfglangJRx3ghVb+x2RwHMQIKypNBkUY2wVqdSQvm0b/GKW6cH
LUq5E/TCnck2acPlWHZuPIYXIgP6imkObtvhQpj1dtid6TAd9ay+hI4o+DA6qL0m
VMhkId43COMJ7FbffFBBNQRmsBEHe/Nx2tVmMW/hWKS8MzDN5066GU2u30ewcKoo
EitWwyxqNDeRMv5uG98SDL+K35xsckC0iKNarPKgJor+wsn/oU/R2XwFcajUN5fm
Vfp+LnifDxDgOka4qfQt/XKXhebV7tFJIVAkfm2WQODhPPuzOWuv4oCuKuKyX1Db
1rNOF1ELfutmN4euMK6CIgBjwcrSOcG3QJUC4tQS1ADC27wwDFBxbIFX0DlF+QUB
0MXjnkf9LV/P8DbSINHwaIDHb4C+7/Uadraq20K4TxRWCCdBdSAapdcnX42mVa9h
L7ckglTQCS0KVuo7LkE6W98PEArtfMEI00qo3Pn3NS5GzY2YE/4okSIpALhjMJcj
9GvyNuvxsRaz9akKN/NhzD2iZALfmw8Be+ygHQWjUjAH9wv3elSi8vGY1pTI7pGH
AeO6OG8waV6LE60PdoAy1zdLdbhdYbT96oATo+Zafasw6zxlNawMqM4jbPZe6ZLZ
W8kQTM8YLNUhxL2/Jpj5vxi715GHIIz6bhLhqCE7y/ysqmuINQ4qs58I2elAFPHO
26LmDVZ60NlALl0qBNs0JZVm+rWB3ovw7VZOqJz/vBf91vN7DZeR2zvVSM4HiuT2
z8wk+m8eM8gZx/8Vju6f/+jrh5Wz08B2i4JYAag6OIEI+yF7cypdceSTPZcGhE4K
1gjUIFfzwqjU/lySrscm7WOkehZbDBICrRiTzqwjRRNug8CoQlKoHrsI1fjD32lG
pfMT3fHfBeBpjMLAwBAZAHUXQtpjgCq8PvbLqBTZzx/arcnScVprEMf3hmrog0C8
UnzEhaPf0dnmu3PhmMvZyi26sCmvneCThI1vfJjDBWyReXROdeQ8brT2f1pX3HBT
w/S5jGgJt1ZOCkiNCXCQUa2JrS1wGaa1WqOBnK3G3FAgeMIuy2BzZ7t+mZFcG44P
bYj/7s1mlo2/e7gYAjsWD8Sgha/7ZkppODbT/+SWDm8mQP76il6LNU1I55bLzBXo
jACeUQycTYY8inUPzRj8WtQV2sQNoKQI895MEdlNh6zutKhmTOD9euyH/S7Qabbl
1abUdnZ/bu/P4wL74686o61/NqqfCT/QSqyRibXcAMOidopyYIRlk+MzVFGsONNc
O7IQPzvyT8VYaaEPBAgak7XYsUOm3eikT3XtP3VzbtCTPV+sdzBAKS5VGGnJqTRr
hvJ8p+uCAj67IAz17Y61pn1561HPgyIvLqnpTQaLawVfbiBedIP0zojY38aH2Wc/
HDKGnBbRkndpaD0CbnymOYB+o99enspt8LSSZ0WjT/hzhxFiYsvh/zzhr4narFgI
JjnqB6KbMUXb4WiIR11RkF9hr0tGE3meQkehR7VEjWsjPohC0kpPtk7cXQRa99U/
DLcxMtQP7DSPX4sinFPa2PeukoC6Usg+Avnbad0GhJMojP4ipulwk2PcJgA81Xw5
EJiinjdvDBA+RtcjXrxdQMqtYtcZwzKCmMMxpsUv/GjB+FZZsMpOvBg6w11z3C/t
agMoMdnau9C0cROxApG5ESaEmLOZtjdD9vkhOg91MFdpQDZVRMzcYnJpzTPOxmQo
Ga7RTI5mq02q9cqPkeVePLU/jMuaR6Pk11hP2N+lZpwdA0BcLleo2bOTBBU/oV0L
KPbp+1gvomUcfa+zxu9HFDdI8F8NjckdDYu+NnUwJid+YvAVgpACgDWg0e3FPABL
jnD3hm+TbR68y9eEyG0N61yIwgZvJuEOtK8PsTqQk2cTT2OAdAnd2+GaWpXZ4TTE
AxvrAh7TMCjs83UX9HhKACMklTPCPCv2Cg+aK29gbyQ4U9uBs4FVPe5iSEDJ/7dX
1t9D9xHTevc3RqTuDTaBdEG952eGJjz1yYenQhFkDCgwnSBJERFlSTtOFwbNXSkG
QmCkFlqcFbWGuQTdEFNaeYSXEbsbTp8dEWx1L49tFIn286dhZFGA02KMhLfSvjpt
yk/2wsbV811byURabw9DLJy/iGH15I+TN1oJcgI5LyDnOGAAOCyv8wXEcCrjrxep
POug9poNMXuSX9674WCwJ1dK+UEtfRBhBziElUkp3HrKSST3PLK386wpYnH036wH
AH+o2k6CpWRDyYLPKa2LmPYql5rbBmOmT9YN4XTODtxQtSw4Cuxe6363hQnWRupk
R4c9NcDMfjB/ONaL0pBVMbIf32jGLxplvlijVz01sLMc3hpqefGS7if4kzt8YU2V
dpcfelZ0CVWg7/BRWJEeVQwBPnyC68dEswmRs8/JIuQrfhVEZssUmZ7wwwuBVa7F
Sbe3kfk/guKmnEGzkMAYnQpEA34J4jG66qvRc1rO3of+DgzGXPcpkF3GS75ICZUv
b/0DALA2FQQQyr1XdVfwS/ft+0+L6iMohZ577tZ73ExGrj7XkLSE+T19Xd3fhhRW
g/KLSqdXay7tOdCK3TF8ly+GAcJij8t3+01QZlgcKRaKqbPzcIoMmmC7hxtkMFMv
avOX9D+CSoxO0LUFRD5Q/lIDLZUNa5aoZa5hEbBvAU6m7H8eX7uyCVuKXRqrengb
UDwD0r/k0vgfuQHzgVIyv4tVQFheuVg/vD/DiZV7RtUnYw5OliggLEjG7Hw0bgZZ
tF2UybR+SeE05rub6Yyd07hwZXhqlCS6SW3ZgEg2WweGx97rMt+MW7tCe/k4qq+i
e8EoXigjDHYPPn5uNdHib9RTCWHdxCNu2MzTFchBTJ6pVsB/fe2RImj5wGA2QmQG
mYhWMzre7AeQ3mSIgIT/48fQ3vjJVDV+shrxmb5lZifC/d4/puIKo6KptTmOHAkj
HlTfvZM0MTLSs2hxSikMAjNhegf0uXD+vV5vx8Ie3PHvoPrz/PUfKvoxEu5TvkIp
PF2RzaB/SdDXfkWeDlcm7B9Y/uq810ucCFTWI85jAx5u8G5yZZX0IfFssEusl16S
msFdDv7NInt5aD7V1nBNyjbeVrEpxDvWiaKd01hUWX2+7v3XN2u+flU86srhTwSb
kYG5VfUdg4ZzdJOLlvyezUBn0PwCTQH3i9qhx/rnGnQLijsrlL+WL3TJs3QfQD+X
bttmVvZCfyfq+qyI/i3zP44MHRtCC2sBtF8zoTXYdssrhTl4qHg1cJOkND/g+DkB
JQuzvH7ngH1ZI1jiZz8di50uEGjJAmyL2NeobdlHOJbFBWeVBsLexCJl6v+Lhkbn
XnAwt5bbQxXGEwRuoLFQoMrwCzAOcHqwnQrY50HgdLnwhhu9GQ+nmw12bJyuVcLK
/8tk7IjGXlmNDGgItYXG4ikjshQee8Va74WfYaoq+sjceVcCm5lGNqNIGa5L9Xxv
j9VdewOC8etns+nISj9PLH/4w9dn9oOR+8NuH9ng1LK1F9TRESCyrBohc1CUJgFl
zjUk9fNYIioHN/4I9iHjcPJ9ESY+OJBupqYOZI/a9nuiEdC8kfQJJ7xQia8YjGIe
K+BShLEzNjhXcrkoQJk9tj5Vj78bf5DHay9FsomijGJEpdvj3Lx2bWY6EFvRLTZf
A7QFq1tVJ9NiWLXP2AbNpWuIUYGCOB0VSLN8J1gZHy5O5FsXvlhu7qbJBYuHEYiW
R2l9+zvxjw9sHEvDSKSR2RFWQFtixrJAJkg2StGvJfM7qjvHiM2trycdaM5sw1QN
3AYSPPxsfXxusVV67YiEycYfbthKMvmScsxHPDYSRAVG5keM5Qkqq2rLhG6FQCI6
hkledZSGTLmjGx0llTjFxpsz6ZwCWe22x5NHkqa4aPH3f5kl2IINDomMgM+k9v5F
Lkn9S1UsZz0u62BCJlFiH9+pwJdkvoWgDg627HC6pvBBogV0i0k7AHFj+XczO/5b
Ua8X7hqNVESGYOQWj/j+JCwBKRGGZ9IogjABazzYK3GFR4tpTFpx0X9J01fmdg4e
9eovNvf4whPky9wZ4cbuvNIQzKVJ751eUGmHsCU9p5k6EJivkZD6bDsf7Pm1IJuD
Ke/VHBdb0dhVAmNx/eN6Yn9cUx8XcShw1XDpqtondBBAADyrxGf3qPCuZlH1VN7k
vLiCHw6GvD9wpmG4Mi4QMi+xXr900NbRdAQPBx8xAEnOyOLgVWPN4GUqAXKtnYbT
l9EunsQtdXGzpc2Ql7nRPnjOQe9a6koL2uE+u7dlsIyyh+Bz908cIf+yd6tY9Cmh
fLpU2/A8mzX00laVv5B8QFa9fibxE2Q2N7VmFpd3GIdJSDfaIwPEBBxpg37SEVY6
JrCAVkH0KMfLJfxdQwyexDisKEOqzxV+bo4v5si9TFmkbv7lLfzAuSkQ+aoPRwEC
6Cdj+Fytk9vYb1g3vTJOv/zhXAPoqGOAP27kST4N7C26h4942yMXFaZXOm6pOy5K
/evLlKoiiHx46CUhhupVFhRPlxKVahbrp+2mnSP95wy731FYOel5USNAPh7EAbQI
CNdwDV33w2mWJ96r6YEEtR77fTSEXw9zuDe7aybniX9CDUlE3U7S9eWgxaF8UTfa
TRpabuA5UzbdOf41V2pilUWsfNxb0JLiDfCw1jdesp5Lm6k6F3dAbx2b+NbDcdUO
WQPwfwp4QKCngExEFc/3I1ABD2FB4V2kdx7qizfzQyC+1Bqxqnf83c8SSSomXKMn
ve35HcuH8e0BEz4/HNNuuRE/GxVvkWjVgwlxRb030ZrlGkTG3MOS/DDDzD/8zVHr
MB37M1yuJl7CP0wenzk2ITCWBF3ooB81LNifPIMKrods287N6qXOZwjwhaD6DNtC
grcMYPKJcylv+vQZ0SlBGfbn61lu86DhpVdjenlYEyYuUU8WAQqslaLN5Gk4lMMB
cJODp9EtjPW2cgikGwqIW+y8PFvPIKM4YrhZJmb5R0AqzR1xdZDDpD6K8pb9nVOQ
d0dkuyD0q2YCoovmp3aAdF9Lu8ubvDQGNYEpp3uPAkTnrU4vvNxcw/GXirJTIuxT
DsiDly/GNnrAXwGNhQs0ecHayEGXLZjfK9pwy4EhKP7wud9Ke+Cmn+XFN52f7U7g
UWxfxpz365esCKG73UmQkwbyCGGSrHrZJ6He35tZWeETFwcALjNmoEPswbCtaWBp
Zvt/rdW/ZjyycHp+F4utVHLxJyhG+1gbpfKm+lQN1QSTBovUg8ICZD+49zNrxEUa
AYoW3aFUCU7Kfx4H+Q/N/9+SlpxaXbadZ5DdADRVY8HQYz9G8zUs44+L7ffglrIu
leDwogQhfSIDMBK2BQwCMEzqXjD4UHwM9DHx+qJg+G7mP3snqBUsgqToQ+g+umGH
0blzBBIhVcjcqjPgGOv96ZYQeyfxS5duDkYdOeYdg39WCvdlepvuv3O8k4JKfwrl
+vTsNNEUDgHUeO7II1hITOj0v+djmxD7rynuc8jRjXG/HuXd7rmrevxLUcOqvsWl
5LNbw1m13nOc4pqy8JNoVEg/qqvxu/b8QApFQ67oBFJZ2bzYmU/UYfg65bwfURLf
nNyO2oYTpO4GEvXDHiqIQjSrDe88tlqvcwCwed/GyGp2IT7ZEfbv//e3nzcLUmri
BXg3U85O2oEfekWriBV4arEDeFgLyjr+f95i5TNC1GdiOG81OEcIY6442hcDsgud
8F3jXlrlTS7jWvPQMARuwvUicM7toJaIdivj19lICAcFaLYALWtIRZxDOG8GHbb9
gHr+FC8aUgA7s5K7qd+umFAwRsLxz0R1QvjyGLa2Ift2bMSNNNUdZUfYeDI6WL9f
pSw88QItT8OGv/zxGLq1h4EhuX66Nc3Tt0XJZ6NfBVHqfjV5pRuRz7/3tgIVJlao
R3NPXBw/5OrJbWqC/NM7pagNnmHdpy092ptbJJYUBcCoJm4mfF0Fp3JOd5g1V1Al
jzahf5O/iXaUbrI8TBDqD4RPZbRgzJhRDzwdLix476fN7CoYRxBEhP/FqdRzsC4w
zDeKn8IS/ywikQ5RGx8zIIqMEAU7QErFatkXTCM0R/fEue3XOnwqBN+bmyy7JH6G
eueFnHeomi8GCjImEGAv+eA7ho9PEaZtk1PuM2Q0YKT3uzgwxVvbRpUoHeZZbEzP
WcwXYJm0AU2Ox4rIST8FTV3VmWiTxwFkx7NJHfBQ8lEzXKBCiCEm6xAL+Z4gKBte
mC7wJbQFIPTeSmj8nZl67lBBlz7W269DTH2cecfSPsBIdl4grl2hFrme7KHfrqQa
FgGm1vzRviedNp1AgoqgwcRfHYPqEf/jOuZH/HdJTpuuZ6FbqhRqsqQ9IyoUj9mC
bdLC1zuMb7bZOcP3ultWiWCDxbSHtdrYsXKHN+iMkMXaTpeIhoMqb2Ys7NmQrR6j
RWWoECr++KWtPPKr/uhaTe6m/xSkcnbQE7agA+9aSqD45zImjQJMUDxv51zYELl8
bywAOQ8ij5sI+2Xe+FQ/gXN+1Wl92RdNbOM4F340ZiJvgL4F6kHtMhoTyw5L8E8g
diVijjaQI6jWqFSd7lN0KgLfRnTeQ4u5YiqFaVFb3cUcZRc5H3QbQ9D4A4fJpH7T
T6qwlzihq62VT4sBczmeCLkL8QuT2kIdO0QmScV6ZlTKOhWtRy7SSXSys99xIXOP
T7aLCq1+YPe5VlBg6rtFA/jRbQLpNTyC8cJy5El9Jh/pG55BsjLnSXaACwB+7M2d
FRBH95O9/K3tXC1g2Jml1HVkpDCgRyTRahkk4xJeAm7lswUtslf0y1VU1CjtPc4d
Lb6RljSMW4RU/JZWXYVvepn8ej6fI1LcdRf30qFuEf7qj3WiATmZbnuNcYHB6nAC
VU2IhgDm338xyOw24a/e7CE2JEqWlu7mSx83b2HHPudyoUmyVSSDKA4y5R4PDCy9
8/pG8vj04KCEIKxCfqcZPVxL8dJETd56rbaIqEbUs5pK1UqBQbGnJ4rw6Xf5j3tw
4h4Nv+cGwIGktbukvsLfZgQxo05RuwC8L72wP1kTnFTBT6/uTeRyzdKEUqMcB7Fq
Pt7Ib7GWOZ0aWgk6AwcdgrX5WbXOjXlbiQU5kbSfuFSB/rW9ZX008pXAYX1ItaeT
UGIpo3tbKwGyDx0zu+ca/JKGaXZHvG+ePLHKvudkX/prdrAdOrS1UfisDAW7wnLQ
s3Pv4JmDbNjRLy0WrII/Yr1/faBIGdvjaQmseg+FyeztPZ8w90lzPkvxTEAhMoEt
psxP+5phPXl8wByXk8HMqdON7wIcZb7/cUsCkc2+D1kv9mKfGEuUl5Ns6+cfgdbs
gtzxoeqtUbXPFSl1w7ByaLQrv8tCIMHxQxtWiFlToAXXuOS/JBdHUIVRa3RHh6+P
hOhl7qcb7gOKicPUHNIYVH/95wPZukiUE8ngY3PK4JX/q2ImzqPVHHDhz21Z3vb/
byTlw+4I+KAmXidByPKJ1cxabQdKUfaOYiBeDCTvBl6XI5p77/YKaG9HW//XcJ3P
DDu8vfP5Rs/tOffae9ea1om4CcOU+ays0HmUtyLggfzUWqLClFbDkJfmED3mifzc
iodJGUM1SttlL4v3sSir7g0UxwxIzm3ipvDorMkyjBWRNVoKHnWejS960nqjUkC6
v/ijWGQI1FunYxD/Ncp2wCMmlQ3fWTig+RBmpEVNYR/hRU572wdsRkEf+qh0IgpG
sGJRbM0fSR3IlT6NFM9B82xstO0Th58r4DoWBGMS4X0X0kLsHNLdnxUNQt3xMXVt
M04kTtg/bEMHaEFinMYFwLKfKSR7/6V1iKEONJw0UTIMU+2/M5lDwzrrhwEMpLCt
PZX4q71QSq/vthe1PhthMXZGSXWapj8lj/nF/+OtrAWkdhoA3OzfuGoxCK2o23hQ
mjtbKixpmlPZcBP/aHSy53y8B1evxE+Lbg5onutw0KS+iFzE8VVI7O7U62fLS6cM
fZr040WdKKQklPw8E0QsST3lzhiy4Ut552v/Puq0VhaUjtIl+bcH8IBB1orsgxci
r7iZPTzZzy2mqUyaa9MBvmP53whGwCT8SylDETRzv/95XYhZOdG0aZO5HlzFe/VC
8EJTGT/sqPRGY43ouY0BexrMTfFy/g0k5d+o1iTZYzoP0eompOHM6XepW34wurB1
I/BbX5KUgixMeF91U+NoEbZc3vIXC2ZodZwty/nLP/ScmumSikaWwcwk7hdqW9Nb
BCzgqcUmdNgcltfMygcLpAbxVfNxVsbZyHBUyGq0tlx1zX6muheoQyScshtMkJ1g
XZihPUnAi6BvK1NP6WHRjhnF0CVpMZ0R7Hih6G+416UtM0slVVLNu+vpRe0no/r6
sz7JCW8ZUt91JBAGKxJWcfR/MGPRFv05jkLkujgC1ldWAMVGZt+bdEv2f3Xzbcbg
9476F1JPrI8gyjL8OCfVqyJvu/3jj5m5ejb8btGSA+6x1cZUBUvJ6+Wpnu0Ew6cw
P8XEm4AMChoVtSI8zSnaUslQMVvQeLUQES5ft20z70AYIa274AuArlvd7uHq9r8z
Pe2qNX4EfLUCbJUYBMXQtxXg+YqoanwU4ufkUZk3PceNQnC7egyDI4FQxhpdbuKY
JPJYqt/I5i5AxkJVuA/qHvJcu5zr2uWcrKx1BmU2Nc/k9tcs1n1r/SU+c7ZzBjjG
pQAE9LtuOocmRdkfP2A864mVYiMJ/GdU+eD7v9QIx8t/Sk1rnqtBb2TpirFBNbdi
1ZdyIB3pY1YaV7rPZdc1AbH31IgxMX1yUCPzGLd2zZs8erjToe+oVV58s4SOfzq/
zU7/zm2QSF/In6GrDTbi1tYUopB66iGZmieMNdykQ9rSmsfBUUbr5JvjRyd5PzIA
IihS6OzySgkkTx0mAkYDoBNPU93cPR2z/3zYuLbHqJD7yC/VBBkAcFYxbFcZ/vAD
+rIVxNFkqPn8ivo070ILqi4RjwEJQjFnIl+jDctNo8K2n3Te4msD4iII0LZNXVTw
rbWyE8VuB7RwuoQF77zqm9xr8JBQCw0unbx8qhqh7+hPH6l3exf58RPeH/D6R0aF
4lqhIcWwY7JrkAp+vF5K/bWOfyaiUHVpkKKMWr2aBxHWF9Wf5gGXzKt7k2GLjG1d
SeL6f74KRIilE1jHKqGdmuntOt/0lSAgcEoRlMK1zcZYH9mYfEuU2P9CsI7MwWkV
1C1YvOMlJY+I9fxLjozzx1C9df8Xc/+s675JLJeGUyT8zt2EwuJ2kFdUmcfJ0z8x
b8gQp/cEu51h7QTM6W6Gb/3VYgA2aNsL0QKehVObJZxSBhpASbHdsDZp9mQa+kvQ
hX1HZNaU5jjY7Xq1S+tVSJtm955TOQqAu7vEkj1jY+G900AsuIzcnWbAgCyak6Og
ZJR8upkxC1OGcDGbQSrDonGV6BkYUvStAJSGh/eq+q2i9YPkofw1PKpxy4y3zFOX
FxQf9vZOvbOBGChivWnRnBb89MhA/B6ANi7wIzgnzcG1YHnT+Mf1wfZZ4Y0gnUmv
1ApXSmyUeK0oa9+pp0QJxsxtvIQDcvBo0+tZe0lLJlwMDjcBFOt/PQtH52bZUjlB
J2mtkAxF/5pKBOH/C4oJAjR6L+srn7UicXHWGOPAdG7xYEzlsfsNVoOYUVRghGmc
3xs6tVLmroNxemTTWLuN4eZm15B+ir4+phTJolLnMJHglSmKzyvaC0U5XMlxc0Ez
jeC4rFU4iRshTKOJLGtqQnnI8YbRprpBqvd4Jl+Z5wAkvB5bQtYECQzAYUHrDLv1
P/lOHhS/i4OLSB/CeIKVfFKXDNAJb9ge4u05TTpnSMw6R2qb9sHcTSWLXA9zcHm9
7I0onE2pqf+bV9OKRPAUvoCUckYpHB7rTWWz4enhyQW6K5mhj5yiFrYQx6il2PU0
IbBrQvp9MYJrmwTx+dggIm3ijJM6iV0dH878uPFj+psz73cVU4NLfR4Gpn8+87om
cDh1CzIDZpnnV9kJdmzEUsi5bRhXWvUJpmdM62Clg5wXPVwUCyKu4wrxZL5RtGBL
MJhDq251z8WViogmlboNekB3TyTFdBIhlXqosDuxQzd6MBxGsqjGpPQgb1DPgyEb
0wvvXymzkPrC125RKuumg3V64XK3JebUNnnIQmhxPtX7VOPMfRtEQeqO/m4OKTQI
HkZN/5cjWMON69HpeEFi2+gehygkIaCuCH5WCmMjZfA4wk48LSXTUwfTGfrH825c
57PYw2ltG2xvx95JjPFshS7Ta2m4C/AMn1sqNbHOXQDoSghumBK1ufo79dJ3twzH
pXWVkhDEbPj9V83oTRzwfsaf9OS90RvpthBI+0yyInzCOodND7FdT7S1fKtG+MvM
MPSFAr3W9v21PHjqXZ4/TXzTRaNxtz3JzUXyPMEmOzMNum/xPJaWxToMq4wOnRld
w6RLSTEM7Rc3Rth/g0AcCa36C6Y41S+aKmgNyIcI+W7kZ4wxPHDCv9ErC/gcD8XB
eEwjWyUij/HgwFtk1mYRdp5yrOLC0GTA+xqx+fSsiLj6ieBD/70mDsmaBjZqRFsX
7g4ixW83LsAmMHDummp7EPLMEVE8NrkzO1zbGL+ZfaaOw6DXbBaShn1aHP/V94X8
qfW0WFLtYAF9vAvBqJe3y+TXAwN0VXhTSDJdxIDVJmNBUKnTt3eDM1RE18fUrkl+
RCHa1xXwkLo63k1+xOq1qX12S+RJgNrXviJuGv3UyMXgPuxA+Kdi7rU3SeetELuy
SkhI4dx1oi5AV8tjNAMoYczMvS3fAUgA3z4xLUoWI3m1vNBsNnekpCtsp5oxeaqj
gnfblGqTHJBQB0S6Q2Mh6eGGgh+xEibrR7IwI6cBsl0eVmtBYl55vHBU71As+kBM
WdZFghAJNzv8ylDLfMUE8xxjYNC1N1/ivvQ0jqGXadZCv3VQGAg2uLNbMYdL25+m
UQNsT4yBltjboOS0rAqbapPtUoW8afOJCSPVUQJbJJZJuby6c8npcjaeaeiPvCaf
+RuTbsbuNOzOiADd/0PFkqrQXoAt11BiChzGnOPc743j2WrlBxiwz4pr42oBVn0y
C5HCwwYQ40ZVvm4ozzhIAMADLtNindLY4lMOnKf1oSpDW0mv8z3vbnG2zdCH6Bdk
bYNneOj5AmY/E3+YAO6bJGpsLNVB2niAJ+iAI+Uz+WxCkpXdUAlkESMfKmNGWPrk
TC2WHj0aj4YS0dI8T4CTLTWOAXwGZUWTB8ftr/p9wBB1MAKSDie3ZEK5jOp8co2p
5f4lnc9reKKFkHLpAQJLl8P4bMANVWcS7XTiGQSdwKSCSNgLXyJ0czQ0wRUxOJQl
quyCXqiD9nBU6pxmH2ybuWARJ2XKLs+SX6t0APGlukyzyFOwUF1oxtLS23w/J4b9
2d6mzXi4GBfFbhKledaNAEt/uG6pBhs2/THX45YweNs3S60Z7VWmtzyOwmy64dN2
RkL4Qb5jMkIrK3tovL0As0lq0VSpxir8z0voY37V0jA4lygmiaPRa/gFRM1vungm
iwg8iM3TUBl1W9Nw65lxPHbRRQmozkxWw1gSYks68SEgt0wuPsox+C3nzhfovHlA
ZEyJscEX9+vnj0ZiGh9U2GYpHZPHgAHLsFW6D9xnmKhZsLVo91/4qOMVHd0wbv+7
vWZFPp+/64rvhYsqPHbuzjR1SqyHXPSKpvayVjtJelHJ8Fs26XYHGo1Of+8+65JW
/2vwPbKnE5ChDkokGuGGl/dqyRAAT4HltYR37p4VVqLyVzJ20ElfhH1JYUJ5kuGL
3uK7wkx3VPSRnOzDvHv3qQYQqwDchOxDU0E58sCrrabR/ML92V3AUDzXmg/iVHwf
WQ5LdA/gmBcEwduxD6mmiTCmwnYpETQgVqni+OYcOYbFLmCV0JiKrLqsHPxYGE8W
S/7yfqwhrNas+OEy2AFuWt0NdmTuF8FqRWODkqFiDZsjggdVOdLz6dbYzF3Lneae
JZVzn6rZe5KmRVlAkuKupvVDmX3+cax8aAimdEk8wWOrAbNMnP+Vz7L+VK0GHcMA
vV3UWsHoYGi/pRb12Shvf88Xe9qEIrXXFas23sMQx1H5nqcPrLdfe4GwaB8kHCJT
SdaIcGJ1w3syAw8Q7gBtQHqMYqEtIDgSn5gUsLQcwd90/qGoYG0+cJvsZzS0UZAC
V9j7FNwdFnfi+tcCyrkjuGv25gwCh1M58ViGsh8JEymHBHo4Djb61bk2t95nxINz
TzJwIZzU/tTexwzxSCArYhG8/yV1iACxUgytqiJyee/TDGMDweD5F49tdHBfH7pB
5kJWf259OIBeNZ1b9fO+U7FIi2iS+u0uLgQL3xSNnnZAuYhNniXGpXIwKNwO+a3n
fcRqjGozNayJ3lcZJvDeNgTAYkB1aW0E0VGg1wwq0u02tUhKChB/fcHbQeJNq+ve
RW41cwmqaz5EUSpGhQEez4FEICe2hmlLdXSFjMN2Fx1x3zJprWc9gaLeJa5aJ0+U
WBjxAfBOwFT79B9vHDIQKr5Z7IuJ+oamRUOep4fZIeQpOYakUYH8PZK0JgxBa6J9
iBJT+wb0qcvxx8Vs5EWlRsl1nATQfor54nGaBTkY4fMI+BRXvX0IT1C2gQPc2gGa
ZktN19lXBlpP76aNw04XK5K9X12ROQ80OPJC1I1FXPMipiR/wLcL4BkUHKUMAqbo
Dw8jqM2OQar9Is/2IwNYokKM4vz45u1ep507NLGh0nsBXfTxQOvx/4SIYCf+wZNv
2SyS/SEcEvbyYBiUrH/OF0KDb0OK5eu3W05enu6bXlCN+i6vjDTfKY0FmiF0RuyX
a3PcYqgwUV0vc0ZbKpRm+Xaw7/4ygDCWwakVuVC1cIBZgxO1AcG/kzzPv+Ot+9fE
sPiEIjgDC8MYlusSenvb/Ns6Rdg5pgK/dnOfG+AILbYw9pB6ryq/PepYL+t5MCfc
dfx3LcZWSHx/gqpEWPtbCpYPVh/QnfAan6gnW4UBfiv2ELKTgLIX2f6oInUf8P9c
+JJrfEh/ppsxT0kzeEahAHSfIhrexI0GTs1QGWp0L8NVbMUiBXGVNRzzc6Jiloe9
DppuRPMdGTULVFVqalMVatkq9zcnp3anUI1JZO8H8nBXWJ4+VTctsC407NFVfXNX
I57dNMU1/fac92WP9LVEaWMOdv0WFvRKNzEIMoJAYJRFhAMSr9Z202easev57TQH
DDXkIF+1v4t4RTBsBOT8ha6Yrl1+9dR4cTYN4hbkCjDrVD6XkU/Hb1AANFaRfuhu
Hb5EkwGrebbGgMzVRPwoZcgnA+5eG2vAm1FS0/MAi9deJewCppdkTDxw2gaSrhUC
riwKf9Y9wlR/96DuY30+gJDeg+5KFEH7eX+BWk3IUxjfQw1gG1B7npyELogG2Flv
QGTPSaiqYIPDkCZBdwRS9CdcssPQwgY2iPjfhb/PJ7eeP3n1f83K7Q8BprnkhFc5
MdsQh8VUWyb6eHik+oQoyD16+lWXNSwN4Cud1/gfeNvgkiGD+rzfJ6x6knLaHdwQ
m3eYkHTSquN7coYvqg3CkbV5NhTK14kic49ilk6w/15UPdybcIwTbffok+I4UZhB
yvPTyG5RUutlbTclQv18RwwV9//cfp1+HgztEgbuiH7J6hcHCX/lQETkhzFq4LKc
HjfOcKlHYIAGLZ9/IeP2E5OgdB3sxuQva9ngAjIsJwkF40WghnqUzbadJ0G9cTXB
BVzplE3M6m7G5DFDkkhoJ7LxRRj6zEjSl0FGHvcUC+r8RgUazfJ1CYaCIhc79jFC
O3zOy/F5LO8LpXq2kvbrm+zf0tGykUwNY02Rn6SXxQxWP4wtIxYBFC/MkVWAZ6ab
jfWKSaBXm0qkAQjieJr+3ndY6RQclxqPmroH7rVsgnwRli8PoMCKWMg7k4+80g4y
WLU3svyQH0BKH3WFoQAe+zwmwYjsWDO+SGGIdPbe/xQ6KRRYmpAx0DbgEorHESl6
WRBkowZWNzeFWMgoKirbc8rtrYhQhssk28shmBxyBG8oBufkPWdzKjfiKyJa5AS1
HoVLow93LrLeP6HRgd6+5YW0WfKmnmXQVuh8vQMlSARHo97EewRAKqdFeWmnpRQw
2ntYjRM5SU2N5hoZ+vSBrc6MYD9mJlOJJv3CmJGJUtNPb+10AnzZ4/XejENrtfyD
2u6s7UraE8VqtC4p0Cki3KP08rW4FP79lPyOlzVWwL1+uic9iDjFcVeRtz1ZZbNa
j/+D9nLdtY4rcxJpeHzOA5zgodBKNqdAREb80renoevZFGZkAxa584RMzgTVC87+
chhKiuwa23TQOmqI9iVW7l1+8rAC4jbxEgaTXYcaI9rG8Mw8dol6DboqAzVdQPNf
NhjfnoerV207Hx3NURxXM7xZNgzusSKp66O6ZEF5sQDEU9Zn9nKiiGuja/envxSv
ub+dJ1xE+fU/BPwOtU3kAte3vvsENutQuYvAerDgVu1Siv+CBrvMLMCnAkBxwvrw
HqcwzdrbPPIQC8KUVg61H7rAvJAkTif3u6VfyBc3IQFBNzDkENZGOW8BAEIr1IZb
1ElZ7PJcoGyw//eGdTeLOq+3jGY4EMm7ZcXZNVodibpv+nwApiEQT9EYSxJR37YC
UC9cb5aiiUCTZaotkMkMgbccC7a3ry0Yt8hf1VQ+dyOfw9ABHzVHXeB3rykqGYAT
lWhB5dOcwQgmDu0p0XY9S7zrBqazkAySTy3IajH8Hp/hLgvkC6VIoFjiqgpbpHIz
rN3FqbkgXw9avkUL6/XC13PC/B0eyHBE6AZDPNN9j+CTfikmnhZvjzQOj1iJybrK
EFzkjzar3p2NF56zIUQEI9+utJwQ7mV9xRTb2XpDm6d8THoDCT+QOHwVY2+KbikG
Mzr/HtDO6c3Lhm7O39vxyQeFSDhfSFroOqzgqeuBFdg7puiKfmngHyZNGnC6rNNl
GsCuvP/+Q2TXra93vi8dfCUFZlYt7D5UGsu78EZERaliHzMl5ol+8lDJpeUIzLtR
jjokTUvpbdgxZaRiFYEHN1+LM9qqX4m97S959ssrAqysFBTvbhQP7mAGZS93TMdI
QdwMjEs4z5DG4c2mkYjIQreD07aeh5dz08Nor78FpvmC+S2LOhSxAZCcwMaS+lPl
WhjA3HIvt6NBHZ2zx6YlI3hxVfrZwojJ/glMFtvfAB3qWvxoq8jeGRtGNVFd8HY1
6IO4XanV7KWOyDz3UZDRp9NlkfNRJP9NsJHUSb9jwaC0Wqqhq8p+ebc1Sd/N5Hcb
pbH9DZm6ojJDZp5kRBjPfPtL0x9nzs/GfICxJ9SbWg1lkZwEVT5awtL28K/2acLt
OIa3qoE/OjlQcPVH1KTATdoIfKAnnwMWwWaCwz1AVVPywPJ/YR6XQt7Kl1PMHWoc
tRRDGpVJ5qweJJ3pONWWe7HhHcuVosws/okKxXvW6ZNwjL8Oi3RgFsb0RjZzvf/1
kssiapWLoDvw20+V1bSUiNvIcV4O7iYNTzIt5LMznnptkooM5sTmgcgK+3+0tpjS
yXxyPQiaXONuUNVRQb/fYuffx3MQeUHukfcOf3y0w7Sc70etqO+SghtdSE8vdnFV
9t2QeNv9csbThmhNfPfxuH56mRT9xnYE1GLe43MLD6P8SckgNwT/4NL6aA3LUrqe
85RpnmPfH2yBciniUnA8aqKY97NAMmhziSdVaVT2ww6aZBbu2VF0Fnos8kbhmA1l
FnmynDEJSR3O29mGj+OeVDaiYudEa3nUiLVDkdJscER45LZkAwpM+3Yl8piwvqgx
TMIAmmqO4kPIBypt6xvIHGDmDQMlUz4SLiOgh5GOj3M00/VaHZJaG63dp0qu/Tkc
PFxd3Ea3L8NSvkiRfgUZ7jL7hfwDElwarR87BanQLLG6rE++q5j/kp/ZWclNald8
sfd1gxpWzmOA+o/2Zu++kM2Z/IMsxScMf0ng+YEwQBkKju9Onf58keYqF6xo5BLu
HQdzbbGe6o7FIQqlK/boT2FVafwj56TnI1zhtwCvFFTgEn9xi0BpMps0TDwVCYnt
llWB5PuDBj4rFXrh3aXSD2nUhYrBc+TzJRvuNTgIVjl0XVa0RVP7LQX2J3YtSYBh
GaUjuMa7R4NBmoChXcCjekLMHfCC+KEn6Wtjf2qUdYGmtQwKIkXyDEnRbguWjaXq
iA2RJR+WE+yvGTf6dLQUQwG0G+TEu4LUcCgUzjH/fFVaohdGU4rkMP9nURaZVjOS
juf2n7rzDCmI1uq6id0Pv2/VZYWjfne6YOS9kAmR5PqR/PqYWlHpYsRAxkwG9Fwu
SpsXfnl0ZjYLwIs40Qn8idtIUVl3srhsYOZa7zyyuDDa4yOAdgX/1dteiZhVxc4K
V9Ve15Hf8TunKIIJ1uHbxjBDf37l+puZM5n6LxvL7O3MajKbCv4lQS+81q2aoTXE
FXWMd6W2ALnZwEHMLhj04ta1WU7JEEX32gzwGw5GDeSSBLDyXY4Y786kUVqMhW+m
EPPo/0tp0Shvkdkw3ZfT4o3vQIy13kimh1K0npMJqfNDnqpksaObxhuU+zT43juU
zc3y526XK/bcds8tHDcQ8ltkZU1eOzHob3lHzONbpDKVqPUsgk/KTBeLWsbinLvF
KTvO1Y2ODKUHtyq2iM9RPPcnxkW3gQRHfh8gUnjJMHRqqvw7MdziQHnkChc/A6ZB
h9fOLAidYZX+k1PGNXfZGfwvVoa46tvzNoYTkeQzAhLxBYIxbJp4yxZVeMZ23SyH
TCgfNCgOQH1/YQUS84J+WjgnqAbpmFTl5OUzLNeT5FOKev2dprHwyyjVpCMluH5m
CIIcicNzdXfM43kjClJm8JrtMocqFtSBwpaWd/ae9caPG3l8Bp03i1UEDQ7pWn6v
Jl4HPwbAlUj4WKdDl+iPYjd9YLwMEqUeS+cZesr+tpScU8VwQZgraS54evaY53TM
kNP4lUJmsqSfRpO4g2VPQ1qnWBnASIitcAjWo26Wvjeu43fzUJFXnm9Vk3PIDMOA
kvWeCXTj7p5UYKydsyiUri11zOl3IbQ9rOjlSVzoCdogfIvS1x+UJS8qA4sJoTom
S4pKPLT+mRitFkHD251cbnl64OcBxhiiJskeh+bEklhnpxpVpIoXgSflNMhO/zMd
odl/VeclCmf4ZfI4M+Y4H6xFwf1KLprYSTZt94gH005dqP6qDzim5dacKkzBnpK0
uY6GYD726s3OqHquuzXC+RNnlDjJZqCYU5MSLgwD1R4D0M3yS53EyjZlmX0swr5j
6QD2KSgTFsqp8EXI1vioV05VoCmgOkazzrwURW95UUA6HIJX7JF7/KlnnG+Xap+Q
F5Q8mBHLmfQZ15cZ8ZE5fsWbmN97Pz7u361GLL0rndF+7H55NjZpy2xp0osWsN5W
HkXXUMq0KDn5J2UEouejEnvb5wAKv/RwUT0KVfez0FnL0E+ejD2F+10iIL/umu0j
rWoy7FYO7pmZmHfturrevSYuyYM4iCrGrWmBcPPZNeMYwER3op+RXZN4f89haoAl
7wVeZjauNQiVWCb8wT0WqRPRInku2UFJpBBe18z/3ZeyHcBbyAbLeMH+D7yKUjVA
Gq4ezOQ8ejrJ87RH0NmPTacMdOfmGkr3IY87zdzwe80EmNmagkxuyyXmGkjiEx3X
EYfk88j4OoTewGF8bjihubRKRWahKJMoua3hlgiEvUr1iuoYtM2jt1qrYY8Gux2d
6ceQOev1DqdNLoldFZKL9inaX3GAdwOHn9JD9eChO2+cH5YYHSOAkNR441FASiUT
fjMpWKR0aZQnz9ghYK2dUZeAoKjyoEOUFK4xiQUpXne90NqiQf7KXl9o2XRWWcPh
X2/xvOAg4SW9HneXz2GEAe/NsybPL5ZJnedmdRUf3Al0QJuvKqr0J0owafxHe3fx
7TQn81KRkUemPAaCXZ8UVD8KWgT/jkuoglR/vQX/m5oYpQZ8H/H9QuZ5LbCiMMBb
MCjKPxg+nW39LEtJ37ZT4BF7bLh1AFRw0Gbw7XtBHkM4aGx6Vj1YKdWUWblIC0CC
57nSQItC1zIw+DiZcIVPEx+bW7/UgpKZ4sLRXXuGj/46KBxLVDuy+nZRgq0lwhdv
tE6v6NpMx9T14U+jRvpj8BtMuwuemOu/uYFVUr97YBu8+8AWFmvMsFWTDmJmJ7ko
6TRxCyJOTdasVk+H8xCBkNoz/SW8SGmA7t9oNH/XTJOFb1Er8v7I9JHt1dRHZ0Gj
UMAofAUHhfDy4awLdLpkszANoQMPh4a8bzp9zEM7DgNOpT1dB/z0iLaQdyfyI98g
HGoqTVkuuobrgr6rImWPnsJL8Mp3VT1cEcCfvtx1yys5jFJgqqRIOYtdmzHzoY5V
/tR1xlEUB5Gm/yn0Nb7+4dXNHX5cJg2Pc+dfS9UaeiU3XYTkcN/+If+K2OglSTGD
uOzb5vWSIoK36pexgavRyQkG71VojKl7qcTlvVPzigJHYjZ2ubqEbe8uknlaaSBj
QVxuTJ40QJMq8KgmU6oPrIikDUXjrbNGAbKUfcudGCMe/TTnfN3Whyg5libDkAC+
Xv8Vf5CTenyCbXw7oUhAffsmkofKKI7iSwe+6nLBW1hWkEHqavXYDrC3ug7BMW2R
rA6mGcPpZ9L2dr0pSkhB3q4/N7BEPnjhREUU2j2ho/fbfzViS8VGOJZoqE+sfmya
Xc8uIOGsygVOYAYX0md4vtDqE/+tFJ0f0DlpJsd2DAveznVi35A7qbnTEcMiFDud
ok7EhRbD7bI0iv3FE9YVgd2KeRd3RTWFLW760g2V6YgrgSw0iMzlEG1rRQye2U0v
aV1+k8P8D6h00IgXDFHGY0CbQvS80vqNXdboBx3n+i9FtBjOjS+NivhXqrvSk9U6
2RGYMaNR/rybjQNX4kIubYHMvDnZ/RWSiqpAcJBoI5EUepTj0CCJ/+Nahx/WK27t
xrC+Mf7TTw8X65Zn5MvWoSN8Sb+9Wvw7xe81yzP0Ny2dGZQ/hwx+lX2zGW6P1jhD
Cl6ap2deQyxOuMybMCAMjbtuI4eOw+jVNfuGfqOZPTdPwijOEaTIvTj/qWkFDsep
z8I/AhwRtsCnGlz4pi5KVX1QYPuKQ0/ElQGeeiRRPL7wRxGNFcddob5T2n1RQmx9
x9gx4j6ip5kGuVKxOGfEAfBH/lwu4h56HEtcpag4ybst7U2vO+Ab9EAM1XNk7InF
SxEsOcYWbS80hTfdhYOEKad3mXjJsM257cQwWpki9KmexE/e0ltTOspbwJ5uaWoN
jPwvNJVfrtVKtE9rg/WIhymJHeYJdySE8amFMrjiOZZdVG41vyNwnh/FEUkS4msU
P7iHGcp2oe7kgUWWSrE3lzJ6Gjn3x921j3x6qnhoh6fOJeqtSYOH/5h5RvMjWiBI
zIixrHQNRw6fDu9M6vmtyXIG+R3JC6YwvoTR+OtIKpUU8I47xQ2T6cYBfHAZj+nw
UCsOpIP7Kk5ugo2UBqMy1XEpPhSeHbPGFvyC5EdkyV17idySfjovPMZbIGSlyp1e
6+Jdwn9xYNLDMpPlKC8vJYQnsxbeRyskdBenZt4QVrQqSZbgz8O4qXBsEkzSxP1g
0la06NTvyk2UhbaIEUrIBWe7+zzAFt5+WqSlOw9cL8yhKIc+2osRCWEbpJMxtFJ3
aNrLADxzOB9h7OUdT/mYiM1/rYKk0WagMm14HZiqKtcKaNmj/bKVdYQ5BoM4y3Ur
oD2AyoxjxsZrB278fvn7QSQ+pSC2IiGdJYH5ZFW8empPrQ3wfrllSb/p7Y7LNKh7
obC74rsUhC0lrxmfomqbHUOvGdE61x+Z/+Mqk9O+MIXxTPVeTncYVM7GnWGNEYYt
OrCo8J4Z7NY7CkuZReistQ+2Nf5ThfewPwb9hMxuL/e+x2kGmTj3wffln8l8usjA
t+T2yAtgF/umrSrB1Ckv1f/9Q20UmggIkW5Cos8OAsIEfm3eVp+XVYsKaB+TRgvg
Dv/lkXpURZWr/dU7KN0jpnl/nh0aVp2gqvXZUHbZy57C/HUYYDn0I6dE1bm8gHv5
ITfnnGlJK3ZPbmbHVJ++LFd25LuSXPxfax38eCLv7qDns5/foiMn+h9M8GbgxW3Y
Vx7Zp9vsWJJO4G3wl2b2GwUQh46SAJROXdNlgx/69LzmxCrCXmYBpyN0ghBNRgtV
+/ZrRpwgaepr+c4o0pa+3QsCIP5YgODNiLoRiJnDSdZ1iOT5r8fmF/cuHPe10kEi
OVidjqIRH1NOzthejb9NctbgTJFZXX/j2c5GMBXUhAbtsh+5IeDf+zKyu4j2pi5q
0/iinEWpyBLSzKHaxpmanl2WOXfJYaSxsglIW+DvufpYmlC2sLu1ed4eXTNV+KVO
XvP7KPXX+ixVaPK7jgG8iu4sByBe3VKEGPWYTAD/Kup3/P6DURZIVJqJXkXtKcbX
/Qvg0leHv2YyYs+iu0k02UYsUbOxmKP3US0kr6emfZPAJvHJeiSYrkeQ3BzllZV9
Zt78ZkfraZfZLDpej/onbfUhyT5pDSW2exjCiReLMlaNC3/1OEsgjTDgOIoQhqil
2TjMg542gXcmpeIW4tll8pmHBqDL2lZpKjKjk8dXuG0NoSub3R/B0lYWn0bQ1Q31
ii9AJqjoEdNPX+kDun+PeN33529LpXFJrlhmMG00xxu0zjrWaYMw15nRnyCRD47B
Ht0pNmou0ccVv05h33+4IKFlrWlToiqZip0I9QkjID92Zg+IhXKdrWzPcuRZt24r
qFRWN3tX1D6QrONF36FpODt3FMoisLgVCuhzfMgswOGd3gU3rxjGZcHsLaL0bOu+
AtjFdvvB4N5uKvahsXvhYNljNMBpiWw5X04Yb4JyyvRitjvkHh7Rlg5LZXLdOQAP
vwPAyXBgkhXHOTKchJ6cIRIGrjtGRQ50kDm8uhebvO+fd0OYgyhOZa1amy3uayhw
bLHXW0I9zxQr10Zbz4nK8QtE6gRG8NtPBESNDAheZxVNDIzTOMaE0RrS9X8q5w88
vew9CDIFMmjP5l1PIV/ZMgWnnCkh/7Fkfvd+CXDx34ENiaTCeCxcJNojqq1B4MA9
H9mpG1lYgGiv0uiucHJqK11nhalbwu7CyhZOHZNbwGDmIKhNwI0HqFzdkWpJrGPD
ODcNqVO7u+yq3wZbA5+92kF1ZUiCI8WtPGRwwiP7/z4f2GHIPLmqBpkwvU8W/fX3
GKiB7F1qpcnSxs8PMx/DTZRlLr8gS0HV7opn4vaUNI9mXhNIXnvEARHYVuBYVsPu
lsAaqShzonFarWTcR6dO5yoo7xxzzkt+qLx20WrrH1RK4+4fy/UvUMQV0tNie3XN
/A0iaaFmhctowwh0+u+STl8nEidw9RFkmKMAOwrs9Ds2g7V0ZwsPTwUJvZlcN8Zg
VEyUl0obW2U3URHeCZ8KAVeQrbzlT1jDS3gM82zyOaNscu4ELYMhJaIn7OPsqQpH
+ubCS2n5b/dju6cCanH4Y0WgYqCufp3iZ6TrXq8j49gjBh5XG5yUgeGYfy3WnDMj
AichrZZtwzzEquVIch8fZP+S8Ghsb2qtsG8N5a/Ax1i0A5Gys7XkAj/qB7O1hnhe
Z31ooeXd5RzIa5M1DwEqMmgm0ZzyMlQ44S455JwDl8UEuF7CChtJ2APOBq6Qkgci
4OC92vXbvtovzcSna/UAoJCfR3E4/z+j9NcUkhqK2YiqaFRb9J2LHC50nMFv8Nz6
0opVVH+Bx1a/N64D8nDxjUCAQD6dkukMkQI/U4zcAtBMfWsT6/W3O6/JS1el70+D
dh6JgYUGSvyAiiVLmQNgVWW48DJ2VZz5simOE7uN+PrQZSXEfCBfjgUoVeCsMkw6
jhY+eF//gWbv9ArbPoxkm+ncVVNlw+6+mv2QmMuqUjHdkmWimDir6KLYbIN4MYRf
Q1PSnHTr7iUl5PPGwlfT4uFAp2IwN8up8f1FSy0ilxhc8sFDKFRji0tAVGWPpDg7
OfUYygI5MjgnrwkTEOSEE/UXynBcR1nkWr3U08hv36sMKXkLQHBhrXlh+/C881t7
KHVwZThqSCnoncS28T08+q/SwEFTCKGVnjWJmPANnWrk9X5WRAhHdaC8pFUCuMAC
LJ6Vh/f8sJOf9VrZTDxmiRNy0WW14eUw52lfMAJr1c/++PTwqmm9rOfN4EEjkqRk
cokIcMaA4dC0yIV99ZrUrroVTwZzCesxBjU7ZvgDLQavoFR2xX+NqsUSpiHvux2b
Rme+rj3/K+q1j3FeVYevSAnt0ea0YKsm4QACGWiXgvAh7S4kCrIcrflzxZs8VY2N
NFICXH/5hI0TmEsJwq5roSKJ03IhMoMsR3vDrZVgwMenobnZrTHefOg6zz97G68Q
7Z7frs281sdTrHR4kikdO9mKLCvSAeoo0wiA72KI8gt1uagPTOZArte24E2Y2U0Z
96SZSd6ScorefWxTlkD9LSr1oC+NhfpNUU81o240l9ptdVZF67FJM8LlErrKXPfY
sms1Qomo+AcE/g1lx8leLm5vHLzqWif2IQif3/FzdHX+AUyKqYCjZ70Ud3Bo/GKQ
Rox4G90sROAvgOwcJAwYegUV4tNV6DNIoXCNCGyNsp2k/v7A4mRgXhwF7TzEmvOB
1ZaSKKi5q9gnG4TIqK3dqrZeOfWRdsc/Cenv8RFiIDnP3bzZz3de8+HvjirGraT5
eeBp/HFTPq+PZmDHkhM6winud/v3TYXn5s8uVXMUxk+Q4SdLgv+qzmnAuvrA06TO
wk7IOj339ZwmZvZuQuHmFCibqpacKxlE9LsVn330RIRW3TtbQl6TTrpoQArhjivL
XRpf8yAWJGr4qyqpfLU9QzFbwSiTqQ+b76g8/MCY/1a4e3yJ/jmxp0HY51C6hJnK
m7sahd+DXgehLPayFqUBVOdBRAmYpNs2V6yrptoO1K5MvLgJXYj/0BtzL9LbhtMr
8WtwzXDf6X0QjSzDLGV+CJyVFct9vQuOeiHS21aZvRywCxocOv5dh0mbox/Ah+rU
DckXIkvhSbQTP0+cNRmu9y47614lXKQiwJVSKGL+f3wJg68dC7DcqR0Td120T5k5
WlHyDGe5QItxREfWdCAcYihuK1JBOodiO09JSRFhVwCu55rMPykG72eoXLNx9HfG
HaZDDLvuwh5G9n2D7b1JCpcrp0ImGKZW8AYmAeU4v7e4XGSc1CnWYVnmi6VbqhSi
ZWigbqgvV1iMyz9TwvFS478pWksK5KBjn/9oimDq+A1DFZtM2gMynMot3Z/wxcwx
5C7tQ047eYIYxxettWGmSwHcmTsJ5GW+DdO3fr1JceYuOm6C10GkF7r6Awxm5L7N
m/gskdtItjoFUBnH/rfVNI1TMrZii6XfAEU0frwEXArrSsvlPM3NlabuPlO6NFaA
mz3um+i1QnRXc67LyJnf9Ea3Jw3xCEC0XCgSaZvbtfVvgshH9RhpA0fXyr+Ql0re
706qIbhzRn5z+JanzN6wCx5N+0xbCdxP4KoEzPPl6PTNnlrdj9W4doGJV0d/gdC9
nZJa+agEYmfvW1FxD1Cfegb6YA6miW+KbmtKFWM+2usUvCsbEdgsPA1+2InyqK8R
PUyEfJK11PEcNLWsqzD4acOIw3iGksBhU5QpSQ6zKSQdzZG6kKtTRGcD8s2QvxOV
cJhCbTiEbrgy15+MJRgZyZoUe0PCi/vTG64RCt9Fb3a6MDyT6u5Cwb+rnXBSfhYF
ODZt82jJFLdQPM0dkLQxXOhQexKXbTid71+Y8sIHzioyoism2WxZVpnYpUwbEgoX
hoKuUfsWrcKF9tmToAw3mWfLB1rk1nxxwN8jgIN/3vXTvqaXeRSEcOJiaax0btjH
elI8+zOkKFGzn3DVkthK2u0esG/6PWSs7zu2DNQAebMPw5hE/un2DMd+Ocfhn8MF
xrAwwkdzguT/brGj+LmHw9THfrrslbsKT024fRG8w9919v/REfeEcmQJjCy6A2xj
QecruYrJNPb0C/HX8dyqckXLLc8S3zjBttCpaL2MhySckXVYvnMFzzwbKIurKCj0
lJEAsnIHCEP0XnsvAps+MHlCKqLlLfkDVU4y7y8Qle80ia/PstR6xf/R1f+LRlAJ
y7wR56hTx8tPCSv7/D+wRjRdDowdAjmzDqunu3t3BhdjheLdCIWzF0ljue+HEFSQ
3q+kLS1Nz4ajybP1wdIegKrWH/u5qi2tADLj5yQ6Vwp4m/LuAFvrw19+GPd0A9gX
Ib555SU5CaZr0ufvDr64hUE2i+V48Oj6S/RhVRaPEU7LwRDcnO03vaiq7Yok8/U4
jGhNMKLOGHdttRaKOzl/XLC/M8st7yaGfRQqGr23acGTt/Y4eTemzHzFfxauAd0H
7RkbNuK60IIhp0NbE7qV3QQeFsQ4WcNDt+GvRMZA+oVaoDpI7NUykYVlxl2RGvNi
ptkI6YXUfhJ1opsz6dTCHmaNzDE5y+4RTk3ooSZVCCKPIjdiJWbx1euiaLxUI0R0
VZiL9A52PzXGauxgKDnbbbxTiabcDxJO/l4EvWNA8q/+F+yBF5+K7YnuWcFCGG+w
baiT9paZnvilouBAVDX+jKblmahfLXfqF/kqzlXry31GNIa9gIf1L1WaY1F7PeWj
b3FfvccrPuxXC0mOpZwHfzDsYX6wU9mbUMhl6awnNd3DectRX477OCQZXJ9+fyYM
F0EdgJKwYtRPCH2YAtX2J5bMHgru0DGmB+6G6YbWxOw7ZgR6iSmrZ5N0lb8YszyP
3mgAEBqDyTY2dFfOlcrXjvUAOQwoYIiQ4UDnTZUhKscwO+UnEzY902N6QErTDu1U
Kn1Mzo8tHV7IbQExGnLnsIuYLoZMSJOeEWSMzAlpWjELux+QJ7GMa5+cqCkQIF5F
QOJ7j2Mo+kBgyjhZ33oz3IjvRSCtUzD2RCBUislDpZPtCdVDNxfFhoftogS1gW8L
FlVeKucA9HhhKOm/spK6vi6O2ERM1zBmscoy51KzLVmFmoRdVJUkgXouBT6YBIp4
RORLRUAoJaei5S5jtBKXSsIsQDGNDlHr8aPRligpB/Ici+uCZ85Wsh0N2diSaJLU
Wv1SiFm47e2ldz7rUPapyxcEElIWE9JDNJPLlg5Qn5f45zEuJzR/1hy1sSaP9BzH
aaYnc/nE586XBQzglE/vUnkfgYdOzUiJkfs/6+xUOndZHcyTPVHhlyUuxFC0jrNJ
m1s7iNLB7Uf8wHkot8l40+R9BIGFW7gAtB2D4I9CRpiSh0txHujjg85hQGZf86It
shZrvSyIR7EtWjuGc2+UFl8RBnfHrXcGLlLWxRTF7cupyJwFlxumMoDdeQzS46rM
n0VFrb5xN1IEZF9MXAnlX38D6jcYZCj2iQqeY1Ot3lOUy2fQ3hsJnAuvWYlyF4Gf
U3VjMobIjQ5N6qjg9g5o+nDgl6+t19WJBpvWOfOSby+gvq3ST4moP2xtLSKKV4B4
NAI/B2ejUpGxx9C37/dq4sGzLfwrEllhy5h2gw6qJc/4hbEW53oY5C8ga/ClmLKm
QrlNZHEIc24lCWFYEliy9Ln2mmfDWiZJxzNXEq3xOUzwEVUI7nc0BkS3mILuieIv
NGULTDURcEAkY9ymi/nqWsTSU0b3CydCHmu+MqBuvKuU96sqC3DPfdGymuw68dh2
sTqB2M1C/XkCQjczVMj1abonOI+YSiA8PNjDCEudQnR5KYGmnepssNHFSNI73gWB
6Rt0L8ExFKakGSxXa4tUPwgSU804LSheW6iiKhGWTa62yBkeEpJp951E4c4gBrsr
jmPG3Olb6NiTksy0MZxfQR2X5Exs0/EKP8We824WKJ5MLYfPlKyLJTGAQ+eriCCK
kZ2gBeryMeP1QaVw0MnXv4A2Uury6mxHXSRNs7xWGWQ6oaB2B6RQvefUboVyPYaX
GSkW25DNA/87Z2XoSK3XewmabPZkiKl6rn2FajWdlSyhIkpIdOukw2VOmBgI6TFi
M0MV41qi82joELPZyp5VuMzt3fu4arZF16AzoD8NiCNWYluXoEZm3nn9RNXieZGv
RcF9sl5GzWKyeXdqs6lO2tJKSwKHls8Dv2/nVX/gys+R410iXAP470wHCT+voQEt
+HEq4VNR9LDGotmuucvkOIeL9S1m6NDAEfMSbpaCWc8vHhtc9vl8HODbvWBO6H+b
t2Jxi150m7O+2s6Yv9v2wdGrQfrvp1BZjFDghg1E9q6Os2Mlma+H72t+9pyFE9vw
5cPBlNvoFYSBHI6XSgFO9cU+BejtmGnE5m/rtWKJaevhK46BmTApdiouxTyHQlfX
0ZvGXQ8/elh5zjhOHOj5FoE4mPSxuX5GrrC1v8ySx9IBIMfFiiiySw//vjsXG9aG
gesKxrCsUtaHD/eahYhXSoAQMdSliN3FjZRvHFbI88kKDQ2lu5mPyfAqxL+QkvTr
Sj4JEynDYa+RCHKs0YrFetZQONHqBccpfqzMFY/ZEhnQf9VHFzJLfIJnZsJPtkaR
/5oo+lJFczdqPoaawH6ymAc7GnXjXCWvYSfx6W45YBI0VmZ7ptzv2OLr54unPnAN
XJSS10756/uH59vb35VPhr6hbAW/WAj2H3t4suBLKpuyYR2NxqkoLLf2NoO7ytwM
OOpyhstmOCKTJtByhCMLxgHtCEXzPJt3jRu/hjYH/w0b717LLxHBaIKoR8j15YZl
1S7A+lGW1xswTMhDjxwTsmwg1EOHxWfLp0TQ3XizD/AqK4sfNnkWlvnYs//WaKIx
h60qQkTtIdlvqjUp98czkuXxx83HwdrVXwhya07qVaFIoaHHGOKEI+eX6zLbA4sc
RJfqEc+sFbhj2SKCfbgLqwJhq7rpzD5UHWzB150ytHUJg+Pk4Fm1erhndVP0GvV2
vJZwAuq8/5P36uDDjvH6+Skc+TNnG00nOTV+PB3jFekXZvt3bpy6wRuJtlGoS41C
A9BagZ+/gwhjS2bg3TPnSg95qbGR0THl3z2EbXfKOTFxvDNkfvtC/e/bLSIukF1j
XfIjrh+IoJOXGpZRP+0WY5RzqZ2PauR+BYTyNNpZZX/8jlShCCiy2HxIBGvNuZf0
Nu2TCESs/EB/9KPXJsUsS/McowXnr2Jxdbco8ZjeAwk1nS9kgzL8ynQw+ppnI1B7
GSqVtaybvnFHPGw3JzQ8d49jjPs9iLqpFDHUm+h6nF8tAo/h9MxaJxxwp6auQ+0r
v/HfGHb7m/UOQ51EWuF2fZ8ohGag0p6KjDGGcWTmyz3F/b0Wr1J+Fr/6Utd+Xc3k
Og166uPQxcNY/eY+CmYO4HDrMpTSpGXnAEh/7A6ypMqSYL7jonmbAEsYqhh11klp
KmHLt2J4vaFIOwJZdLkaBFbtJxBTXt+wdsOvde/mM49CSNfHUKOKdDe++L4TMIhe
lc2ilPJ3ksxt2QD41D0VqmeGDj158eQ4lSZpODLXxZiCJuAVtoi1kwv0CZ/UmObv
zY2dN4YNMvJ4ELChV1sRpQ0W05u7WHDNtTzK67XuCP4MuxOtGi351JEVzVTpEWro
Gl/XRPG2vlPOEuEsNesd4BOU6HZ1JCHw+vBUbTz1ubowYYaNZ6n0ocZ0Sp8K5+5l
EMLW6+CrY05Ibaz4cm2O5QKPJs2pyyqAyBf0zIgkkk84V4FPL+G4/lAbZTVjcNRq
4Fowo0IV4LFP4t8YXrcw3sN9q+FLtqOrD+Ij3sixBU0UAGWdtPAthV3Wo7+a6D+2
gKYn+n9FGVkxBkxoB1jfpvuQR1+14l5OcpfGutcRn5eSjok+iQj5MCS5PvzLcIUN
DXjwCDUaBH9epHc/yT5RN2iMQkWBKERo3kRGgyEoJtiJusdzLGzyDEYX4fT5kBzi
K2HJyj68/N8+CsIRABvSBkGKg5XjsA8N4kmC+sLV7aRgXiTKS3Xt56BzGQS+T/JX
a9Hg4LUDgygbG7qfZfmJdj9hNJECwundmGW0GSiom89xbhC7C74th2YUE4gSyzhP
9XetGB1OVcNNnpfVkPEu7aKb44KA6wLULhVZTLHNuJ3sQA8kPu80QdKU6iagimeo
tBTdVtXegJ+0VcwuJ3ekIPnr5/TC1FW+E45flI51wtyumEdgZFGZlWvok0dEwDGO
sWpEBFOuWrRLVEL/oeqU/b2G3E2G20D+PZr+QxVw9uVwhIu8eyiwsx/+FxYSxTyO
1Ll20mxyO/dmzqOksZK23qlF59OJ6yF++Dbr4/nQxGYCPE53ifqjiBUkeOsusalb
LfbhXmh6ST1u/JNnvRUtlhUBZI1bjXlngJzju2ROQqY4HRC94EBwVDfFIKfUeOtT
UNw8J2+4lSVTQIvBCBFlN0bwcsn1GnkjCg/RzSFI1dZFAWzs4QOKn8ZqfGZj+j/E
xXCH38hN6N3fFGREjYUg+CuihVH0f1PGAEhOF7xC6PJwtxy2sg969kB0i5C8xz3y
aF0UTBVgTGGQWckBdxoOiJjqPwTy2sypUKd7h7rffLV2DGVxMnfKHLv5xgJzpJkW
pH+Pd405gBE9LkPHxr+GL5e6d3lqCWWzlI5tl/A123/XkFB5giwVTUJE3lnkfO8q
Hva+T5fqPO4hNx67e+cFZKYvjVrideFoWRswk6aldpGKjG9y5gPboHlt8kWG9Eiw
4rPf+FEY95636qxdIj42e3SNu0Iyyx0YEy5cjeEtIz2f0aBO2QilGdPoW/xvzidi
0zw+0KWDHzYWvssEjaXkfcQfdlur9upzUGsU74lnBbRySHOxkKSOAEskRirF1rHz
ZJSbTvDT3JHq5AhJ/UXS5lqO4nE9frPnVEN/lOa5uBlYV7JIbzRYYAM/Z4BxdABq
rlTNa4II74JqC8HHjOBHb46tMpgOILzaXdOJxtw+Ww/YQZK74WpMtYOCIJnFbLD3
xfvzOU5SrYorc9P2nQnBYGMc2bmRUl9dAMiQV8E3peeu/rJIBFQRp3HnqY2lpIf1
xf/qVje4wegPZLigL8KM3dhMBcyju0B5yqT/GGOKwQFhMenBfcjU6mwzKMq4EyXa
pC+UFgIJJkbam3E7bPqFDuXtlCSO6+dI3ymh3WH4RMJNRQFtm6DaRrO7RJ6+3g8Y
gb71IShhV1dAZo3wm9DIeQhD19fx6PbP2EwfEHsdC2sFCOLtzmq7m+PmDBRLTAxA
kDeRd868HBRzaqQYp4Hf0m3n3TeZkvOMfs0QWKPoOjS/PK5O0Wl6yhSpAV1q4cnQ
HTENBVmRRAJYYdrwBzWFPc1GczpqsAzG5bMmCJXiHbKmYECxCCde7u/FT1dADBCe
nKcPOp9E0lvqUe3P0dFUQSur4lxMZ4Vc8/1GKyIzIzxZHK8OWXNMhw8fFe8NLimT
hqnNFAmD/t6lri02/eUvd0KjN8pMB9rbpVjYicD+xpRonA9e/QplhRnf1L0B4ZjA
dAyfZ1xt3UjjX3pTbd2FQo1v/ZT4jjyWhbkcAY29dwAywe0mgac485yu9Aoqc+dr
fU3WwNS7Lg/xLl8Df+z8jFO1YXiiS1UZ8OdLuOYo4w8s2XvrTQog/zPUQx5SY+GW
eRQXqgUmWiaxaG0lVTtpwtwIQNjDHQQlnI6cxgaIZAeGypYriNJ5ixzcKun0AjKB
6Bh1A9Aho85vrx3sot4tuoxFD/a8FwVfgI8VS5/pa7cAff7a6CE1r7CMyNUIgXu4
6GGjPWLn3frdhwAxFbiPvBFPzPc3Nnde5j+qqPj2V/+l5+/LhwocSNnN4wZC71NS
XzbgwINPjSgjaFiLT1+V64Jz4OT5/kQh85S5nPDRnIMWlUOCdvyWeS3gKG8CtU6V
HsD7THUCAtJnzJCL+ec8keEJnvXPYe/qd+/DCTleiBaMtvdWrAHg7/AyY5jnns3n
N694tyCcrY9Z1qdOr0TdOEmFdOciGa1k+Bh5Ks3D4rkxtA7hhQ8jfm9CN0QtyyKI
JXfT2x7f/UWeTxptoJyRafmxEa9+ijbgWpALQRXyc3Voj8EoJhlMKypwcfykImAg
91nLlvSCv4YJSHjVGNg1iAxufOeVl7tEnLZAV4mqTWc/AeVGNUQ917Ic9WLrac/q
6tR/O6ldSDXShUB452pRI2eFb80KQPB72x9GtqeUIXk4jxaMo6psZ9oGhOu8i1NP
5Ibw77QVzpgx5LeNsOAEvMh696oNCnMgqVcektZKyOPW3xE4IZJmtP8eqbL4PtOR
Q9j6hfBR9JGRI7kuTNGmoY58ahCyZweiZgyebeMWxRJ+vWV0Emvq7sKMij3JB82j
dGkU52hEljotnM468VZIS7PJoyl/4sM1ya3OKTAUIAlwNpxdR4lC8GuGkp/e7OxZ
JvYJAqayeG2gXZrFOs4rE9rJGUeT7H8bg5ZR/lGIzOQn9JS0Guxax1lKTxjVS5ZJ
42ow70VZlYz4Cqbisn+i1gtuyV4hu0mKM9IOYXNNBZ6cKrV7Cy6biRy9S09Eswuh
D25EXs0MJcV3x9PE+Ewd0B9Qh3QjxQbQ7rGMVwsbrf4Epccsr734wCM4cdbt1w6O
sKfF9pgR65/7eq+3AF+0fSu4btz0p2TDdpiRc/ejep0AIYGzE1tC5MIYuAllXBCK
8JxKx11I1INQJAnY1KBgAtIBm9Tpj8+wWTMBCVu3djG8UNbH2+hU7Z7jfeBYHdWC
aR5iyp9TeOaoX5nqgpGaMOSDNSj0hNbhTuFtBti72Wll24Qt6EUYRUdO9NvhfxK7
d6Qq/zXgsxIKxziqh96rsiyL3lFSyE77ctR/HYdzXeqSrNfDdHUcsxM0EesVX2wi
wEgQz5rMfC0mtMtHAb7mLq55rKRoeBhljAWjvCbE7YZGKSwHD3nB+0pP69pdfwrE
OQPuUcndrw59puZ8kyPalr/g1c3MBBOOz7xFvKI1e3xzmHYn5LuVYwEUU/rLiHNj
xXDcZr1kJiDE31OCwtWNKbCV/1uLoTfIlUqON0s36/B2eoSnSG9uQ3J4GsKduSc3
gEHojmeSHa+jy0vWSOan4oipF7LvzRVkaLBRCuoR4SfuHkVt2ky1AUB0k7MBvGZt
f5ISIYWYrDxN8GfMqNTs4GBsynOG628ol/6M9dWMYGvZl6BPKTXTJ03DkftMiJ8/
vqAyUcMmDPQynMuCS/weQts936N0o+tO81Gt2a1s5cc2tNNXW2t/f51CNfsMyf+w
ZkdyT298pjyHrVRQsxpQt8oMkFMm0zZ9FUSPc9i4Kexzt+rM7i9Wh4D1uztT5DOX
mDjjVzmOEiFhP/PzzfGSLJOX29spha8WIkPe7sJZMEWDMjQn2lxVQrjz6JlmK6gX
fkmsXvVEswS21/TpcEk9HFaw8zVGDlhcP6UaXBZTjKc6jZB5UQtL1bxi1n4KKsBf
CDdlno56Op+7MEI+ND+fuyIuFQqF9wY+LTfIEiV0kUahvZFnt6g5YWSoc5y14lPw
W/SHY09DDptQa+R9+GQgmFDOErGEB3zqEJVqr0NsLz3gWjGV4Wp7iw9Tqib/42sa
3RF94okX52uWcuQFSKZXZExaGWTlIvZkNNQws599eQcgIp3vYkz9PkPa6rTRuHqe
/V01km1MD0jOlqWQ/BhckVwxjAIJg3hF3U264IT/Smvcx0ZO7DVGa89Q3OaAA2zF
15b55yzZYk+o8rhmcpVfuPaRkZbxskIzVocI+rwTzLz69xqEMHEbPQG+6v9kcN9J
hJOiTd/zah7knP9NQ+u0/lX03jqH7v8+YjvKsZ0eB1CWoQnfcZvG/ZsI4Uu0GwHZ
Shfms1XbG2y73GlDfDNfrkvcgeXI2krNauXjHURIbxRbM8Ia6mroKxsjBN79Lx0S
NnqTPCvNARtPPwxEDmlV883xZDYQjoVJ2/8M68e8EjVRjGfluHz8DqyAUG/ftM9N
Vf9yazjXDXuZ+NgPxsTbpc9wso9ew2HGdgX4TKIalSbPgNisrhWWScEzR/52ZTxx
92sfZtc2FYzkbQjlFM3O+12SJb9legpZfBKpQ6i8rn4qe64vPx4vy7Q9QIn/bXVt
hiovkyT7cWVRO8PleKbaTQ8n/ua4yx65xUdH2tyqSC59t4hy9ly1LXlKDHX440vH
QJwk1HkELiOg9Nnc7Cs3C9cz6HtA3568DVpniOn+fIx9uzYEc64qXKxgZnd3wnOl
GL7taiq+Mtz0xR1iNzmdcDrjvqBTBIbwysMOTVbSbOoUVgMuGZ/6HrtmPZYAdlkN
P1W6tYFp77gq62/J2ZYSWIEmtpIebR2ZFhqsmBOpOR3ejuAMm1kqdZ+mNgXEdezW
QnFT0Qy8VL/Llt/5rPGI6tp0WinQwC9I4vxc1dnnhxtKHAtiewn+qOUR/cIQFFZc
mrs41aSCVxwKS/PmiDRlSpJoepFzvakVCu1JLMoZAFUqkA9fEZw70Aeya71L8auf
YpptvgMlt4DdwPPwP9mVqoP9I9n3ujxnUC5tnOXVQHVzyN8XYzgsCLxyEvORcks0
spIw53xWouDIF1+1Ll/XSziP+bVz+EL9yv0fNi1Ay+AQ5wwHensUJxtFwsKr0Rit
5tXtgvBikQ0Ioq+21QeIcuhjaXw2WngTf5dUXYd/hzPYroJqPVm1sciZHM+w5GKF
BrjDgHVFUuSY3pgZ5CnHhCRO35IMzBc4nSO0PZ4uDziGkxy/YXUrgPxJKAs1s7u5
S2eKG9cvPMb81kx/aHiJsS81VtvhjKi11fMHrMJhdGU0rIiw/c7HZFF/y4RiWCVk
/DkmJeuggnFe6imeU9cygXMKEBv3wUwIMf2J3X1BT6ABmah3dJqlSIJidP5zMY6O
Dh/9pURLqj4yB2PyNgX1dGrlwJtxu4tPpYcau6coho1iZ/7uGFIuyEOHoPgvFQWI
QvJD1wWhITiobG0JoiAdES0SZsi/J8cVNbUC2n7tKoYoNsnMlB2UtC5BzW9UgNwD
u5zmgOCrcSPPaB65M9/dqMxXc8ntXQE3Xb37vXd0PGMQMW+7fkt/zEZvb306pZbr
+0ORLn9821qlb1s3o8V0gN7uOb+EViIbR8wiKQ48VDKWi5qiHQwd1TB0UBLj+dGl
2gEsxpHfdZKeNnGvNyRodiMqXeZSQzBU4MlwZYZLPkxSbjtNC697NJXen4vaW1ue
Ni8pe0mw6QA7olPDc4s1my2ygBSXtfzezh+Y8oGrYlbZSirhPKhGBuoZl8nrnhPE
ef2wQ3ZE71woGryc97ftjBj0AqSqvX6p4TMg4T2NEjppoArCd2EcYVAZuvXceUXk
jBOWL+RZubRDiuhn/sO9LLK8XjygjpaFyLiz8wygwFkBbygBnQTycTjWjBj/YnXe
On3BePhqrPa/598z89I+JVLcH6qpCm6IVm3uf8L864EsO4CyoeLj64cKVkm30riq
ibzohpaTsE7ivZ6q3wPFfS6UjnizC3A2P985yNhcRWdthtFpA8AtCYBOB0GiSriC
1s8m8pSDvKOU8NUfDH9Gx+MkG8IVPvEkOjrBuqg081vkVSMeMjAEjEu6QWlLg6U/
08spfUiU+6O3VXD2OLBjNO39jlV4l/L7sswR3Z4D0zxYjI3PGX0E3TmkF43cwSVv
oz5yZoinB0koAono7nwmhWOzjySkcRFlZhZRSYCzrPhMyyacjmmFN+MCq//UsY33
sy5/MZS3U/ZToHN6DaamKpveuBPngJieKMu2/E1bQeXHa3QK7x8WpiTbvhAggMwB
PpdJOmtaiFu0cbLog6HOzemmedGuJDp8KBQQz+EqJo04ocNSJxS/7FlARgCZ+Vfl
gkv56hx819ts5qCeO3pM0x49PUM+aZB0GunSkN7Dix6O19EaOH6Bklf+1i4rU2qL
9rFeWOdk+bqxEwzzTA/b1mAhSJHws/j2BjcxxRpWGol6kQKrsqVzv/xi7PJq3hWb
jVzxjsdLhJGdj4kyIVIcLxbZ8DYH26IODs0wQolYGHKlaLQMyxal+CRbVkE1+rAb
cQ9FGU6we0EBv2ZwYP3S9tifw3kjjvn7aZ0KeIYL13SCOimwtjTtCFOZJxEgqo5J
b7TUbGgWL5q6x32BC42nftjkPHJa8/6hvN8NBljEgTNeSDAz8jji9Loipz6jwuWX
TKvTR5qlCc0HBRd1wQsq4U0IH0k42//+Y79UcdN9wCxVHO6z7Kp0VxabC9V9cfTi
dSs++JUW7Z5gh8uecOL13g0rRfQSbs8Cyt/ZEJLGewzzOJfstTG9hBI5ZnIPriRm
jR7SVndNWuFNNki/moOUmZGzpLgILr9tkJB52YH4zvfDtEKTV3Al3f9dpMJLel02
8tAwim63/2Ps/289WrYiSRNrcHbfo0UuMHgY+DGV8NoddVE+q7XZJiwOm92YHC7I
DNX4hl+PAOuOUXkN9ftQB+OV+pdHg7T6M4Cw+2wo/uGSbbZ5LDmYBwxNJdZXclwe
okIxNVGcDo4ruR+FNN5g14xNFXvPYYwZSkvhpDXDK442iSe343tIAlhEqt2u4ohr
lyA5zQmh73QgiBz3BC3MOzDIfdQABQC/T6yP0tu/uDiKN44ZQe/ckIBRu0BwyKMU
bjdze86HzJ+xB/N49caVRue8DqCZMT4zhHCDlHjK6ypddgCGSiso5aOLsrV3d/lf
esslKiYHpepTMEuuidjQFTDkEezUtgIOjLmZm5vHYhvgo+3qPd5EgGp1u9wuwrjW
GnvZVipkxXtV82tmkY4qSRbFaXNnT5fSbXHyIo1P5rPItEk46n5Fhomy42Fo2OR4
bPL2DZ4CpBShqCYvVfXJ1aKa7K4MZ4cMLSfdFUTkArV5kwdff+KNhDgja3R8Q9wT
hkSIgoAiHAiZ3QPbTAdkOpeQHx1FzhKCCQIId5BOaXvdVgwaYDJ7pqAgEDx0fIaZ
e+YMcjIQRYXeUapMcjBA+3En/Q9dKhHZgp3Owf8JLPi6+UjXfQiRQ8tZFbcz83aX
xO75annDD4cv1GOYTdsKkCybDgLh63AP7lkE9cqirJl+e3piK4WaMIi3MI1rLl60
ffbL6ihMyp4AERFwN4R+NTEPfVQdAsq4qaFyQBEjXR6eH6PeC5m58FCfeGH764oH
MTJ2cD/Tk9g9oBiceMG7PsYkGUF0edbERR6qf8Qg6jxIHzOZ/Cv57IjSgjyTMahh
6z3CxxIeLWwM6xPoBe6Y4VSoboDR4p/XilVbyMQ9AqzYoU2uwsOhD6bRE+kQrG6o
DD92Qmff8D7fZW4vPth9T950gSsPcc+Xk5pFF1oq4FppzdrlR8sJ4AERcVAvX2Y5
pkFhHqKWeax8kQ/ObaGzt3PTVSYxYfn3pzHZOiVy+4olMAT4WRn8IJtrgvJLaKKi
zxaDzorpblbgnmcsr/AoVk02an3hWWDYSiwLDcaDkUhs3GV+VR+zKcCgZMWav0D/
dx76uGYnLUEktFmGLRgtPwplbGsXBysHn8a+Obxk2qc1RjG7UgWkzrRiNwxcbYuG
M0zlEIWu+eJSZ9T1CiFGPlxc2a+7IhZut5YIfOgNnRkL2h8BteeBkWotpaqRGPjx
d3N0w/X0n/JK2f9DJJDg6y74k4IQ7DnBnA/OWUceeSn/4h+dcPN20hD8ZeFQhWMf
APab+sqrAi4vVddkuJzYRPThH8r5mJkWEFTdQIyxDyEnZvV00s6YpAXi3wjCz6dG
09JTg9up3HrjxRwPZuQQywjxnDoLiVnQNgTihy8W+JaqZTEA5lqd9c3MiyzsxwHX
0VzvSTDD0o/MvXC+16CZu8JhM6m2wzkhJZt65dZapUjcRG/hELR13NTn2G2uF2/1
9jJzB6hgLFDTuKmee8v9vDszWr2upVi74SPV6DAwYNIIpkfIKSuRZKKsx0GFhN1u
0n3WxHRUhQ/y+OjdStP6Ct5kq7C+H0DFGOU7jumjpKP55vER5iFsyDRqS22LzkA/
2Xh1SM6iVz8JkUAe/yc9QAxG2qLJpCDVSkJN8ihobTcnc3Lygf0FLmuOhKPbEyPx
cFXFU8hICxDJyJCt9wuVH3QOWOo67E+ySJ5Uf0cOIZ7eeL1Jji+R+K1dBTzb1Uu9
j51BUJZCn1ilkJEnqLv2/i1r4Q8h2qExO04ckPkhD1N4o38AMYaRFdyvUdLCDDvS
Q0ISnkhpA1Cp9emuthwHhkoIgnJ8XPoqo4dIotnjwmwhiRsXwKS+g72dBXOyK/ed
52eb0cza4PZhj72sD663XcapqqciWZPnXudDDwJ/FWDqWKu7ZV1eHzKi6ocpc4jK
O30jhwi5T34mZpGHfWicDV7XKpOxYfhJHTAeAFbGV+5aGUgBa0QpMh1VBHj9QL6q
Ceombnzh4n/iA0cJzS9Qkm84b1iYdt2vllaA94vHhu1XyoOyev2ImhDiGoMS9xYo
OeZAhIku2/fC1AtTIM+Y1W3wyWahRF4dqTOaERdw3hHR4BF+gb0COidjCjxvQs7F
ZZtnKga9sPkSQLFVbwxC+4HHKwIynDx2wuQXwj+gBWlleBi854BvSIlf28YdKM9h
C35Qs2Mk+WlZ3yWqI5t3bTl0jfgC5+rCoGCF1u4O6KUFGnC/HMxZwRDm4qjPnK1t
BzEfGWrD+PObP7SuF/bZ7Vzw7nRjUFl1DnU/rkQFuQBsbNvZhxhWV2Km9ZbHx4XJ
8QbCgaz4pgj7B7/nUTaEXgl2cKasHCcCci3rQqUWrLrXxY+Ap94oQS4j8OCwrfxg
jC41znVZT/ydLrf/TNA52o0a+tChHV26+HcqUzmWbxoCVlbLD8TfCx6b/uZdVEZ5
xH7mk8wXvpwDz7ffLLLiAUIOpq1O9iEs3v1KJatScDsE3JWMyCw8ZhDQXTl/fWFr
nF671wvc86M3pg7nYLdw8EX3wuekiAxqa17UYG9SLxWs94OcOUtzJmo7tF34Chg/
FQ/+DvmkKEdgcCBLnL2tiKhYQx62dbbYA8JomLbAXD3+yvtsfBQLWXdEmrtSDC8D
R9c68/b2SV43KK+Xbw/ha4awZcwlGKbsExXBC+3sYfkb+D9yxyOXeXTgMia/44s6
lo1vR/QYHr9+0i/Hc/inyOdTHrrV0vOYonkke9dodb4crHNcb2MYVXWLoAeFFWus
XD6M9QuGSt9BVPYkuGoIMCAqXGRSm4FO/VbfxJKqXShawdsw0Ss5WtXAhCLwSZcl
pOBBbdlMc/nz7ZQW7worVhtctQi/sm4BNEC7iuj9PoIj2wVMFAgYi+dINZG5BAaN
UbPJs4T9UZ09fTZBmH8KfGFiz1ogLJIrvGecnTcjcN8eTR50B2aEUD0Fju7rGJ+B
+GLkX52/A8uBrz9jdlrEQBlHxoqUhOf7gtxYcIT4GhLy6srAPYr8iYtJKerdc7MK
NWNQrewIDSKQBdRH+E1BebBEKZmQ5HxWPbP+kXtMdUMHEyU5TSt8dEsqZk8XuHIi
iBke7ocLGwH+gBFwSeW4mUswc6V5qO+g/tmEd60O0t1VF1LihY/P8mIm0xgUpYXD
ev7zE/CoEUQbEEfre0W3XIkhs/gf6ish7dflAFLcZl1sbEhC6Zq0KtRYKaIH+xeh
Jj0vxWHIXMReUw3AMT7zOTaDyHImuVYLO4YBp/qP+S0VJnz91p/LR/+8cP8K4JXO
PVLDHKC7gHTwUFNP+JVQ7fxClLKK9eVcu6hHcRp8EW/WkipARDzvRdf9ykdbm7mF
d5bJmw9djsEl6uMbFz4in2CAaogyULoGiHjHhrNKCKRVSpUYob9cRB+Wq/Z7qA33
NtyYWE/Xj47KBbkkq+1fQbDtoIa2Q6/RTaUcMaQ037j9wAOg46sVjozY8RR4HDg6
GlKTlFTYrdU9s62UW/JIvxPlH/ZPigbfRMcpzbgsoAJ9kBvGkrmY2kg/7WUL/idB
1wTGu0VWZAtcCPT4+BQ+/nIxQvJfvS7briyvouu7vG8OQ03cXB7KURV8MVy7Gs9G
lRQBitGSzs59IK0C7ZXogkZbqn0kFsrcwR949Q8ZivSLmNREFoO1aUGykY0q8l8K
3uyotI54Ssd5uwRSqgDBdyBxKDmFQXi4ZKRWCsNBFISoD0wB2vS+SlIt1GTziZVB
Wob3Z8jBoX4DVk3B/SgHUncy0AG1Oz4wTIbaYcFq66xbnSxPYK+jNVIWQb1JY351
BhkSp6tk2AZbfuYzxSF4u+3W1+XebWyiUmEjPWuA38LCxkEm9TTHIGlpi9BhD4nU
LCXODUyfmiTmVFN/MS49/ogICBybiBsNpSB1fsgC4Zs/H+eTbbsTIbelSInx0xx8
2mk5l40+awyRknX+uyVqjNhZ1/0w7txF/bjxkwHbH+seXI+gVjjrLszHbfzLkVxP
GH7hsJthTv2lSJiTOYoksaQoPon1Cc5p1vvrV+gaGD/HEkChgnwkrAb65lBXycYL
2OjrXCTOYIlm20SgnjY6PEE7Y4neStDJuew1V29A0Tz39tOqjNiPwgqszFdw9e4q
AkJM18QPTstocAuqxqEaeOJbb+UzviKUaI8UQYgfQ3bLbhbXHJlEoCeikIksS6TG
aYbiHPXy25odrfFyAQxWCg6/jhjhXoQebhabBOJgT3oh63ovdG703gSCcKEa00/h
YvoJRQ2j8eHUxx2gVjouuY+NZo/mSXFa8TsL2E2/2FeoOL6d6ga/CVkttMTsXUVn
6hSyyzZyxtd+zC9kxzeaXgxui4tvCHB1QTx9CLZPlZBR44R7paMpgaxsuytazkfp
LNudO2m3xKYshGu3gZhgAHHluvO8pI70VVRQb/VUdyIZvFMYppdXK+aCmTTJjB5b
GuVRC1Ac7XhEhoqO0HNY42B+xbQwsxpIxk2g8TaNYw/qqcnJ/FwVssL3BCv93mtI
b5LRNsBQPb8Z1eupGxRILT+lthBatjSKcRayvddLh+yVDGI92X641fhlmDm3LLYF
s/sx5TmHLiBtROSNJ0l1ITNxLM90K4SmKebJUm9uMR/Uk/WKdgbKMO7qCzCo6SbG
uzbtFWSclpTZBzs52lYuyJ8Nv94Uj7Vi4vflBOlg0D+nNZ15lsp+MkDioZQcNGMm
uuESJo3h7OqN9nrO+SCtilMyq9j9H89fhLDnmse1qLw6tTkf+h9QY60BmDw+1x+Y
Jq+qPuS/jSOpXvmfGYQk3+iinPpL0EYa+SOM+AyEbdD1tNWwSVMvdLqo78xxJOht
7ywWvAfj8K8EEb8EIgyy1qZu8pYZZHwnxFVf8pPFxavYSgalgUqA2beMxqUGmw0t
5nU0gmFq/ZR7IShP7j8xutW+kQW14zvddnamAr27BwudsrHwAFCEGDcXyMmSIY9h
BUgFN6pHaB5DzcjX/aU/G9UI4Tyc5tWLbQqR9j1WYYSfm+Sn0GXpWzqVpnZKwJQ8
s3BLOcjyBsIEt14Mx1HcCU8qEBEva6mun/ypvewuGLRf495lsVUor9br+c9Xi2pH
VLCsoRwTHc5/1SnzQvltn+z0yS/TMN915QMF60RGDcBxICX42eK1RpgjRV4mwgaV
UfWI5P5pq3z2XtsbhpUX3Uo3yQZFuWsFYxHEDaPX+hOX/dJmtixJ+QZvPE5PBngG
FR0zuvI/DJHnfDny9w2/ENy+Mj+lKT48lIGKMANk/CEGGgV13UBjFSfQU60eXgAg
CbTJjeigtWJOASwi28wkvdqfDr7RCsORsfpmZFzTNCAS8yIZVi9hj2xiAW9Jf5DR
QU8vb4Wb6B7ntwn6Q48PzrE9FyVYGxgW2b7tCgzAJ8BuXRwSotHPVeRVLFf9TeWq
QXrtOymNDfCTkrMdU8XjBrkf/+QcAjOGyzhlYQNAMuFWlkDkkI3Kar+06hEyVa13
mkAkJ1dxZsHq0f+iNdui8n4U9f8gEioYFKOtQb9Qi28vHkTORIZQ9zWTRuWj4kIY
bgz+7+ipsufz4JFGFvrbOQhr8MXKp1OhH6KSvNxc3Smrvy8BKGEuRFwDrYUWdUhK
EWUnlevyfeYzwjxcDTqGYhj8OyqjC0G5b+/sqZBFkuPis8eEnCS8FS/zZRnw8OxA
sPhi2TIkA+2BAkrd6/kzqH9XxfzaSGQiWjDTn2JerYKzYoWRdQXhNF0GislRJ5xl
2hfTNvqm8RZDZYc7Wc/jDfpRvja/W5bcHOBX3LPropVmEP+FVXTFy5je2U2Pjg2a
kNnu/8rluX6pIcjRQgrBJhLh48SUjrHDakaCwntpMwDkbAQpt5bZ3oDJr0GvPnYK
z24XGIvpMWqK6xhl5Yg+ePoLxIcHVYwVHR8QIm4tioNc4BuxCDjmzDBfPDfq1gwC
lPalBi6E/hpDcvJ2UqgUGdBCgfelvvzWkU55QyOBjtvXxjDTr9tB4ud3rT/k+QIU
FkUVH3tVl9rYh79Ec6tKrylIBbe4q+z6CQYUWkXWCkNcOmlckB5bEEOF0vLD5qny
Vg0+t+okoUHFr8W4utSdpoq370u3Pi4WTbY2fJRNS2LYEDjd3fLpAzg/OHtfGxhR
UwS0v9XuSboBzdGBZacehje0TZFi5OSqDOCbJr1DjFO0KQwjb/cXBmjFuGGgnZ/I
xBk60D7eTvwH93dV/GmYFCn5qZLjJv0FG/Vm+LthW8CGTp3NJApylJthzdeW3Hsf
PrNhJ6HBwwr0LFgB+lS44NwVfHhHwjQfxtcUNbOktNR2EsBjxV2/+X9P/h+FxuBL
HSFsT+cGeK9KcskxmD0b0lSrUnKNEHi25CWXz0C33PrjpK0Jt8Vm6F8RsYcAafmm
G9dCyFPUEw0+1zrUsJO2/vOqz8RtdneUzSGZtRpkiP5afdDiirQDzxcM+B+Yhtlf
09iAXQQ3Bmo9HY1OrT1ru5egBhDpTv9EwR282IndbHdNu/YXYdNT+9Hclbac+1n5
R1xr2gDDsDhZBxccG/Bmi8r9LTqwk7ZV44C3YzJ50TBB1FnXRih97DtfSVSgq1Xr
085MWewqabILZNLIWVjHSf5APomf9e+/8LCJ4hPeB3fZdO9F0HLh0VCqi9Uc62D8
zX6HSbtq1nC4oZrna1Jl6do88ziwGL85LIWSOgFMceSBgLvdri6XIj3sQsDzo5Kb
0bxSxfLELYuqKfmtm8MME0xZmY1anqWttebwmKzRFjwskiMfxNiIb4XPOZwbi+M5
RhspDps4+HE6jrVj0T5+8DSYuvS6TxZwtJ6IRK/Ox7oeD6jtJ896A0c7sewaH1Gr
OsyTqCpGebVfzJ7hXa32eeUKlMX6cylvUDtEAIGPhjWD8o8soYRBspveJsvR4GEA
QinCEHcklEpmnq7bDbuw0ucwP33sBT+RJZUFM+e1YL9ztUeoM/we3g8D1kxp8i7V
3oJvVvRZCBZqk34KKeFD+7bMN1Ifolgvv4coqof7SNZ8GLkjNGl2+RFrn+eOszJ3
H8/S8cWOUZaHamHwaa68aHaz04gvnO+iX04SV03pwGGOQctbrbX77/h5Zrbw1rAA
WOBOeTFVADRJR1w7LTe0Rp8QdXefjwRn/R/1ym7Z639n0ob2Gk6PvyOMSos8p5hq
Luvk6gECzA5venHh7A44I5fJKEUnM3cezyXAvR/ap+7XdBd1pI8oItYyWEnXmUdq
0BaMWhz5N6T1+qrJp58mHMP2jHUv5/plbzQfzLqGxL9Ub+mwGOM3nnQfxzigbrZp
zH51sLrxzt8MMNyDQhUgDe2anXBkw+EKXtm0sfh5plv5Iwn0X9HgX0t2tf950UUi
dDMbPOD5E63Bps3g/mLZdF5cjyb/d3TbOcisvHb/yhYNEUZgP4XSZi8huBj1UUl8
ONvZpgzVX2MMtCLE1FBwwvw0WtduZbyVlkuQXK5ked63DKEsyobmnIQZQg5aYyzs
Hu/0686VHyI2YSKRLq2uiEKuxyUZ19lFYwlii0wFUxJ/X89ylxAWCK6WwwMwk6li
5So2lRoxqemq6HRMNon+TWW8HAPWE6mg9tgYTkf9d1WM0Zlu2EGg87OJXST11Zv9
h9W2vIQzd+3mXGZU7S8G56Z3iSyZibgX4/XHSNCwcINrUChzqcoKi00AWjlYJeH7
w/5E1Fyoj9EYtoraLsL/za6uEoOD51xX7CLjvhpoTWoODhrByPSGQusfftaYz45m
Ak3rbexK2S60OKHV1vJPVZf+JyEvyUlN3YNtqlKpsSBCQVBiNAR4e8p5tR9xVa+5
Xe1RJktEcNIVI561cew7reD0e+YCQn24deCxH3iIWLKrve9KcK+eVs0ic/Azf5vf
JRTdqy4jPo3CWSKG9uKMghCb//0tO7Rk7FzepzcL7ALQaqdeUb6HEMisAkFTcQLY
+JQG/y0NCeXbTkZ/I6lXrRwlUcHTA83wRQrcPqtI2608q3zy9WOvrCx7z3VPYxAF
YsAPnM2WsEsC63RAK4keClWAJcmcbv+fPs1mlkzLXhVW0E8Ix8HupCd9YFBDZG9C
ckKq7RqgZe8VY7mEk/mDrkeueh9XItg1m0+MXFJGJ3qo26ArY5ddsYr9lQy3NECq
hERusDb8iRnNn73Cw7oCmtV+5xFNQr8DPbww63i/NtjWvDBfXQbe2mpCPOBtSpSz
T/fi2611yF+58+B55w1MEvXDP4EFLPjgzF+q3TBw3HRdV3oiHYhatbyQlQzR7Izd
rlLiKqiHGg4QMPUceZ+0kuddGt0Eixx6eCVevEigUcDq+Csq+VQploa6oexWm0r9
GGhnZW8yEckkkiKhxeoW91xSNmiX6k0/KiuuQcp4WswUM7emUKmYc7k9N3MLbLAd
npaKFlckhekvNqNMniMMwupNlL1N75VQe1T0mH1oGzIbRCjM8Syg7iJgmjkImg+8
KezgrKhI2J0OF3WFghjTTqOWhIjTkvHi3+Pe41yZ8nF+0UERHTgeU5C/TKycnSf0
8fKiemXdKOs9vTV1qXoIG/DRJhhnDcZdEju2x462p7GrJSWeuGUHfu89a2bj65QN
p1uO4qwdlFykdZotjwux7N8uhxz5yZg2oOwWNzGb56hnfpz26/swJY1mYUeZK5r4
ymsWvv3Rp7nH5vrO+5qQGfML0n/tcnnBT/i0l0+zvygOV/W0/g/8yyRrqAiiHjnW
Jr7052AtXCntDeB3r5zxuKZmcgkaniJlVB8ysK4Am8F+EsCDZ+kzYcqQpo5iZLeq
5GJWZN5+R35+q7p3qf6OouzG216qoDiEjd/2MECNI8pc0+EGeqmWhXGHVgOjNnTx
QsmyMjw2tI2UJLDJ5Nt5HUk16MLBdkrMK40YRWyfIm240T6+v8QSl9yROUSaL8dk
OY9KtxfHOwNbOcTUL0kZctC6vY3Sxqo/dM/FzCkiBSv/kTvGiMK1fMNXPp/mhV9M
rhgQhntbYLErC4VBeKR7OF1zdcyD5ovntH2utUJTJij96jjnz6S94OBry4pnyWjG
TVbCZpPCCHah5TJxoYf4u0EJIkZ/Mm6c0v+IwZIw4n2HIgNoSUCw2oE3fK3P2QHm
dchzswfI1xd3SAMM1pDBVlN/hOm+fV4z9+KBX5Xkr7SXKH/j8Fl0TSqtdXK4TB4N
AV0VXmgcpTjYcuYatN7fzMnS3DdV1bEhQ8U5SPnMSukCNVXzLQEgTx4K7D6V9EPa
scvsxSNDAodJomlaBvs1NVQFNHyYV8rr96ZkJ0DlRzlAOC381LS4nX55lPHKrVL5
jTdWS0V3Wlsmusw3AhbmzlLVPbNVtnrW9u7ax8peXb5e7JAKtpdW5Li5qkDsbvgE
LCM4LTgQQncGTPxZCxXSuQmHw3f2qnhcQ0aYEwHYBwJjqKie1evVItGVgUo7olUk
m+jgwW1JuuLh9l/zbCk4rbmVK2CevTz0MCvYbdYOhtEadl3es0GQr5hdX9iD6kR+
YjBaDG4qKlriNiZVVNLe1AZv9kyAqQuhSlxKUVOfw3xfmeDdepVNzTFFgQoNJdKX
8ZmLU4+OY6T0MTxn9fmIiTBCQaboMW2pnsP05qK/18TlFbOg+AzDrAD8MQM6z/7s
oyJyYKgg8qk51j31IOSNlqLvHetSBhpVNOlEIL35LihtFQRZVOdw3c17u+9CAg7W
UW1wY9NGvVSXB4pG1+Zf1kDkvr6afM/cSPixrpvTORWRvMldTI9RkP/RIRC1PChK
BzkoXgQWbituPS/rrBWZ5ykcc+ZlE3W0pBHDGn/qPFdAXn+cOKk1NYimmHSueUwD
4KBBnQaFxPJIOs+oy//tD+mbs+hxDTKSA9rPwpWzNF82bClsX3dM2FwW/BC8vu52
gA3RjjwAbDR6P89xzZ5hw4334QYFqc8uncZgMSwFqp4QF7PXRgl0fF73MlD3ehao
dH12KT2vSTwgnuk4EeNsoeyY1rlyWK16e6aAULS7xCpXEQIzK5fbQCxOmjJ4yLx8
pVhOmYsBTgzvu1205tgBOvS2HAiD1sdWyM7KK0EDWk55KwoARAPmFBrw0Ji1DfFX
s/WrumvErkHL/taqTM/U+PA/SHTon6dMigFeIpxPqTqum85PMqWDpoyKcPWR5dzb
F1PCi43KJQzZsZvLsMtjzX7L/CCdLS1jxLRAWWkw8edq9xXfmdBYpE/yU3Fwk//x
1kzxGPBE1gogYEVAoWWSCyF8s7ljfRqCBu+ZdI34IAAPI54DUfJVoZ7zMADruN49
W7S8RfwdeeMYjEBQ2UT7nwOnfo+QNDxvHAvUzUNYonj86GtO2piLucZ10rBCpmWd
5cEsiqt6i4NE8W4hwnhX00Cmk5jE5zqpxbqHP4gwNAJqX/xQMkqYqkxzswqaCc2j
BsBTDSeeEoOceOb2FwLalVs/NseQG4NzYwI/0+r8WtAM8rLgQ4g80i2faB3cX1dm
Tx8W/LDq0FKKbQWZIw+jI+jVKhJ9M029VQzS44g6O/sSBFp4xWle3VTgXE+oN5+O
tEr8X74jOLBK2EjMzlczsQERXwh96iDSxK91sYNKEXxoWfnyvNlfYiZDY/mkAJ4P
Mgx61lueeeBE2ifiBtK4zB2A+4ljnMx3rrBqy4CMIMnZ+maOc1j75a4Xn6UhCqyP
t7xwTpE/WbAVlZwrViRIARa71valSouhqeGS3sPJPzzXYH8p1s8ARBYUiPzyedYm
5+WWJUYVkhaT47YzPjkeg46JjQZGtjhGb+acCSmGLitGPk8DUAZuQ0G4J741FKvO
0JFzl/hYKmbGiOew57H+uk76zK2nR0mqZRVfo9ngZVGGtRsmXRGZvoDutm2uPwv0
U99wv5ZMArOvVx41DFWeJ6ema7mFcVhOAHn2cbJ3a38XSokQlUwuYweCuVv1jSh+
5U9jqaKJgY113s6/n8KT+RlDEY64Mh47nztKQRYoFnSkSC/IWwOIfJXLBJRYjU6s
LOw8mHsN8QD5Gs+MnF2YmAN7+JLY7exT6HW0StvUgAWUeZGBFdWQ8LK2B5p3BKU+
TmRaSdLUK4xrWxIDSjl/4Yu1tcwko1LqwLhkyta92M5eTWLitofqn7dltVbJjeft
NDK9YfuMUjZD5Bbe5ZyGFkXq1A83H98W78rjHQKk2qaViX01BO77ZjtIKDjwBdbl
DdrYOZ3P7j/Y03V/r0V2Kk+ggpDZ481lnlSNeRfsi3DpIiO6XKhMzf63ChDofao/
YPQcfslc84yuqqIBfEg8EzCBU57ax0uPd3dOFqwpLNf2y0HCztiNpp7hGgsUZ7YK
SvqWDCNLEQAaNJ1ertyz0oKCccvovcEgYefGVxvO2k2c8MKSGjXlU7HlJgcBxF2K
zfOfwUJmx26Pa7aV+D81FD4x0BIp5/txoE8lP825ho9ESK2s4JKyYBJ8lTgklNvF
hLBriEsNesr2Q37ejbgiooews+EyydGJdNAck68Bu0JyA5w9Zo2B5wRl/1HSj3Gu
gZTPDhNtqby5x56KPJOd2AVTdnhjOuCZSiQSfGaRfRTQ5b62Sc8FpAuSeb/lGIYY
FYQr5i8omedhPP82u9LOtYkGRIuULY87YPwE2duUpwoG99QW8UlKC+DEiwQuMkO8
jpmnln29wezOOf9JQvgLEuHc3tWUaTysmr6uZsokdxBSJHSc3/2EbyaORuGJ//ZD
qAwVfNCGxlGtTS697nYrosKo3KShQNDFdRwvaeM/LADyQmd7TVG3/Lm8txfEmkdB
/5+Ipj/fSXVt0GytZtYQnfkDjMRDDkVmBm2Z9YGUukhaEtZ8rmPcIYr73NS2jbx6
z5TbzhDGwHdw5oGaiOMhmStLPkbQ5FafIeEOkhFbIdAEfvY222Y6b5w6mcjwlpZz
I86xQl43AUgGL+psH581hXZPJJq5EJ6yvuihBpoX8k3WrgllZ2y/4NFFzPfeTAlM
c4j7iAhKbPyFohamOE+pGo11jricMk17r2rxC+7Cmm4+k259WNyVHEKVNFUVb03W
lWU/eTtirMvRedSKIygPfFCzO+LfxyXfxzdUbaSgYN0VILLOiNrft0wOY7oCNb4c
tPsROb7Qz2KLSjorsfUtOZF8qi6MdSVDp//seiOJNcsqMIgU5b6duW3MBn2+o4h9
XVWntZnLoVJZZt2cUv/81Ku3uyscuMNilIVulFgoZnRpznzOuuQnmQVNhsiETrbb
TRq3c8rYQcxYgF0o+8vGNZwv5C92+rUXA13ZQFtz3bpeTwRntVfzRpmT6djQljh/
3A6qvJ0Ui67N4FnhuQgybAsE1NwVJFeA2dIYK2maqLV/htGDR30h0ot80aEse8ql
MKgnfWD0zu/lW3EPJ7A718fLCBeo1ug+7d0dCHNYhcqsOubUhWhefg4zXrNtYmu5
gnQW03fsXzeMq/ZsJz77HbtlzKkf5L0QDZPWu35sbmGEH6Q9Jie5yho63PHe/C2z
vtZVFvlZMR4Lk+7+LjU+I37cndsOQtl+ylaYeouKmvBPuU6jXiJXnmG2s9os3crj
6DUQh6dHOtR9YZaaZgax6A+uXv5/xDZTcEiv3AyS3CcnFle8Pp2E+VjzumlGEqCU
CGNxZceNULERa2IwCxl8SjDrkNIuBtesoyeIEqFVKFAhWOzuYFkUGhD6ffqD4HN+
dGas13qwMPGfAWRfYWvEOZs9NzaCw5Q6hmipEmuLX0I2DKvHBLxEjlicOITiIXxZ
zsTtUP2cKC/d9DOoj1FM57fr/voZcXfc9lB2No9gQtgWc4wsS+Okw7t0gyaBgig1
3Fdnix5FsNOjhVGrXpAyUk05U27LDu4kg2nKGWfbr9IL/ss4/lXryWhoynRFr75X
2bbd/x+QVJQLW2ECd7mcSH/BPMYiYIDv4SZ60kvV8i8B68eGt32U9t2sgMWVa9Jn
0p3vTyvFBoY7/+XsipL71D2pZMWu5c+K2Dy21FdIuqVVkTgzQewYchNJKaIe7mjz
TnO1erU21gXY5sU2G2//xVKavsGhG1XDnG0461OWYRRv1WkRW4Ii+l8Sh5neC/WK
ufR0zLj6RaJXrohNHIpU8GLhQVyjYCGtuEmwK0WH4hWapIq1KUTSV4xmt4aPgj5A
IAZC4SQxfC2UXlRJ3UI1ieBdRJLv9rB7R3QuUariJMFDy4S7Gv9gOm9udt9IVTlR
gOcA58+yWq2k9CyiA0brFK7nMfbSoV+b7wsJJT9ShJUk4oTXnVuRuINB5xpUci/f
PJFGzc3K0AhM2K4UCichnguNpPZMeRNIp+05fOI2beWchNP7qw5clqSKGyYBeLwt
2Gm5OqXDneubWoXyDzAeZl/pZZ6kkWj9kVuLazZOP+qta3oK2UaCgaIbedp3bY8t
Y40SFK3WddsbR5q+ESn4B8fY8f0ZD5nJdTslEAmU8yLp8flNLMWytfBLLLeRFesN
qBpZ7A3hj5155ADuu9E5Aw==
`protect END_PROTECTED
