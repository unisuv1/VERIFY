`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p76TjdJRxhUHfT60HnEC+57sgARqqRiv74GTaWR9NS/KoeHGk4Y5DxFAdTMSF2Mw
L5Wc64VWtnRWmGna5Q1/od6k54XPjjv4Ggf2C8PZuF7KzXY9CHBdJy7/yNiJS2ln
/CYGpdVSxRCYHbIRhArsQtci0uGQigH+zC8gCBCEnZXadZNZ9Pjt4i3Mm0L3TErY
2/4SrZ+Vwl8Xxq4hN+JnkawxhvpluhxG3wuvah/o8Ihzz5CsCaPMeh33ro8NFP9k
aNq/JI5ZPh+/9I0AvJFzWuvLe+1icQl00W0UIgLcXcDgxKllNAMZukY4AL4BG4n6
73yDbW6zBR8vkjEiXh9WjHI2jdxFR7HO6r3MMfbrI2Ir0fo7s6MWYRApN1CgZJlh
QEOH2EDaD5cNJoM7xBuFMvfsb+J6jgNcPJZIxJeAbWfyzN3kwj34emaZFS8HuN1F
3kR8ZPn2W6d6YP8cdkCaTSQ7wvuaXvwtabXi5W64lRoPoJ3s0ptK/Y9tHG94aZmB
EJM5/B4FsYqr50rCoXv61kEUelmymLFyXz8S4EeG9WR0OuTVbl+CxZQCTopYGw/9
U/E/LK/G6j2ORcoIPRd4U3i3VNyp7Fs0hRiS3F42BnT6A2Cn3hoc1cZ0OzwTQsZK
EUSucmyYYwLQFlX9Uk9Co49yld9WuM71tAJadC4b/oXHUW6YooERn/LNBu9OyvLA
zP4KuyWJBcINPGDZgU4wSli0ShqzI9Om8ajpRjN5xPBWom2nlXzed/NwynrIk5D2
+WkL3QYDdEJ0BuTfNNXEiZn6I6FL/DWnkfRHLrfLfirx0XCMztUKM3MH3GTb3Xo8
pqX3TC9nGDPViokCfITGyAZ8y0yXQ6Ias3ZhJAjUVYBM0MB0rY4Eulw2ictSsK6q
ZSm/v1EAiV3QhN2XqPeI2OPkoj3+1nvDyZaTjtLCI3LzCTa5rnN0u3S/DSqQhB/n
NY92CfRuRzVBTNrx5h9VbDmFQLMq8O2RgO3g9C401WT7EinVbk+VR35padYmQoFa
It3roLVg8E1RVlCBAK6vVOzGCup4B0b9txqeDWlgEr0rZg9vbRKj6QWXuAdZjD2X
CNSYVaYPinzx4l7x3gW/C4eKJeodaXefGSiuwo/F2Fhik053Seis38HnuB8mzrYj
Ksz/Bvt4WVbf3ha26nuC8rE49FOkRnDRKkIl1e3F8MCCoSRF2daSFLwEOK/36zRB
DwBqnEtmnk0XqnywgaIe6zb1gKUbk5AhJv5W5do8ZxqSk9br/hTZwaF13oN1fD5h
wR5R95bWXtXJiqMdQbfZOb9rX9APMaKtHut5qmv+IlxEfIbWObMliR6OlQZAJgH+
/U7wRaPqxtZSroqcnXpx8gGoGPvAFbpn3Pdc91BpiiCgIl2B+CJbwi6mQ8hdc53c
j4WEancuU5A+3Yj1L/TxPph29Zq7Yw+6aCKkCEcsRIbroiONkK1MUzj+S2dLT2YS
umIEFsoMsd0/Heo8qkpxKlIZallEy8wlz51q5blA+/vMBABEVsft5k7zdBdt9Zn8
QnRKohxGv5r1R6qWPjvK75JFgn9csG7sRCPWyyTahsiGdazKFQtLkxso4SbgbZQ2
q04I8Iy2EfxvXCSj++/9CHNJhMAaUVATlHtZNPj/5OV6a9TQLCGL2CgI8NlizbFa
P1Uyp9QElFJb6H65f4hw4TxGADbL3N8B9w/ZAKh16frRyXYeKLvcu6VyzZqesywq
jjZXpqVy8xEzE/xixK6q1QS3GoSLiELI/tsHiE/6PKfy+aM6FXHXaf3w3dpRySqj
JOcic7abeWXjaSmSN3cGyozyAHRuwnnsfvEO9NQskSiROMv6dtIT8RlN9dGm9f35
JnoxLp3MKjyBaOwG1ccXIToaTTi7lBuHIEqyz/V6m+OamzQcwrgAaDc9HqXFwcpG
Hmrk/eCLAq3Q7LC6Vh6XBpoQE+BogG5S3vZLHOeELQ+Zi+D5FN0AsZ5i5lyqX3nH
73mUA2q3DXzj30hncUvJx7B6gHFyLhFrCIexR4kV5TQ6xx114CCbccnnpHsSmuES
8706EddxEJej+F5l80rNo3u3q0Y0B90QPCbwIXL0qn0mXFb3Z0Oqe0+fLIMtelfe
mzRn8c/VeEkZKvehssQ/xQ==
`protect END_PROTECTED
