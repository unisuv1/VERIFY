`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bB35ssA+pTWae8j9+VBNkppz9SFwOGDNOkw+vJfTu2Talf9kDb9SMZZeDZeEuP60
fH5+CRpq+BWiX2wM67k0mpu8sWS0VP6PbsUBzYZATzVt+cfleyiG1ojypsU3hoOA
I3+BbvGw8sSJDqddcS5lKwar44sXgvKxgqlFzgkQDK9GwaTp6DwxegRT+DjcR0B1
KxQeZ4jp4PGNG7gcQvwcDTwd+hHJINTbwyDpghJZhFX08wOu9if+ftgfdlRQuDj9
rm3x1GkTLI+mU9ognrUYVHwKbU6kFaOCSNpbEynsoK+Yjdup57sZsiuxzVbBLrUh
fHPr2FeHmAnpjOzVGZhNavT99Q7mfrzH+TC1jTxmLPiHZGc8cf+gMY3AhBAjHaQK
LDvUa2AO+zaRc0LY9dgrQHaJMvyLxc0EqxJn/DdlqKWpj4lEdU1HY/J0dk3Ms3hh
QoaIv9ZKinMFJfs+BDgUTfL9Hc6FpnoWP1KestCbDO0kkSVLaoIHagQtc1OXw/cG
DNaMeV8SBM+1CEYrDR0mqhSXBJr5m10wSLnmUWdbzVlYJBfehEeudvSWflwxEnAC
gnvr1qfcZKDXslVYa45Pq87ULJKQPPMx5pwBeKK3DJjij64viDUC5QP8AcQ6gpRn
qzen9yiJJb8SplOPvVn0aj2xgGLlvp+NVJZ9o7bbh1afRt7E/+TNG3tmrdF8IJ06
W8uV4VgJNjQeI3SU5BsezaKycU0wB6gc8Q5iMG2D0NFOmaYdPmYXiFZuKATJuYXh
AyxiOiXaP9wmosASEiGqFlhD3kbc8gwAhhH7p6f/GJ71surA75p23YXHqk+C71Cm
xpT5kwQLwFBG08aY9oV/Z6JsWHWWNljVuRXePdQc5k/8gJYokrNzKmqrL1AVKy5F
kyOrygkaz3O5OHe/eY5GBtSwwHQUMrtrSCpOyg5SF989R9nLzY/AigPgJ/iGYunf
XcAlZYDElI1skFy5QP0zzZRb31SAKI/F4P3d35Qs7RcgCfbwCs7ej2W3TQnnP1l/
es1OmKJnp2INjp7CYknzeXevrqlbYtPuUsz4G/bIJ0ykON7cqc4SA7IuerpF3o8M
TxIhf8DTfgr1KFU9Jo/2lLYfvtiZns+dyPti/iZy1EPW/8DuAAOOxMNn1KQYG6rG
7OQcZUGOfANgqbv4FnY7uAcxGS7hrwuaf72knw1+RtO4GhkLwmmipTVloQPaKMxx
9Rf6ukXA8JWo7UdwGxFu+azz8y7/h6V9tQNwvZLyEDq3AzP0IZsYf1Zn5/a1/nyG
kukDHR2VR2gHc47ci2GIOlaYnC/dZijHMRKlExjJ3rhl1B2Jm0UMwg5f6iI6SD+w
ymhAh0scuxkCtVbHng1H5s1JpbTdzJcFZvUM53sE9nCKEgK2Dvsv30sTxqCtzSXA
BPPIyZgOl+AMAq8p7QxvDOdtq2QxaegLjNw534blyq4uz7uMiHKx2/fjEpdLyL0p
AQQ1OA0dWr1LRMSAxfwzc1g+zQsno0lfyRkpjLZOTYc6B5bgdfvlMtyEekMUKT7K
CfVWfPSjPERscpSKvqrIi8hDmarK3X+iWMpnw2JBudT+Edigs8w2BX09HwUJyn3B
UFKaDGxCixsbdkR0avRff55uzKrdZUKmt42FVVX4SQP9cB2AtQBegR7dqw7D5gmB
wmTBbD4UQqJQ/NocSIVaMPRoQwFbEGik5Ulr3vvWNXYO0dCZ+tLWmFHkCvuq1RaD
p+yvpX7tGD6BT6qpc/84eI35SrYjoDjKDxGCR6uezYwyeSQQYRUuq6qf3oNU1pzm
WrqQSY3CdhuU0IgT8VeL6fw+JKcpQueJSeGNiwQfSI54FzzQ2OQkhzdiCmF9hDY2
mxts7w2bmhg75iPIAeFlQG+A9Rb0eWyFGPaXhm+ViDQgDVMgq7HM7xHFw8n9VtFt
/dFrEGe9q26aHA0m5sZ5RssanFJZiPW4MAvucE3hrxxR2oZUGg2h60nlkqnIyGj0
4uLK9a8wojo+A7w5yigpVV646tbVCT0I+M0qYFb3Wj77aCL6HffWZFb93wmX25uK
/pljUGkCciEq+IBO2E4yL/z7ptw7rFCSAd6F5XdAAJMKeQYJd8plR0RiwTZGXRGa
F9XA7NlTbmkObFoawh6Zr3RYODDVfObh3fjf/bcRF1AcO/t06DJm8cOsSaCUbvuH
ewFUwdJ0OEgimZBIbxX+vxVxGIC7bzjjnQRCS27EMJUxGaOGz6vNKxxxaIPopbEL
vtHYSU39WBFvCeKyRy6eis80bZrr3x/iVOUUxTOJrowuwmjVGbKJPaqCJxIUapPg
8E5Q3K3LwKzd3lIfj89MFez+//bCfw+E+FQzn9fOgPnlbxkUWxwgLp02Ri4vqyDo
TXg2YBN9N65KL3N1b1uxqm6VWg3ZmqahV6e4+kP5QhBcWkdzKSY27bL61bRw+524
06v9qYU+QIDfMvtHlxbdfBfJViZSfQxjroqJhtPiKK5qkKEDzMPSyWjYXkIe1iny
IuZEDKy3xr9OfZYZNYSqJ8LCkOAJ39k6rfXr6cuxtID63jK5Di8JZGeYgAoOUUCw
XGma8sqoY1CQr5NuIiDA4AHLAgroS6H+550cRM6lkqg=
`protect END_PROTECTED
