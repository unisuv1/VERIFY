`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bc5OLqN9FnYa3zs5GpAgeUmoq7mRjuViQClXWLNy2gFBW67BMA1G0IjAANwQpHU2
Z6uQC1613bpxr2MRyx3BYFgXx8LXisa35l8e1TNsoZ3MNkE8HdkU7LljHExQdg6e
6GiNLOBmz97ovgoG487vtrnQioh7y/guYLHs7tQ1x+fUVCzWHV4HDoR+kuCgG+2R
xBhY7coc6ixIIppX9dR6dp5NG/sUpSsv4ArY9C1b2ZK7QbdUU8Zk8ybH7f/9Mgo9
NjkznzoPqQY9mrciZgnWDMRHGsJ9NyjhGSKUFvCIowoSO08jnC2zq/dkfUfpHYQ4
kAAvjDIE3pt2jyi+xfQAJVn4jU/Rm/6lD2W4Sk6eLXXvA0iSkPoSeXVXn7G4jfOZ
q2SHLTl9RADNmvaluNKKrRq7nvHH7UbqgCm7nG2ISMBdZdlvtilHWGLD+WsHTUgQ
L95Po6o1KK8y79+pNDcKNA==
`protect END_PROTECTED
