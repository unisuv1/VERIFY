`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ItmX2AvFBO+D48ezevzRBxCXyEX7t61RZgtqRpFbKGLo3HY/5cyXRwsWYTkw+Ts+
4XomE8Y/u8UtYEuxm+dehAzEXEnJyG6wbbqaP1P/RbgDM51W1bK7gFGIJj0uI66/
U9GNcLMrjfZX1FHYZ/t6JnmobmQEUgW8lWuIOYkDps/DoYaXVbDycEDTsZ8YAzTZ
xYDLruFB7lD8IeTB7FmuC4i9ZlbmWjFN23UL78r0HNgvnPxXf2xaof2zsOXyOV6L
hNLu1YJc5hpNd5WWlgDZKIcr7vEjfhugKLNOENIofiGVx++6HGJexur+EEGqHZxh
bvs+alNOhsmxurgAskPEHdtKsX956qkaDI0oJuy1k9m13Q3MPrGZk0OKuCGSaOPW
DIlAwBm+cvmieeYqFrKXlApQiluCFKhqRehijiISA40km+zPfZC9mo1XxWZjFsPO
lBxqMyTsXm4iPkt/V1TXvq9DtrDcjyS1me7TMKHkFT94HQugPjlJFVjz+UjNJMHk
TrSFA/+itDzXnbbTSwNLtb+MsS7gZlyGIsHn9sPP3WFDcHZpKUwX79bkLMlELdCD
MsqWXdvH2xPvImAu1QLUTvUZamr6q/1Vj/jg8snoTiG++xAshJFMygoCNZotgjNM
pYn2QQZY9Hs5FovsC4Xl4y1HidtRxUswVkjwkovkXyXYKKeX/wEpMfkE7WYHko2f
pYgiiu/3noQGimyUmPshOiiVaboKxek7Ua2KjA/XJJ2zceZfz5IvaN0lrv3hlBqT
rBSE71tZ+IvtSr/l440uKRa/ktyu1l+T31e6wqX9+Mu3+BvaaPkPsBvdi8LM1CXl
LDDtSCncjewoyf/c+6vn4sBieKnpTfl42pFylqoGRTvvW++pz9q8wY0IRfIvJI94
/uiePyqQr/3x+UmyNOGr/Btb+ok6gTYhSVAYxpQx6npHeXDqux2vFOANyNt48SBe
uPCnWEZibxtYH2X/egjm7KgY6WchzmXTIxRA0z8lEeSdhZLkfPCgxCwJ+sNUrvs2
rCka1D9r/Re2rxN1HQrL2zIQaMGXhQj0Pwmj8GTGTqJ+ptJa/Wc6YZWAZmw+cp55
mEtTmWqhRBn3wymGUc0Z921LiNsivraThPeGxqKzV0Wru3Nsnq8M/ldofhB+Aoy8
Hk4ptAbZp9tScJzMITbBxGGSWQ9UshN2JmgGWtb6gDPKsFWXb7FcOqxXYoxv6DiO
UArv+6XX/YOUgQt9urTcRYGvC6MaHBFkHyIVyM/u2X6NOTp4T464tx4aWxr5Ci//
pW2BljosCM0lukHmdXQNJ9/Uw2gmGtoPGnGaLwQVvXEfR9KpK+daP759PIlGlyPU
yxT5xhIrF15zLeTpAdVKnS0WZXXn84LxvtEEf/1jcfYljOT8fe69t+Ihuo8BLku+
gc7BtBgpWVvZbQZq3K0dXcflJ75vh7msuwNS9brZsgPtsg7zQVcn2ltzTKVE/DYs
1anFDZ23CtAlszizU6wP1gTVlp9/GYENhxVjJEvuHPARTuc8IzteJVMqehk4ZyF1
2cxubjcC7Kg0IkVv/EN8geJxR9l+P49Sq5fJcDgNah4FPB/1HZgDOxaDDcv3bjvM
bki4vKVqcgR9U8hFaX+kZtsVUZhOghRSU0PYqdkLykhrR9VTf5a+zDVm5dh/KR32
PTwo+rNrDB/tGpvPKmB47fioDO9d+Fn+iqw/OzReO/pdlP6Fte6ParDw33eJ8EUS
6lmJWP3ZO4T+ZKF+okHbPfh9FX4jBv1eZvoACYXVQrcx4aQEuhE94WsJa+XpuIJt
7Ecc8MX8eK2CqXr26ciXkwrP2NW0n00xhpJje0vqivUFXeHTriokDy7f4dqFP71C
692M4xYA3gUom5cIL7udB865x+GAaQgBdIomoGfebD2b1Bg0IB2UUpkj8A1YRLvI
SRL044Bnv9E3V92dZQR+t3j8EKGQkb619gIrCLNzj133Rb3Q8D3Nd7xLux2Az5sJ
JoeBnAIrcPld2rqvcFKOt7vG4tbPaAmd+EymuJ7YhGXaugRsvcgQzedzA/4h5szv
vJ7PuCaxG/XO+XnUc5NDLnoF6/Wu4ZYroBb2K5CMwy1h7yfNNXNLCvSGNBzXSchP
B689BpVCNECpAZvcgMp6BtsXIZEUMPcE0CIIj967Dpgf0uBrzLMvYwotL+3phXjx
WFf0uAFaR34svx/c0iooXApBOyY8sOg9IjdQ0ENfX8mKB04IXwvHY+tTQxVal83B
B6I3EA26wtyFPXFvL2CRPorHmoB+R9OpfhEKgkFm7l6ku0WZT28N2UCn6KsdLi/J
ccybdPVYU0ircQqdy0xrZQzfdQ30SW8mxoSeNm6z7ttIe+mmeKMRp2ieBb3k68G3
+tCc7bnVcngHngaJf5Psby051D7r6d0hBUPPvHOBRF0+xmKaU8bOe1Znok0l8bd7
JFYd30eCwY2WhYOwpMemiFuGO4OF+LdNgtxTnDTWrludbKhgYOblbs4fN5cYvabI
Rs4NpDvTLqjmRBiAxD9UnxUxKAopteRd8O7V0FewW4AEyDuFWy1uRa7itg5IMFS7
Vj/MnjW89GRglqTprsx9m8cVugH9zDfkPTg3w3zlLI02mlJZ2XKtUGMpm5EiE/SF
SCfGGQGDHxWYwgnwJDxQIQ20QWwgh6cPjsaD3WXl94WsoLwhva+Umv6o1sMLEw6r
hOsCXyH4NVG+ob9JVAdv6QGrtIADNn3Pp8zmD/VrkC9zGPUKlM4NVAGIbeU9RjI/
Q/QEFH3Fp61hTZevMVKyNXnoxXdAWOMYkqgzFUFyIqaQgt4S/M/ivlb7M1hx5aTJ
X+i52GVVLjlPNPJKL3smD8OCpcNTBnxCVkjQc8TgHbqVhzbaHAMKVZwDyUQ66hOb
3p7SzGzJjru+FYvsMXJiDftCnFRteAPd+XvZ2k/Tj02uJjO/ZyJVwGh5+LFmt896
VZRat5XuPNxdTsXIZHgdD5+EhcV+FkTWEdY1SNCjUk5zUFeeJMGGxZlh6R8xaX0a
9Z70T/UYGLdgV+TgqcJTtcz6zjh9v2dV1qKDK1cvTHq5pVhyQIF08H4pT+rcCVz8
8f1DEHn0RuMeqLUjprqMIoERBUh7U3XCmVevJ4fscEKEverO+EJpIJzQHqNpH61f
4/E6TOPfkDjDdKTsisiuH18fRBqSpKt98qFdYUYsqz7SZDkcdQSjbxUSOkWfwbaO
sXzkCSRpFWF8k51piZolmcHK/W4i2auwpbHANpuOsr8Avce1Lt22pPPOIkQRrn7Y
HERJyWz05XVXr4NNUpkkOX6Bc+ljRSwFY++bd+3qSyMduK+4OPWck1RofnqJBvqi
pB4WV0iCTDaP4xkESpKROXM7c4g4CxU8A4s0ql21Z44YY4nzPVdztxduusUssvz6
7xhZNurqLfih/kfky2vHhrc4YUUzIfSvYNIkj3ZfAlroYMgHhiMvel3CwhuLij01
uF6FxnqNs+rClwJF3GzHLqej4GdKI82Sk7ObTtJA3lZygKoAyrxBAoFMg3ySG95O
V8HyQJkyJqZdyVe+D5rR6u/MNLbIovDmuxGGN7Zki/1Mkak/mvK28q+GPYskJjZy
tZvLHffha4WTWVGt/LsRmbeKHdPzf/RpDkKtAs231TsWITYIO8sByvll7nm8Kqmt
LEz2Qc8DbIgnBWxu0GhW5Ohai6hELAFlTlt9ZAyz5u90KZXHPo99PWsXRJpguPWK
p7sxc1WLeWdvizadmZPzaXzCh4fdkeG9Fz4w610BpJoxuace7YsPp1h/IA3pikv4
CH7ekXmMUeLnd1L3Utv5MJG4v1PuZYICigLBCAo7Xp4UCYKpuhtoaiiWfAVbZ0lW
fDivAvaQhjKXvtR6PKb/6UBMz3sgtQrJvMXKk1a59Qfg///ym4szw8iEF0szCKe/
2d3kzG/Dlrvt/TZgUE8xY/O5lfTkCeLZ08HxLhtUk2JdNv2dEqG4bdfAWV1LxLjz
EL1+kRHZ/FT+/ecHVVpH65xf9MGUjpyL70aMGBf9XpwByXqj7/fU8BfgsA9eX6T4
GMnZTA7lPXorAk5KVWHZUFU0O69x+qKhObHML1WJSQhN6xk2n0VUxyWXnmwoRhT3
GikffKetvg3UYz6jtOkGrnxnFxdPt5LhoesegEnqaUFdnqeUIQxY2XfE8vYmIJ5D
5A5akTSS2Capuqi/4ZA+sNiSbj0Dj++NsMpBq2AycDA0SlXQkdWoAaqAxauXc1/W
y06pXqqmMXysPg1hXl4F6L99U2x//Xy9BF0Zaanffw7+22fIJFgGoJbtStSuw2Hu
4SAUk2JoloV1lym29B9/JImMZCHIKPY3aUhkkYA3kxszyK1KqdmuAmdwJCwDHseb
PT1Iw349sBimNL3Sbf4pCqTxX/CSh8r57T0/50RJTMdw4lcXYomFdnDcS8BjrsUH
HlIyqgXyLjTW5Z9VwOd2hK4cJAijYB+fTjfdnvUPRlLLIVIxe+M4tjFWc/9Xmiy+
xy/mcSuHykcN6S8IlalrGTP0PM4iEnQDJ78hUTcd0/5YL2yzm/L4AR9IwVmILCad
wvFKQriaYFqLn2I70duEJ7WBkxljMZkH4Xdbu/oUO2WXzFP/xYDouBj5PAGL4GM/
V42UrFXcJobTecTsvaoLAIRN72eXcpnUAL4PkWDz0IOYMMP4XjAz0zgaEIBIY7hh
xNvQ3xsmSvT6l8kSmDbAvz9FmMJbnjuRPTwkgOZGObvwgO0wjzpBPw0GnQ6QqeM8
1UyP0tD0GVbnBnLbKardhsy0ncS0RHdyVEjmysJkuCDS24g+RpIWI1DeMHQnO4gm
+nSnEnsrXakiad1llNARaUQeJuMnf7OSn9b2Eya4OsdiXSF/akh49nSAm/HyDX1p
RQ+JX8xfdScQl0FH/HneoFirvXIJk073HKZOZdQLdD3nJiDVzRxuWqtCIvvrudYt
1CwHc8SuyFu/860JQJorHhdpnX4qSPLf/yb6KJGbnAnwswDumOWKP+0eTfmDPIJx
OGCIE9adj/T1fKmeLkTaq8SvrojHxzSh663bo1O0B7GuhBljXSk1/DvTkrpVSpgb
yfceMsCN85AJKLTTxVRdMeQvkoFYdrSky5AuaT23Tg8bWWUEvvJG4Ff0o5iqnmoy
8zajkx21aFIjCjb0WCf8z6dPL8tIiV5AjLWbgflHCmMtZk/yf1GKlp9p1ngb3rcy
ZR2Ci6pMh58vC9kgtcX0JyjOChRM7cJ19dBKsbZUPUP8W532q0V2Cx5L2wJBJueg
Juq3rwgu65/quscm3qWClLpMh3MjUcPw8znjm8AeLyGXiBQ2MWqDvJniUYZSBOmn
OAnCEi719pbFBeaaPB6Gg4tYIygrz7EuEja5rcWZmkAdwgSUKOZ8qoxerJaOIcb1
oXMAWZXsGtgNvvyMg6kraibwikdO88wHE/Do4oDMecPw24vYZka6crKZ5MJJrL82
sV5dHQFxqiGdLL199ELDy9RCPNWkCMWatKElD9IsmnEdC69fw4qIBAjFQimgOAaU
oGJWY25FMk9QxWzOf6VrTK21jQkeCQ1fj/fRbYt69BvoQKho+0xVNqrJ++3kHNBg
94Ak51ObBK5SANa3DIDovYL3u1hl3+R2nlWlZen/+QKBh7JKtxPoTLT+HAfJTjzf
uG1SL/tOZKK06ftnpdT4F+WtzB/2b/5G/hEmFuYn8gZ2HAh5a5xDkPIzENg+aLFt
iT3AKrT4ElUi5VYplMySFHaIthfHnL29rXcp84N/gxXqBBQ2uhO9LxfUrIQM1+Up
8wLgTTiIQdRXQuIrqGNIU0H3h3gUmHESmxIcsvy4SbnR1C5mhXIKI1jFGaxCleNc
wLvh9AD52uYrl7qgG9e3JXTuAfOUkm1VTH3uXktDOMCpwwlCV1F2CQ4GzqVSxigM
ZId+OtTJs16+llQqKC6rsNL1rRgPc5A0xPpyVH6Nb369cQ1pJnr0oqA6CBQMlQIz
Y8qkgjoUGryUmMtw1NqTYS4c1Nsm1v8L3O0cst8Puxyk8g0c3Z5+j3Bk1+HLk6hJ
qjN739o/9pUJBijtTx1ZwoVXhwy4TwOif7VO8Y6oMJTh3BErvXS5Lu/vfi0neE1I
Vbt28O7d5BCIOAUOkfqhcKe5t/w/qmyWHvmKWqxSSIge0ggIUBXC43/Hx3GiK/5V
nfF/R0Loz+3CGZPz1AJB8q+Hrpscc8GEIhLUB6mGt36WGxe7XOVcVK5ALvaASczQ
PRvdeWQO7v87KILAFZ7vv0JWOd4GaANyPQGVBk62NXriLeoe74/Iv6e3vlYZxbaA
oi9+2A9pM8N+uJUzvkp/TK9z/KIHZ7GBA95kjOGcKkio1iP1jFUTF1dHOOx+fQj/
pH2jhfc2ag050tqxLRTi7wsvXzQL/IFxWKxW2a9v3JXUfXn56cc9v4RJhb/csHQB
NIdBaBHS63EnnzNbJIHAxVRaN4cqZy4WrL+IDUrCxzzUU3sRKTlUlJloXCQQaGvX
ziY5x8tn/UFQlNv177Zbik6b5at8oORriLTXPZY4JsTetgZwiBuDxfkIwZm+UBQh
5y0ZLo5Cjin7yV4strDiPFx8diM4GmUubGd7sFF59VJCn4g9BLo8yhAXQsNOc0zn
bPDbBiQZgdqplyyyGxHGSC0JqaEeLEe4Ekov5Fv+r1gqy+4Gdz/CFDzPicpW1Rie
erj0uE0g7dpuxI1vLMC/UqU3eFG5c10epzhoKDxYSGLdKYUESeC6YGrxNKxDAuMZ
FxUP4PnFcBc20gJAKsH7wSnlpyuoQc3NToh8gxzP/VaBT43SZH1vIcxqnab9b6Bu
Nac2lHeUOIuPkIbdDJ4QIuk1r8mKSB16aPfflOCE6/wOTXk0s45D+DKaaUA7+43i
mH4pXJvACeVkDqNKxW6eKM3XOiQpqrMp9Cgsq5V4nVaIfA6cgNtHCetOeLkNCUes
unZw+srkOk9A95fTZfGO93npuWCeHjHM11u8FXE1vD3wsIUuzThNYXM9btKXo2nC
FkitiNedSirr0bV3h1aE1GbIDxizHAlsdaXtO/It+cv7l8lRk+Memz4YvrEnJ7r1
P4CZNtQ6vovzklq+l8aYPDZN1aJVS0YViyNTCnSXbsjuMWm7ijlSh+s7ZY3ESL4Z
NRvo0jDZm9AvcbeI7w5J1nt0ioLzRpMbkse0S/SR+T506ABFSuY2B7m3FF20fgS7
xx82+At8N10ag2/7AhlyjiPZr1A4QQHv3InHCmhHF6jkiC9h+Wh8Q038TABFnzZz
nRgEdgjBdfKOwBAI7e+J5FqCccx66gNNJNT3hdfsFDtXsJ1poTUrISEzybRlNxR3
E89LAcRFk2O5XwXu/UyM4+6H01mLsDgrC6twDDg+FwSMIYADmzIg/6++VqmIadsh
x1RoAvgEEb9/Iw3RHDXWTwrKYgyuf8KDzRXn50a4r029EAO9y+SJ8Cio/pjYYMIv
okZQDxM7ONfP3X1G59cS5JeJNYqy2yJc9fw20bqG06GZkbafTYClFaz/KgHZSAHA
vjXBmsvn0UVMyhHVzkWPO/QDQ8emxRvZ1zkDzBIVvgyb8Haz+oLu6kJYo/CfHgnX
k1Ls703dS1WqFgVpDNQ4dduhH/EGbkQyJ4fjGiEr5xc692XKDeh+dAD+Ycc4vSJ9
cwI75Wj6YnE5WC+kgHIfhTYMxvsHwwVavH5t2N41cnk6Uz/IHkn9hZ8DfNTuHt0X
SBp1ooYqS2CIHlUSchEJQv+X6lpryHaT1f05gSby8afx9ILmqCmJyUrXbNHl07uY
Z7+6u8pLS9/ZAiATeF+NRAlSSbA7aZI5GIgTRBDYH6Aix0lhHcL4C6bxBjQxN+Yp
nX30HP9iFbhKnBhxdab+XtF3Hf1BWeKR+wlgpPqrKtyxe3SXPocbXKLuORRhLoDa
upTCkH+4fWPyG3LWFFunGXcR9Wde4o9YqXitM8lXp0D4WqnFkXJT7gxtIp5cFY7Q
HRRNqzp1hQxL5FeQVyBG4SEKqwetie8gXVeRa3C18NHVVk6Gx9dfa1MKIuNp2o1i
Qup2tsx4KRCat7cR1/R+7TCo2bTRv0znhcginVV+6F7z1QqvtupO0AUcYmTgl//s
8OK8iVIZy7zW3hVpr3w66jSL24z0ym7XShMQpnPWEDAsMN307mGg0yDnivHWndfi
Ylyy8rgyMzqZ14fOaTXBOPlXnKPrFZSVUrRo96DTTu+zzsBBL/I/feiCuv0R2z67
oeNz3WcIE6Wk7fR4qcHhhz4tkYG6QW/1nkNbuUdZqix0DREFYosDeWtzP6c0jGas
kZxI3EnEcJ4ePmCu5R83r9vlv7NBgJzNIBwYcW1SvzKiDD3xJdn1C5+n8yMogbDU
NLOQY53d3ZmM7VmvvvVbAg9nnpDeYdoADapAWWmgcyD2rYKpYT9T3jV2q2+m+RFW
cvVVbDKVUUi63+I2S1Ws/fWEr3TSePFFFC1Gt0SYhTM61L8H2Fu2fKyQZGbU5q57
NRqPmfwJdoKB12LoAUktMJAfIGpKWMS4bZyy1eAKLF0iKFupdf7xqdrx+mSJ7gJo
uj1kfe4U3Tib4VNK/DGmhDP4hd2LQXV2gKDYKdwhLUOpuBtygtukY/M46qoXNj9y
Brgjs2H5/SLm1j+7RfslG9T76hBLrYm0rP1SYNQBzpVjAQMX5CWboSR4khrRDVRw
yy6OCbydyOxDpAEYyADRxedEIpk8Y+sx8UDVQBCn5ucVTaW0bEY04dFCDD/lYRGE
jhU61m4oQEvPbbyV4ejdwpY6i61Iv+4GxOZMn/1cmGtddTjIg6gHCZv8WtHjBejw
E1PvXdar4dwIhxMaRtGZRWwnT+f18l0ptPnM/RyEsSq1ckbXG26fhgfrIdj/7pPY
qDZtqTnuuasZtTOUuCRqUyliI7dUKOew/nGh/R3qdpSJokQQ1thSs/w+hFws8eHz
MwegjbLLRkdTZNjWCUuwZ7OBBbui18ZenvZ/un7k7+4he2DGIBGKUn7X4sMbDJ4M
dWmTOGkZxenSl87R0fUzoOTviFkR94rF6falWUpYRcLmZs3TDkl+LmzDlMu5tgp3
uKttu9BQs+1p1OyyLANg/qfDXWolk7BHX+UCR9roqAc9zC7K6HfDKHEvne4tSwjG
sPcyGV/Kz8hPQqNOJ8551zauw0q7DFR/oAaDHMThglEdb+nkJ4rCTX5fOu69hy8H
eZqOGX8UOfCS5cpykxgFBe/zyHG1Z5TGNU6LplaLaIHkNfK3qepMlbElaxEG8fuZ
lgKyzhjpuEKavi8mBLAl+lKzdeZi03nLzVQmPy+p5noVpzXF7rdl1ODeHAtKNarJ
yZDjlM9SdTrzxeOUI40ZEi5CQddTW1jbDFg93B8BB6qYOFYe+2qQDXb9tbbkoVAc
p11Hrs7CtfmIswUNXXONu+Pv7DnRruTaN+BE4NsmSsdZR8uazrk9iS0h/EMehlsm
zT/aO+nFwmP3G67lQYJpIhrU4Ke6lu2stuMf9HCiExCZc7K1WJZ4aP1+sw54+KNr
TyVBdmEp4QvGDVsYV4XJeozJwXQ1ENyWR3CXjdjjzcK/AiqkFWXjkevUXP1lW1/H
rufud4LR8Rk8qmhRYGxz5eWa0wiGH71XvIF/BJOc52PrAnZ9Fonz+hsdbuBJvYQ+
VfrqnuX4VVjSaHcLTyowOoWQ9jcNnH/bM7KGDZCGeXe/0v0kNODfvvrUA5wMrF5d
5s0bZZvbBxM5TNT2K9TpxbPoH+ErIZ8OzOjEfnjYYEIeRSTorMktC3kuvi+wLdcH
kmxKAwhwwcf0Pu771QD7lj6gRy1y2uJPaUO/1Odmo3csxKV6k4FnCWul+Ag6qN6w
OZ/n/sVoBpgkU2JSwcLvNZ7TaehqLa3+jHNs+gTyVB0qFMyBXIX5ZWsPPs7ekPd6
UBMOH1iWL1/N9MO7usVtoh1gR+RxJSudB/+z+yHGDC01cb5Nd2cd3azRAY7n5R3W
U0ip5fGuHNHDygHolRvwMnQeYE/UzcubgiTdv/2/FK2EXP5QK8/F6exIUrfAdppa
Dfj9Vrr7T0k8HDt6bEm2nAoKbY9v/jITNfZVuwlevzIpBYGHm3e8NSVP2DCsFXc2
+84OakMPZW/sJrHbSKVbEyK/q831462uwyYuxczuU04FqfCMMuoql9zbvJVZ/ubr
Fo45jIHckxBI8nRoi18PV1M+NP9TcqckkZHHk0ZTfYWLHjGLkvemz/yUtUJXSUg6
s6SLoJKcd5qNKnv8Bv6T6g1Ba9Na1CYJcCj3re6ytQlQCmwRoV6M3R4LHx3i0+tA
TqJOibglyvB3Gibbi2N7M5LfL1Q4tw9fCWli5vQ5ZqrFVWkAOtqWGOo1bRPfdUOJ
B8fYLJt0XsHT0Jz2Y8PHLTA9KKqe1QzcjuBPj32euyPwt419pRxx1xfOnwR16JaB
yRDHOvN7mgU5h5rtIPo+JxmKFHmotwfxQm9s8LbA3mQj8MXBbH+oSqPN59Vh+G+Q
AfCkUjHR6q5ZDYCvUN2/C/nlq+Eh7CgixsVtVkyiaCQ0gQ2Bc2AkRT4tUB3tdnEJ
+o3Qieoa513RZdGI+NLMmiq56KpqeCQ7yd/sa7LNHWhvIL+VmVfw0Kg7PdZ4gNu/
sYgWJyD3VlaHR5b5MuebvaRrIhPSRYxqx0oTeZEOU2CY4BKFhaYuH+TB2nE4Aqf+
BBRE/V92JCjNIob5XG2Dsqfp2DWsyuIA82Ek3kPhYrtRVCQsTg8tA3euDl2aA5ZU
rG00AM03iTLJuq5u0xiknHR63qUiMa7q4aPFAS+hduXHcWIZKcbXM/54xomU57/z
clJfD9fShnMIO4hHrf64gj2qXtqX/kdOayZCu8Qep+JI6TMaldTU8NJWFuZruNXj
QFdaAfXiozxSy5chpgd9wlaCctd+VVrs+quw8v8SsGEWv5b/0ZEsN+Mb4poUO7Ya
BF5UHXiHbZ5t/lvh3OrTVSegwhRJZPt9EmZhs1zH+GTACXWVimNY4Qtn21qACxPf
1NthFry0qAdb9aQT1+OBYdUuKYsSSuWMViRp6IBXHSvNl98/jFda5EhUzJkUgcvo
rLqyenP5YO5SJOR2n17qbNkKgNUhe4PgYYb0warZtVWFootZu4FlErSP4ncRgbri
JZduQuxsRkZbkrmuibS4F0rpKfzLPNL64oONhz91e79nWvF1HEVuoQX17coXMPn/
OnkdWCUXAPwhke3ie/zxcahKNfkAuxBDOepKPoNOS87UZOgIi0CMb/td+whU+Y8u
qxR3Tkzp2js9R6CrQcTEV6QfNkr7k/A9chAdPxe5g2KK4OHJh3dbpbwCuQo6FV4V
QZKib0JpeutXSJuKwEkN+frJ/nuqzgfZ8ItydMFsLlmqg/SjCjdNVch2Ceb7YdD+
nrZqqfqbk0krD5ywdGOb8ezp7jvz/TlqwzpQSsOUS/Pwd7FzyTXKUAXoxvcYBEX4
za6AilFLCV2qhOc9XPrI35PT2RTEeYIY6DNRH1E4djVEgyUk4D/+d4LaxCWhoN5x
3XwB9B2b3HJZCoWoRZi3LwTI22hDCQ99IAVPIr+XNmKtD8uL8T+MCKWFS6HUMSq6
SCZeZo2XrjrRC7aiLzuhkywXPB622Cius3eNwZ6hTIRjPCU6bQgGv5X850wrpyCd
P5F1j5edzRVP50luvD308gQvBRoKl86t2tx6TvA+iJQ2/aQKDdTAs+4vmlw9ptW1
uxdWql6oAGfPhihfM/5cRWE/RV3/CCiJottW+MbeC6I20pdL/pUT1+HjAB5VE4pH
SArU9M7agsXfxkjEDONm/XDPdN0RKqiYSEKaG9tVUdpprTqJTB6Oh00OkJcd/2jt
OCX0WsBMz0GBkOmw1a1/4SRhjLOKyVVVnhmaOZvZnY1r09Y2RHs3tzZE3bvVx25P
8Gzc8xylvWGHA1pypH1a230JDB+H2YwIXhS/UQdh1z/ifXSiD6a+6e9M2uwh7EjR
4h9VLsOFhQTz0oYzQvvW6HSwAVHZRFbE0Po6CnpEvbGQ2AQLqtkbEX9I8r4Wv0GR
NlouMeESi6o8dZakfiy5Sq/F9ypnMyfFUwvm2C4KvcK/hBiyMqBZ0tiA/8FUadQG
h41NYUeMv498VDfoyspiANYkRHq8K8woR4IHkeGxaoByGKncVP5Jtr23p+DqEWP1
1CPguP6yoxwyLXBpfKufWXDVSXWxPSGkGLy0TFMFzWGYbyoThqXwQopQkkY8AD5/
6j1nT9KWeK+449VSIL6CFYHRWaRIVnl54F+lbaA0rWbw7q0e6yF/VqWOPrhHfc02
hMvd5+7T05Ry5yRlbxJi6lQ1H/Xbj0g/AEpEV/O+J2gWktx6A/Yi+5czzT6lKbIk
/mhvdVhIE5ut2PYfWOjg46ENuu40j2lzi/o8FlEuiARVNrJZOE2fK0ET0Q4caq8f
KwPbVbnUQXA7Sjj5S9IxCBNdO7TSWDdDL3LWTUhuOt6T8NEUxZOtAiTggIJ3FxeJ
z5HZPx1cqFmKYm3ta0msTRzS+x5Ujo3LywPV4fLvq0l/VAYbCj3Hxjs83Gwb6UP7
ycWT52SHohlaCWn1TAsW7Bk76W5J2QgZnGUh6P3euwQ3TdFKaNRW7O7N3tbFSOqV
P1Go/YclYNJ5XYA0+jVTm3fPJXhuI0kn4wShInQbgvMYnCwl2Q5Dyl6MrHndfhV8
dBFm6E6bNYCQTnF2oMq29VI2LXxIQRnFsEhFqQ+7L7w0sPf0QH58+q3meTgZUiEB
xdge1gM/l1PxrvM0W7O5gdLh53/tH/4y5P/g8ORtbVEEBV8UB/FsNzFfIVUJlTOr
clgmdbyXgMtwkrDf+K50wu+3pb7JmbI+WllmdW8ua2JAPkxe0jaSvZEB29I+8Zfe
mCTDtV6v2qO+fCxypgXPdQLTEej6iVNHhakGBe4GMlbQ+CQHgtxNWmKaPrVFiwou
fipMQfJRaxOBGc2AZm+PBtsLvLQ+sGto5TkGZdzDCC15Cipbnc0M6DB76xosN+Dg
eDNU79qglJp9OJX6GSKygHcGkNcvlszdR9MFn9zCEK+49A6EqC9E1a+FJp+q9tBF
yIdfkLGNTS86vcYPbSr3PMPgbTiAHSAMxmVFQ3Ids9jNj7f7AXr+og6wPZ0I10rV
3qnbfbDVhKJOpkPFi+ckEBfKf4UFujixW6EwqgS8HAsfoTw0wJDObalrfZbpFv/W
IjVCa09erm21ObgIWRyk3uD3nYgF3lz8XIpjoDPOV5a8YnSXNQ86u84epQeVAOIs
xkNwv6wQnTcbhZgCYD23ouyWnu9andWU7xfLjI/VrV+XZGmaj5dclvYR+nG5V5Uf
`protect END_PROTECTED
