`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iJvwVQ8FTKIJmRw3SeRRyDyaUxYrHq+A66SLK1gULsIGFSziodaeqDxNU3icYDJ6
aCKKMNDwFyInIcwIlf+8nfHDiBANmbuxKBWqwrT8Rav4gO7JFKly05GWw9V49ACf
ksoZV0/1+di8LttyJ4FZ5wSlfzTmYuteSi6IcTG5EQ2QrnA72f4prrajAhgk/lT2
+i85knhxNiKzc0lqIr69h+Sq43d143EHheMfjKzAQvrkcdEy1nYDyMZm8KgbSuDS
n7cudTQUuxBTwTAPCa1ZrZLtz1NUqbA4HFOSsqnHjL53W21jdnEzG1QkQhpHEl2F
tnY5zfUkzz1cHo+yQJLUoNhV40Mi0aLs/jBlCrqX0yLW3h3yHMTQedo2iw0GeeW/
`protect END_PROTECTED
