`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
xR21zz68GwVjne+kqJvsxjT0ObwYy7WgoQCmG0NwSRK09y1+IDqP5EV+9OIUyhg2
vxozo1XEPnvR13LQA7PGjG4d8VaJ0BTRbG7ZXz2rDUGvK9ex5ayhDH/Y8S2LDti9
HSmvwTUXRxwgzWclkOHElLRt7mkQFW1ujXE0ju4DrVRqXLqnH7tCDJtoQm+Ct5V3
GX1hoTR5PxWx4jSyh7Rwhz0QFM1zHDc8hHrIbEKP/EDfcDqoCfLVtMV43BBloohH
OFgnJAVCyHALp5RZBzooLGvzzkR8jrdAoEW5/jU4tvpiWzNSGMoDkOebioEbQGLy
I0NEvx+C//3ybz/49NGUmsHhXmNfHIjl7/26CrVsdrXRP41IaTP5L8vZqGmCyzoJ
bzfBTjdFcjrcznVPU/ntBlOxuAYVMP+Po6rbUR/1nqgyrXP1dDh9xy5x2w/IPiFo
CAEHimKvs7OppkcuQobIt1xLoN3cs5EuibYTSFerBGoJJD9RHHD5jZKhpM9cz3lJ
3xnuz/OAZqaXP/KQrxuTA+cU6gRPmlXkqhG+CbEXSOC4OU3jriLUBUG0ECnHflmT
Wm2W14dU7UvnavFb+Z0NtYOxj5/YeSCd6G0ho6q2oxRCmebEts/IJLwnpaeqWRFZ
6nzUbkKPDuHBmHjH/YcxPANlqv1yh2HWfGF1LYI3yKHlS/NpS8DJ0GXDAJDMmAdQ
CPGUlwRz0m98VXS7qtmsecpve4dSeFiGDzvInj4GUKKDuT/0PqxJBE4R4syWm0Jp
JMY3eYuOOGbuBkv0z6pOLqQNWPKrICcIQxCldkZXD+y8zt//4W5gH3EBx+U9rwZw
PEN4IeWSqAWe/ejJAxbrlcIuLS91ZxBZiBPFUR7BDzscbb2kxYI+UfI6hXA9EIqS
BO5t1pFB/oCZKr5feT8lzySN/o4e+R3Yv3qpueUBk1EhNccZJOYEr4RHasoVP4JZ
91vvbUMgXLuQZrMsWc5qi4QlyPXpTxqHFvLs99NxQlfkIFRPpDOsF4ahm1eTscAU
SFBY2xllzj+8o39LWauNMVEKT8A/t/KyXM9E7NqmlpVcjbpXdkRN1EelaKhgwv8I
E5y1aAn5HXVIzbIZ/wodi6NMjv5wN/kdnqo1OmPRZGmRpDjjx+1pgbF6KLk+98vW
GQMi4JAV8mn9ciPwuvI0YOhZ+51b7PddoJ6PVRYwqwvlXz/7BqRnsL2xamEiS/V0
f9IYPylGajD5SQAaVn+6BTDLHYrlakGz4tWJhAD5wpUFqaMOGdraq2wBig8HJ1RH
koJtFzLzijHVKvVYt0SubZW0RSow3Yqmpq1jz9dK8WIbv8Ex2FUQyatMj93IAr6Y
tueSgodUu40Odp573VW+V+TJCYIDq0/8se+U55harJa3Svw3FKwu0FOPTTBez8RV
sIAsDEpZWNFje6Tqi8wmVZeV0WZ/cxSQe/sCb4y9iU29H7mq9qV0e0lAlLMAaL7J
Fq8xAaiDPOXuT/ETp1ugUGvw+broK1qj9ONtXX2rKpimXBBfvYPqVDWh5pzzxNXT
3DoapvjyvmfB4n+WiEBVou0WoNlPegGPvZH5Uhlkg3xcF+KbSkblyrd1cdV1Y7o/
Nfzd6TXm2H4GQtXszpVUunh0dVH6AN9AqefhHkXJzrF/8WfrACSWbT3dQ4B9rXtQ
5g0AWBrH6x52iTLub8m0x/RUzD+ASCndloHDpU82n43z71ozIzJuuFBsVF4aDh1v
fug7e0K3wRnv34QWy2yo7lzeiVZGLOow+DZfWgzLvGzGzacaBtszbjyCT7Vl6WXd
s0y+oaTV7bfiAIwuVXiBP0++4TQA2m4sPoVzxEvjBuxzt0wtgdsY/E17tgKBR137
V6ps/ofXb9gu+6uQVd8jF7ElscHAv5/JOTpR0R0PrsnZ4aIAPQkzMlNjK2qveSdc
ECPC4SQStaRuWDZC8k7AwN+SZDpqiucy9myGfp6bEsFNFOQtcbQ3p2d5OjBRBEy8
YEhq59rzaf/i2ba4mTuXU8LoFABisDOZCStxcCDtGNd9/Lix4sToXKNGQu6Zjh2g
pzT1cDn4Yq6ToBW/eBScXlDq2mdLlBiEenVpZTMinbHd2jBok9xoqswzRFdviwzQ
gYImAUK7DB9E6T5/gy9ssczdQPhhUzhz81NLYGG29wF5paJYl1ZL0zCp4ZvGplSm
lk059y8baAeNVwM1j/c4rA+ebmFJPGqdHZnq4DvyiEw2sLYPjpLot/O4t0cdG8T8
g5ld/hN620o+vS/iE3A3i3MX+ICx76kkCbli5/ysLm7ATeI0I6DLFGGjiedXgT6W
5Fmp1QJgNJlFcwa3frSV2V4orQdxPM3ZNF6B2bA3/TpktnNNCCvEoZyY4xZdJhJ/
gq6lCfsDU1UVbh178giFaNdBBi5qI7Mkc/p7KaxHnMYFgdtIgsMHOdnUb4Hz7gM3
h1y1tfToC7cOAXDiS26/+LA9lq5/iithpH/bBubgFoc/VRci7V7ca9ecWj08j4Is
2DLqCOy4LgnVIXfX8BLG7bkjZTCKvvQAi9VE5DDR7riI4wj/FI7PWdpSKOy3I98L
VY5JgEd77Ba60mFQ3aT2QGKY0pIqLwp2aZZm9Ui7sRT23UsENoIRJcx3DfakbiE3
n1Kad6WyhM/Jahe4riwIzV5S9P6jqMnQPgQg2A+2RzVFJ03aPgsJ9VGIj8DofsbC
tNFjSSbjSkmE2yfB2PGwWhxKXUnFXnMHvZohahiBRW0XIR7vZJXSrqt3tLcvaxd+
mb9ri7WMGfKUzRUtCKjjEwIyKhwMh4llDCH/Hs8PYPFIInbF+i8seuF8As+tGOhj
lZ4+uWe4yL7f1gZQW6jsClkJz4fjjpWBi+CnmWMQk99B37BsjFg92kP/dcak4yfq
FMPwt9n137GqaFFnklVFoxZTPLpcmaYraevrHGkRmrzr30kQvBzNEAa8pQU/FDcB
iHNqNUR8rcBHWY1Btr42p/BHS21CHg1YZqfqrq1Yc65CR8ydrcbY9THXKXE+nTlS
/tFgBoRL/eNPuQ9qO5DoAczUpTU1oW4mpkczmfz+57TxSa7jrJlsXXd6mzODHPCz
bVdIx4EhF0p1r2DHUyyiuQfKh4A09TYO06VSg8LAJHSb2xvC/Zca5gi+2iV5Pfh7
AjKSLGBUM2At7ypNwBp69WNEO4Do40midhMsknnbbXFd7sLcSIvqA3ceNeKEX0rx
PnWDW4bIoG0j3Lk2+xS3JRkaKIKUYdv9Imd/LMjcX/U0e8GRE92ewS9szDZ3z7vg
AKklrZmJ1HguDJsD1x+bVRpGWMstjIsYnAo54ePZOtyzJ8T9aCBjVWwfAhlz2XQd
OJliCEEU8W9ne0iFwOh36KOdlw5p/ACUT01CR8kS3WIyWNLJXMwE6lOlg3+BZ2ej
4feP0fsUlZaQBzjke24AXnJgKPJ/PO8P6a7AXl8zndv/JU/Q9iFXSK9A0qIfy1UG
PJ4g061Js5MDsuYet4K0Vd8cyDD4EqYGg22dSCnp60ZEAS8Pol2vEIqIGRGI2gO3
7KoytjJkx/IIOgsgXEZJoVkEPqNtMHzcUg9mdgjVDjQOaz4d2evTtNnIlvBBUDIh
+GUkRo1XGmN831s5B5TqnyoG1cmB2Yyi6mAlK3AJivhM6ic93cKUKCkXgbb4jT26
jjROwqbEH5wmuIhZrmuoaiGQI9r2OEOaD0FFhr+xFTAt11Ek+3Af+sLxOTylOCqA
/lULsXf/0qv6iqSXy0meqLIuQkg2AY21TopAVyH8c4IfOBGI4tW0xoa3xvd3S5rC
bFvRZpB97ZfzbR0YxQX1jzpasuzHvQPy5STPKGyb8wFCVeVe1rzxYAczV4FFFpVR
TPG69/ZWsJv0ft0YVCiISxU/CR6cblXhHVav/BrFzpg5YOcgiQ3jUsuy0C6SCE3p
49yTGvMZ0pQCjF8Bu8oSiaNo86IJsxhxZdq3uh/UA04dLZit0ec0mgk/92pnmVrV
bGrCUHXledJhsdM5FyWVRVo8dXkYPcO0B+3+NaQskkoMwa1ust9jeW+Xgqp/9C3f
lGbAjoR6/biVDcP/RIayayrk7PY/geqvWq+4gJCqpEEwmYlc4Uu7S8hVMOXK9s+e
gcI1MSIIAWyAocPQUec3nBk0wF7B+5y5p59D+ArJLi4GTNCTWxJOOo7F93FUAnFx
SzB8+U2VwtiH8R7FPeBR4QPNL4DZtrmbp/wVvE1Z6Lqopd1yHY8LHMgHYZNjA3qJ
iBZfoPL2ivN67e0g9k854/j5pi0I84NQunhSkrqR+y5w32/f8A1x56I89i0PhEIW
87uG3j25/Q06uyZKeXsdR3iLAnon4jNi/ATDj3VLLTeN4B/jV0TTqEKOWOdDGZHd
8+zapGtwH7KCOVXxlskojOD2wZ6h169wh0u9MJ3QXmVY+pb1FEsz4n008z83b1nf
AdXZHom9R7WVSJ6W0dmGXuM43QOJcN5BzINKEqXYv2YKRUJKGj6u9ycgYhfkdgoP
rBjb4xZekag+TOuZFpPc3E4Hs6tn5lJ+ia2j4SPAU7dPAttMwUYPDDj5oB7eiBoT
FPEvZ4i4l3HbiJmwGOgypZo+tpwv2p94cTfe5njGkGQyL8GJFNXGyLulu/faeawd
mOxLWaGZFU8xRyFADbd/5eYOM6Oq2ek1lGbruQohc2/VsJSLWnDkB9GO0AHYG+1u
1U4XLGCrcNF+rPOStn/BTHdPIt3OeCtjUOzi0T/J138TDSbLsSc8PxxDdTaajn9z
LeqhzvQ9KbYAhcfuGvRH6jWq+nwGeusIvIkCaWkXE8JNc73eTC66zK9r7y0I+JGD
BGPjyS795+fBYo+mj9ivvJASB3dX8gzR7aDYvbLmtoI7GtMsZQEddN5aBUY4kWjk
pxmXt1N9DDnkhNbYt9xSXzeuXVroTiL//IpkGyPol/ZDCQkwtrG8NJQwDlUKiXBx
jXoL7gNDlMGGHcnT74w0MoufuL0GBr/bP6KyvfvVl+wzOE08Kw1/Cuk+gfa1nlHG
y/8kTXIiFU1hMl3iWQ8/MAOe5lfZfo1Z443N5WFeAPFvbNhp5ZbbnDj/NDKXt0r/
X40A2HzH/tDcQmJM/pBB3qBUBxS0GTDQuasJbWgILUbLbaOsPs6hrkr+UuW30AoI
mqQ2MQN8RkVtawZxeH6HUlRQNBYFEaPNB5TLETlf9ls/c+8/WBdo+idd+N8caEC8
TmzG+RZ1mFmTPVq5kpLcLPiaVwGaNLR3MCPZZD0o7+TOU5mLPwmsEUjJGGIDMLiT
ZGLQ8yT8OEVmFxgAfWzEpCQrrJKykpAFuKBGT5Y6+zUQBhinuEoksb7oZTQSzh1M
Z8wgyqGxrTsZQzotJ9wne/pjqbkRwxGcwV4YhcMN6Pps7lIutsOxDH7YdBPC/mWu
D0su6goHI27jScS4aAUShZCobGZ9N3Xfrv6QfKgHpRy7HLtMABof0F6i9oLSyJcB
lh4j9+/W1wcDJRvVL58g9uPkz0wsrB5RcE1IlqK7mssH3y/VwHm6pVzBIFUqrZ63
WebkF61RWBsQcGSX2pHdYY6jsde6HtD6j4mGsFvXlYPNOxibugwEw/GPik4hCKaW
51bDqtBjNYSGGWbg8EgXPduRBXX7bs4HbZAvI535tL0SBeY2FO7KTt/21V6r/4tE
g/WP0sMXPlM6mBEnkAezZls29q6Voo7gh16cAkUivFKyPdWUgNqHcI9P7iA4bhos
OQvNpLQElnhZOuFMM5+bCFdOh3VN7yRl7LxA6Jkxzrn+dbkzCCylEi7NsIbKOVTc
V58RTDHX6tq0cLBuWgw6fEaH1QvCiNJ4nGBt0fB7CeFY9GKl9gNGhoHWpo5DvJEX
KPYXAlmohCO3rv/SRo4TYX9zxLIssptEjrUHUCWCnoHgfuUebG84V7XL36PtowxG
c8xDYdhAqli8MXr+cyzw+fs18ZptaP/ouRg0JX1wVQ5UkSFibvwiPQv+QptxC9Ba
HVMAEHON5+sif5n+KJlkSJXLeCsJ6oM/JfZY6YwNS7r4bDE+4IGfv2Bc8vE1wIf0
ov7KLGiM4XOuX8MBwzsmRW1PlQ8QDYZG0+QUQePAiUcSmIzRYhXZ9EoxCGa+icsO
TwZ19d37AFSsRcbRS899yhhCHl7sF/qJg1ZQ2fO+j0kbeCQtiQc6ZbAxctMg7Z1a
fzEpaw8sEbB92tmxxI3OYRuszKjS0bggccv5Ry5p3zONalnVikcDrI+9TRBO25SV
3x8OAAfUOLUsy7/dCAN+RNQJ4YBZQ2AS79b7etB+ftD030GP1CYDCmfpDWSTPbwX
JNA4vyqEVbobAU/YJqWU4DjCHPXxkr+ijbIZ28x1am1rMdm0M2VdYdTRCm0NPjLc
CefBvgL1Nw/F7ablnMmfx+w4TjudzBwBgwaEyV+181QMWRxGUlMPgp7hEXZcYBgU
YNXYfhTOtHA8utcKvkQzKkV5Enq16EcUVujuk7/uUlTLiJVQ7RKX2YJQ89eGrAk9
5mj3NRvDDf1kf2a3pE/L5pQsDXezg53MC8PMxjVkaUDeT3wPzBp3sv5IE9nRp8o5
Ssv5q+l24V+sNNpgQc/J18DHqcPqwFuBcxz/u/fHqcWDG/mIruqlCbiiSbV5bLfG
PAjSHclfPiNBMCK7tgsWH5z8nG0Fumna9jCrcBMQjuXXFqzl/thKQ71Th8nEEXUE
xxLEBSVzGKnPwWieLuCKfv3cJHCVslO3RrBm3EK3ch0WLIK1u01x1xvevH1p/BT+
fwXr1JF+Ry84mA8eiQek9ctoMzjWnCB1Z2hNmHLBG13ClZtew8X9HHjb4F6h07e3
ntLRfDAwSEIOMYshOwH+t9xtREn9gOwmMPvqXbtBtKWHkyBjASIIVyX9VeaRacZ0
2+OPVdn//f6rLdJHBet5Zd4jYQa/OnOhItSTPbo9+u5qmLkYxpe5K4XK4Ud4ZSTA
6IeQl4NOU19PMHZtIeoBgk3HdMg8EOXTp1bfmuLf+v2n2ZRRpJfxFVdm6qRlchWh
gmEVqBfSoH80i7SdTbxrFLb4RWniH+v4lDfmRewwLVe/QWRAdErcqdecoVs2vZ4I
KVgJSdqlkvxZ/9B+j1hSes1u0ig0PywdOAIZ12zUY2L3cz+v5uTXTjbodT+q7p8P
ZcEb6JXmBHaLU/2fmy6k3V2xl5fiX4wCyu0bmIBbNkM5CYrVBev1K/BDRC7DSr+2
COlR/wi9QGc/ayizshkkqWQuZ0cf91ez7PMigIVxQjPo4ehahWfY3stDpG5ri/f8
Nk07llUQxrlRIX8nWkg86x1FaCpVcuPmKvKuDO12Up4gMb9HUeQCt/or3AtIfyEk
y2ZIL9+7rJWn8bXmRX+TdoDk2Yk3W+35TUOFRJ80y1hT1/tr70/y2IctMIIHDl/t
PTOhSdH5jO023e+q5hco6ycqgxILt/mz2DQZltTGfpMAS0abTB8libTs2F4CeEn3
Iw+1vfpbV2qud4kiXWpxvPyPgkw8nKp3ybvTZJnIZRaIRNqsvrBMcvxl/2qqmHR8
Gg8nqvy9J75w6gbcKiNEI70oBr8Xy0RkExGjbkXKmbMKF2plh4b72kV5x6u5KeVe
kWUaiXjURSXWMxw8SnnIGDZnDcUwSwhI4/OVurK9LGWpw28A8k2AkjGxYm+tgfy6
C/nlcqgTQVM5sskl4mPTpZLy6aGCtG4bguaI8TZbdG4dVtG5sBTUB9WRgjM4QLFJ
8UhCeoJEezF7nLZRglTVbh4emS8t80l8GYsZ7BaUaY0KaVZisqfJwPp/FxFS3RJe
KaVcCzjuK38lWPIRYrBf3756enVdhZJW1LCz8BYSoSk5NWg6O8UUvdFkt3D/fYka
IheWZVKYW4+/BtlGkRBhKZPWV1jcvVwuA1FoIq4AN3B9ylwWDYfySUajZLvnA8qI
fR2AdI2Uiof5w3YcUKO0fml+t8oXvSsAwTAmdlEO/XMJvuccbc+ndgtPnDLGNHq/
Ey1A9DgpyDKW8U1iPFXhPsQss5A+wp+I1YiaACu7s1xbevzz7B9bBIQg9NZq6mrZ
T1gwDRona9aJmxQjIc+FMO1OQiYGt94Df+aduUjbrm2U4LIM5EpVGrOFANAKHOmv
v8h0xCVPH+LseHY7EL+/qL2b4ecuSPDTyqdJBXvKv8vJZIPcindfDxmSaSy1m98A
1SubRiMybf2SCT73Bpa/BZ2WQV4kXJrgl1exKe1O7qXjYaMtq0Pe3I5TlmROAf3G
caO2bC7AUUa4OOEZujweW1maBTYYS5Xg0XfibJrRyHv/t8SLpWDyHp8S/NKKdjQx
iv9NVDUjqCPEOs8rE66pff0zN69EYnSYqSBIhat/O/KG/4S2gFXLDIJd2EfUInVH
6cG5bbNbF3060I6aN71Lq2XrymdXCBUk15utClpUQWirIPOtes4lYpjblDteMxek
ptq2Ep30PedII35F6KJR6/CrEthPBwwNXNP7BPnpZquXYdYwx5imlUTOtduKaHXV
JPl25YGFhV0NGNjOP5N3ysT1WY7jnGSG9nEVltxB0p+3oUQm5BBwT0ylAI2mBP2U
nQIuJAa4oh6TkwMkH/lMhR1CcvZw9fPbV4Oi7LXtx0cugPgAYcL1jMz9Frbuv9Cf
duc5uyYD51sCn3ea6lWTPO2DM9hMCGTOtSF0tbK8pzdUTgL72A9pyZlJ9orL2uJo
rVd/anAJpGQ6qhkWIf8vQaOT1mvjzLYZF0F9QYBQYzSWySFdlqDMAz9XlIQdnhne
OBGrTE6CHhY5lcgbeXSKbjoK/NsEZIJ4Xge/tJuYeylG0m9TY9BRGSQDmRSk2QnG
x4nCsdXF/6c3EzcVlXE8+2/yg4OaQq+PfJx3kvoVQ+ewfUZRZyvorz/g9x0ALzxR
w3sEyLj1W6WQu69wATlfOF5AsPnrn20OQA7aezmElSqr1fwOIM0Y2WP+KqjNP09k
7Cn0bF5v0CDhA3aWEkhy4S7iUAxV3l8vHSAAsOjwGPGhobVU5R3FknWvoH53sFPc
wXi1sTVaFLLo+irspvHnrfvDA2Vd0At3JMYR273c6i0+pBIfI2gDU3Lvw+rtrunh
iZs+I5kZwG/1EEC23n90DtlNdw5LAYwmHqWIwCUsF8JclU8wk9gR58EQYnKiB+/W
o7kzsooh3AH2i8wIP/kdhqx72A9wjF6xZwhI87g3bQPa+KLaKOwzspVy48CmRyzQ
UnOaMCi4Mf2dfUYih4Ir0zT2DW2EJbEEfjSuxkmJZJmNviAH56+InpAH7Ylwk3gd
z5vwsnbf8tfFIN9d3Pd+cWJrVJ2kn3hLMTSw1SmF/3R4fa07Um73SVZCiNz7t2uz
QcE+yWPr1qnJlxYF7bWuWFw22uxEQGQYSiEyu/1OBHEZRX/25ZY0ociPxVXw5Dt7
7qpK8KJkLwuatfC21R0JIdx7RhcKN2IX3m+UmBQAwwipg1QtvL3HTDRloXtp3K58
VVZCshkE0W4Ie3EE+asSLDr+zc6vP08QyIPYCIQUC86UmCh069KdW1Rcv5l+xWPa
nr058XwKbSbNwUuwKoL1itgJXP3iZGW580RPmwXo2EhfW1JKUUIMGCxCk/7Ktt56
kmmZvuM/KPO8GRTm5FP2cx5c3od2ZDloRb202yQYU+Q8Gzjo0Lymt0vnkUshGDbf
tAsbMHk0PINgsCVO1BN2Ecfdc3rrqInIPZGm74BuU/LvgSoA1mZkc8+xYTnSA4GI
WCEqJVTCwxwIVwlGNrrGXu3teaH02uN5IOeL7KuIRhRRojyXjNnXHAhbBvnUdJZV
rQStPlGkTT3R4FSY6mrVj25rhdFt4nXwxiE1BuJIxbIMjr+pmnXTKwaB9G0y7sHj
FepS4RyVTyRbTa46dDHl85WmZxsVuORjBuBbpMsnqbBSu9jlOtBBYwixiGJPEB5N
YO2HLud+5o2dkI55ll0RxUp+xQcQB5xh5eDRv+YfSIwUNi8AE9tMeuKkTOtepuKy
Q5MAmSMDTLEHYevxulwc8oKYCfjU2msU4zgZ+RHPnDc+c0SQjqrM8CIFit6keqMF
/EcvBmIZ+IJeuso35Fl96rJsTgG2A//og1GrvSW3rG2upfb45UxQPiLLyng/1O6a
oC8HQEG2CpIkQzccIsAVoxPbuyQ05kS/drOocJFsCD3sUV8/b1G9UZXyTktZawpU
/N3wykicZ9GA7O5WRTGyx8G7jCWYrzn87cmy2Bp1m9DCggVtGWMsbBgBygEZe0tQ
CQ2mWQdg2zKlgTysfT0Tx7t2IGWYq97iyTvBcrbExJhA2N41ojAG+My6trk42mUr
AG96GaNDh86Gr4B6bE2x26L/B2ISgw36VBLzk22e6/tXHTu1kkWdH1gkMXfBV8wA
POHkXdpV4+IPFW9cOhfETiX7DB6oHGYaT4Loys5463Sjaftw4TBMELO36xTN67Ks
Cfu1kItcf5I7OURi6J1ZItru+zkQRlr0P6cqC1DNmkOC9iGF4qS/qcGyyiouT1a8
6xFD+gat1qWv7q8Se2ECO+GyITOklPXyNzER5aDuJM0Js4nnC5d75OroVEVSuJAP
dd8aGJineKaqwuiraO6OlfZG7eo4KGz5NRFb6VUvmzniSAAznggL46hie0sG1ytE
8swETgfzb+0nYiPnFCVwOJJI6Ig+W2KMlhaQoAFOoYphgrMG/v4fjSbcrx0VrmDe
Lg0aDWyRqwPQXY6eDN7vnxNc7c0zqYnOyEwMpdvrxkw2ayAftnXGue3fzhFVP3d3
ssqork6/P2VHyeGvn0Mk6sf3K6aaVmdpH8UZMBroDxUIT7AlgCOnlaZuI70f18Iq
KUDkZrJS3ZnlR89mkzk7Suw2WiMoexptz2Bq2H2RBrF9P3ag3v4Hm/geNskgZgZ+
gxKZt2kUTQFfocCUZApDoPyVgjZXFzr2KdYrJo0VXL++UZsF1v7aBMyMyk1malv2
ZD4J8vsCUvKI5WwmtBM3I7KvYxKaQXeT8B6TFVhwLbP9sDSsY6wFBOuR4nJ9Je23
cQ1Uq2pnjw44wm9JPH2tf/S6kWq0rb5NjQ4iCB1xU4ENmSIGW6iLoFh40CaZIeGh
8YytRDzaNAu6j+VNYROUCSSxHOEtwjJX3iHzIdZWYBlmrB2QyS+RmkAxLL2En6Pl
rQSEIfH7TDTBJO4RpWyrBR7G8gr9an7A5wD1Cb2oRI7fBU/FBQkdey/elOJDBD19
nFrSZ4X3MZ5trxi2ZnhjhZLTA5r3euWV9GFWVpF6WeFjDqg5CjmRDA+9uk/q7Xu+
cqV9dMNAi20ZfZI5W+zx3XVQPdlfd/u5ftIi/XMZ6OfbgCFnjU2fdz0iGdwszA7I
sJvOptnOyLbnDpWoFnhN+TQhZg0SJR+99qKKBzTOM4Y/QYNYjFA1YJjqmbIpRTjx
D1wjqN1D2C13Shz+IlQZJzSRHk/P+mj69VIL5zUi87J452SxDnbSFsqZWA4IaKda
t5qMqDGF9aftdYxLMBWXqd+O7TZr16CAHSLRsRY+cX+2znDRbqvx/SQZe/6SzQST
NrR3MsqoYboQ6xmjHq7p2dcvo2ix/Mp8jw+Ss57cHyKRcBuCJNyi1JVCEU0PVdiQ
+d2dCK/qtlwIprwrp3RH0yTCICTFCxUaqbRpGMHAlYmJgccXEt30iRDYL+7OpZHS
IVIUNFwhX6EcLTGs5bIgKOK+HurydYmPXz7mvfPPsgt/peLzMSluBZ5h2l3EFSd6
vgxXaR6AAA6K8y8961nQlvJH3pq9ij5yDpRtChI/kMFTegVjPhX6bWfHwRCUdU4n
XFWHN4nxQZqQJ5JIS7icAkWDN0UuNGkQzkMIsyBgffr89IHPd2Dw/+YZqq7MNrU3
Dd6CHElM4199cl0YZsoUSzv2J+7U4dHZmlaDfamuDZygjcDeTGrcCmk5SONHMBT8
c0MtLjtmjZecKZCMJOSe9++48oAZGJtOsw59WolDuBVMFftGM7c6j+QO1G9Y/tC5
SZ4oleBVhSJZRwD5Rbl3G9ngHUDz8nvzs2N3rmCOmLoQ3K0Ev2YbMClZEIJ4dStg
/GoLbikyB0NHz41pXMsZWGGLkZFCJshQhxoE0QyYgCFDuk9dwR9g2cBcTgYoI+UC
kSLZNmx7O7Ey9lohmCxaePRHpaSkTDtbIYXVelFNv4HGnvOMDefaXbCKl/UxZiFu
RN9pGVYvCz4AXezbb7nL59AMFJp7i8jETX2a2ALp9T8OR7V3h8oB+mrUe+AGC3Th
h8aatu5ELX9RVXHH3DsOBUFVSqK48XKivNEgLBNK8RPrhtyQZyAsbQ0Rp/hxoGkA
6UtZWkxIYZogsy1hNv9Epbp4GhSDInq7XBeveDfDQaQ6mvBkJOTenKWjyTv3QaHU
WaOdZyvw8hY34PkCwVrMDNviv4dWq/ctsNU0SOcLzBOVprsUpWR9z12PhZAnyp1V
YSTzjr2KmWpgUgensRs2txtAqYHDAfCFqPo2lnh+sUqq4jQE/nGdu1H5HXpxCaf9
bZcx+XSdtdd6p14TiuwLhLps1QTSbQuWq0Fx6ZkJXuY4GvvAOujw2BeYNTFY0Ile
E5cU6w2eEGHgoLkmGe5ugUkdUFa/TU1Vkab9iqyGhqUXLGd5F8QNQNIYcBR/JWB2
UJCuUGzNkK5e1zwPNJVqw6tJsC4zFnjYvWYGAYft87XJAYJmdzxk4SgncdhwbZ2e
Yqq/U8tOMVy7Kcu7sJMu4VP5dKJ1e1RnX1BmloaN+IK8FcW6b/D1RcTRXnKQGWVN
mWOFFk8xWPRWpc+oG2zlMuj1+i2SG2ccnXtZJtp8fagSNGU197xZHQAIaDIZn2dZ
4xAutI4jINj6owiZ39GepC5mUak1/YFaQHVKRptYh6nPtVxVdjX51+YDkfVh8L8U
VYcXOn0KantAbhnO4XgOCUMQBHAgWZ1u8qKOknQP5kVxyMXU+tIA1oLNBNusldUA
98Z+q8tQb9y5dZZnggy2GTCmM6SJycbwZvxUC9IOosNHuaQgceSJI7CLFaqnE3oo
29jR6WQz5sZHwU6wVCxY/0bxMCKt0hYO9vo6NaVvYoZ1LmxEPG601SWaMd524gul
YZBaYvATBCQdWulBCmL/gk12+2NuruJl4TNWb+IBcm9NmaeGc4CvXQd0sJ2tj+KJ
fb+oCUjJe4H5Q37NTQQ0j0NFQU218mySHWF7fUvDEaTAjv52MfDeIbV2Qly8FP/m
bo3jFQe1TIpuO13fAvTM5Qb2xwB5wgyFqkaaQySBrNbmhy+j5rTf3y8SjY0hU/JX
9PDWL7Bvv574akvrDVE6Nm15Yw2ex+zsBH+cO0lGUhjNccQy8r9pmHj+PHjKe1YK
XJ/EYh/5vg8wvGDj7iHGdrWOL3JO+Jw5QLGQQC/rUWIS7Mkwyju/zKS7DGYNkSel
I03N3OT5aHxzClDsNu1nQzgmSCxoiQq8PkQ+WOCd/lBFvxqP5ned2PmkuuWl6Ggd
5jBeSknz0JQFAls7+XmKR1pFdoaga1wQyqSm307etZaybZLWAd5GPWKjqXT7Pegz
fYlzmvtP3iMQsFrpCj04779zmiyNPEIM1Pfue7+9LGL9wzEhyJru+uMHCvIV6kKL
OmJDRclLqEWBdR7f7wvTJ9P5WPUBTfbEgH/4Fy+ZTAeJb1M6Og4gu2DAlNPWJ0E+
WiTSQz2ve5z4wGgm/ql91VB7x+SMpJ0aK1o+VJYcuXNp0zM4D5NWJ0XlbTSIUhE+
rifHlTSpvapbd8KpssLRh4rB0SmdayZOoALXJAORi+x1SlXQTeAF/plib0ahwaGv
RtvjvfiLLOMwS2iwIqfSf7BTcFC6Qn0VcklTKC/PmNAxQ8EOqkgz7O0+S/8OCJJK
uQ1AOJAa8yentlXBOmJVQ8e6v8wYHltDrpbC1uoC9pQNMQ6TogZ4zaOzTBWX5I7B
VRnsfXMP6nrj9sWI4zWql9pKcH3JDa/7YJHAX5dmOEtzuvZT49UiDs33XpSPO0TZ
jonYmh2pc4ZbfWB9IItFL3cYfNhbwLnqAZKXtGCU+XQBNrCszkKxglyw2g8Pauza
ArcZfWqTxOPC/t5jVohUybIl04KaeTh2kR8lJ9Bi8GnhgUMk50g2d6c6woGfdkT1
LPty0xpFmESgI5lgWBKCdCqR7tkldXUW1w6y+oC7G0CcH8ts/QDYoiCkE4SArvh4
pY+8cF+STVjLxHK55gazLB6b8gxlGS1viC+iv9NFIE4PP2YtzC14O4j06YypKfTa
DG8Dpzk3iHUA9Is+beQLPogxNogn/B/O2bH7CZMHqsf/B2lSQnXUFRaejevbnW90
JTOXXahHjOSw2ZwxatIGoHWmC4elc6CTTuHRTHwvCXlzUHoxC1g9v7Wnvg3IptY8
vIWlLcrUuxL2FFykYwT/w6OsqvZTkG4KZpugt10CV1tFSlyVYkysCajakRN9iYo+
ZYaL+Bk9U54zuBIRoIDDdw+cvQSicnNG4jTMRmxalg4rISoDEKfH0uh9izalNdFN
2EzNchLF9fBJphlk00hoLjngZTe8ymwrk4WNtUSUW9MMdTKVm3NmOGLzAdtd/1ek
xm8nfbNLBrB/Pabcqeazr4kc43B2gPOlVqrtRHlwLOq8Ibpx5yF3Q/nZZx6orPgX
GoWfNFSNABdX40kp2JAwbkdJBNCtoU1rPBGqTltdIKcmhydZYq4DX9TvrGqc7rAJ
NFidzqhQufehPIoBeNPqSv4RVJwmFrtATY0ny167qqHLLSTFI0hS9tpHtaBm+XPQ
tlUe0sIUu/gLOPyaRboJJJhdlpGN6er5JJz11fgGOLVhbIghRgqVJGj2yk2CWXmJ
SBEj88s/YRhjvWwuama0HKoLDJh7qno5Rawy4jK207SsgNhwPjW+B0wmz/tjcqCi
jCTMNEAkfxNx5N6sWAM9LBRwbLf8ApRSti5qg7v+GVec0XkN1nNGbMY0NrIz8qFf
17WBTbKrDYh9eXq6QNYXTB0LSVEArs8BJJ9vZwP9SS3K/6VDtY5MU0X382YK6NNE
IhmhN3z81XHegt9Ej1Fb6DX3v25UJSXjmDTjmEXJ7tELCtCHOyaCNU5bg5joP1Jt
p2LsSQ3dn+984zZoCxmTY2ROpyWYWLiR3Ygxlirb6EJ+6RFRatTwrB3At17ffw1E
ONPwy6ZQuTbhlZgk7IMUlIeMEZdxKaWfdJa4REHFRhYtHWuOVvsHzn2UcRi5QfrD
dmqiGFG7s2DQ1za9phg0HTY6OG66uKLsd6m9nRtnYEBjZYSjILHcnLxcTP3koBjk
f3mXQgh6NTt9iNT/mhwxabamg3/sGOMZL9yJzlF51LiGZ4lVz2yzR5F6xfmhpb4w
0F4lw+ZiMyf+AQ0DsRy5uvpyafaLRz5nwn358zfdspoyDE6KXX82h7pX/Q6TLqnC
c1kJCrzponBN7EHFoqx0n//6gaVDHlj9VyQm+SNdf1U+AOyS0USqu9hfbQZzNRJ/
yuRohKkcDd1LGVlurXw8TU9rzJTLozAyZm2OrQmgo4gXPJj7hgKBSNQQCauXWZ9U
1xoYe9h4sCHi4FxJ1GZWMDhL2VsDLy+NJzPRT1rjuTXDhE/Z8Wvt4UEEbFJ4ibQs
PuKOHMTuy6uZ52iAarg9OgdfwH9tFzRF00QA4bqci8d90mnyt75TpuYKbIkzS8ox
Hfq6bGdRwJrBceP6g0VEx7xaP3okfOPaN9Etj0CgIQtiXMQwswIfj4Qv/UkYSC5Q
d6HlGigGOTXyY3U0P/32qD1sfctOpnHniuh1gKIxcO9zWlSc+IFtwmaENDo3WM0x
WBcgW7ceaddpSvXM3Xa+8lybVnYmIV7ERnuDnHxsdD2uzHy5C52YEHesVUgEfcnD
CoXXAGCTtoaheQNfXnWvmCKezLC/HAbop+j8o+BtwfnjvK82CWwU88r8YtSJEIE2
2ddLJOHXBSoN3xmmlz7yGcqgIIj8dG5GsaifTogZOTwUJ4nVOygN43Oss8rhfIRN
egsjX5hvH/GOrsqqJ2bXg+7J0CuUt9i57aYW7tWAb2JC+Z6I4LRAGW9WyGc5URLz
+/rCHQeaK0YgZSTJ5sQ8etAdfLhs0BkKL+ARSLTeVrPeuk3TiYjm9fMfTgZmliNL
qU8t4D3ejUWn7rze0yIxXJqcP0DdVQhnMQ1PL310b1pyAB9fjNMHjrGTr4AVHBHG
azOlYZ5/PjTosMor0Z5e/j8jvka/wpqZunuOWBFaIQYkiCe659cJ0a40GdiEKfgd
1FRv41vzxQr/Xp7rLYxCPUSlBbNwn6r5sg0xhe0sNVbD+4d8rzbtqdReHE3HBti2
al9pIjBHKUo+z4giqMZoyN2w8b/xgsrL4QLY69I1feDRbTQKHDhG+C05ivNGyhEL
Beb1kukTTk52Gaulgg1fcN0877TbGsy+hcvg9HihHsqJX78BzQekzXmveDVC5Edc
qUmNpGv2Gu2oZFePdk7TVdqqTm8gTh+tmep5ulMn6M/9em/XA5OjiQAxN0Ld1D67
Mq959cnKqcKwlRDMvSdxcis+quYjRyl2R9LxsOCz0R0LoDxNS59+8GJ/vbpgDx9X
4AtPN+VV4JrjpLlQxd9J9OPNM2w2AZ6TPBi5fZvTLmNGM20hBhwKYxmqDPabv0xd
b21lgxd0xo31sY75WLb5JnTMYinpDLSG8v1q4Z0yzjqqZtdT/W2VIBzNJ3wtgFtJ
OdzsLA1Fqzl9Z1W4dqAWKudAL6guuIbmwhesJXOA7WjGtiE2bs9kRLPujBFgaHAq
gU/k9vv1fsWbAq+1xjJ1qmAQsEmlUo9wNhSNgPONyevIQcA8sDTftyh66oEfyQpl
WhQqrbVRU66yYxg/ekhjO88+B440pgW1Jpis57XsLItXdn2iGtUyhNw+QmoLACM+
S9RQ3RAm5FxWf4+GIBgj46zPqcF1hl0pAWcCjL/hfGF04lR/c7Sza/DDPt12zgNh
Cwv2hovDDOGWSI1+Ab1ZgHTThnOBzrCwDaWd/tQ2QhvlYVqswqoXf1pdPX6zZM1z
0I29nwAdKrLNmK5c9i4buH1y/D4DhfgJkHpvDLpQRBPOdbYKxErOLbapy9UwxjrB
HDXiH1thKYqPaoDTszFFVWMC9qIQR3osvVVW3+Bg+wmcls/IOTOC1S8deMoawYFc
2PHcqnbZS0h6B/6jxWJ8mj9tZwi/tslmQ4Ktl33R8/EZnhuzciVinhR+6eXFCLlk
sD9P0cLu4JsTzvJywwOlbOG+f3BUKtV+iUngDJE3zgCRrqG+o9CWLV58BPOMmsQ5
bg9i12uAtlXJdxFkKHIJjWtmTaaywGYB1vEjWelqYsVyKjVIJF8YxG35SYJyPXSl
ARhR1vkx5UEIWYyBnlxeQwPbIKAb1cBSlSNbUIHjl2FomWimMYsIf/dPy/tP6AGJ
T/825+edmOBz0FP8Veg1Jf2IaaVqZUTMg35xZ2rxxw+EvFfgWCCVyWDAO84E6LOC
DdfN4fslGJQ8eqtqAYIRR5D16aAi5cOcnm5125P5pFHNIWNpWVBG5yxBl9QYEVsO
rmb4K38pKQD8eY6x4nBNKCXw6gqDLQtbx9cNF9ZRn/HeBZ2gJPnYWjmJy1+XPpOw
Q2H6U88SwnTaKr3W5cjnqZtHdGye+mRIWrEKD4ZmIwGwQp+dqp/rca4RlGxpaBfx
tzqmXfJGlGPrY3kAHUuSnODvpT3UP/9uZIjegd1yYFLxx0DRnLyvbWts7JdR9cwi
PNi4e0CZYfrB0dgfIFgOp9RDnGm6yDbQ8TLJnREtopojZ5Sf2LShW4R7BEfvmY2h
FzN8eM6EhMhOhmFStZBQ4iE3ovW6hx+t2WatikhSCnfIlVF1BnCPtf5R7lyStlLH
5QderJehcqZSyxCOmuMiPEimqiKAzhO3lBcWfCVF2AuCH3cp6YY/iUQB8l670HTZ
hXnObGsXfkOqZicRtXS4YY23eXRno0bHlsnQrmeCrPxJJCigKPzm4+s26ZCrWtj+
fXJl728PspF7AYQgX8/+T7n5Mzjo0myf/bKc5oLxUu9gHqcIliUDsw14fINqAfHE
imf0c741cZw2aLyH/Lr/pO0JioSNpnNBhz09tNkFKROsTfWLYBZ5dQkA7v8Gb9E+
jpY25HuVvJjlolnrLL9jGw5urtCD7Vfdx4scOvL48fgU5PrsUGrjA5iuE0XVEm8+
lb+/Bq1iG9FX/G0woIDUQE/y8nbtcle2TZixMtZVcRYftVhl41rMNMmm4ekIvl84
EZ8UGodr86WS0LHvpg8AyvJiWxF/HCjVr1iEhNomMH8rJBlCug8SoU/R1RdbWP0X
oeASwtk8c2ILoZT3x+PSqUpSB7GF0tcOPA3BoBki0JY7LhBVmf4A9AX9mUCoM31J
n3dbDY2yF6GSslpJYzL8ujJshmMtbSJrbsmT81jOvM//K8RNzX2+XiPn9oMDHkZ3
jCUP4bydX82+Puafo/dW+1pCZnCXwTJ8UR9O0oqVjiCA4jtVRZM8fMBdS4CD7L18
6QNJDOm7Msl5UYm9Nh0o0eJS6SCNkViU0+eWqFzbvusiKQwW4u2Li6hQZ3lMRAM4
70FwHIsI12Owx5R97OwboLyKAVD5BOlnxaoaNnTnajH4iVLSGlEaxGWvsdIUGFFe
g6ixvu2thO9MN3A9p+zvDoTSN4AYadachUjMOrS8izohuNHj/T9kAKqn4lYnmm9f
hS+s/C4XpB6Cxn8QzGRrtE86qIX2lxHt/ebm/68XhU8bMiVzZmr9crfsX3YTdLGK
5/ZdFUkbgrzI01f+fTKEM5rc7tHEcFKRzoIa5FR1UWdacnR5xzi7BI2flZzvx81B
26IqkhEJmRs+71Fy5mGclnUK+6OKqskncq1wMNfIt1dkR6foBUxAoMsF1BAYQdho
1FdNhd8pbB/nWdafA6LuySKiM5kGEX2Y8rjvqLKQTM8Q4IjEdvnvLGeGXxsYO+0p
OuUZ7kjsevnuPkG0i3lyfaEZ9T1SrFZoVTYOaFUMEdmcAjrpdsHmkpYqBIQLh7NV
4IJ+fzW+QutzwgaBjusXhccnpARHwAfl/Y+TMqowv72DOxYGtjlkKSKgdObrSacm
DekE9ROCvCjWuA+TL09a5wiAPBp3JRWiybLibit72D8SSyMKt4VLiHzCmhu89A1Y
7ViUgXtmPHLE1EU9LwGSanRDMu8Im0OmwktzoYxi5wqZBW8+PydOMFxcBio1ovUo
LpCCQiZAO0X6H4KgCQpSlAbwB9DbSFZRmhu4tkEXjCGNMMGbuzkKWkDtp0uMDfJa
fUGwGCru9uU8JWlP1Jnru5yxMzjFD6pDNS2/9AG0PCmPn1JdRCPSsNPEU66jlCG0
IMKnV7/4z4LmwfapTm6rQ4aI0Ye6y5iWg87rtCM6RtPBd2l5I6GHIpvp46F2DYXL
TBhvBG0ILhd+oqClrUNfjKa7R4OOoljSPTq+SDaNNX2EL9Kzm5QqDywqpLGD31nf
7ihO2b043VD14berM4hFRY7eIU7RIl41kz3huPrKtpuSAR2/0A45cJnYq2xvlX8j
Vd1Xnr7uyKw9NPZ36+ojKNlaHe9Ap+tJ3WpLAAw5wjEz4Kw+MM22D8+7vbimsHdZ
RNqM71239xDSrVmuR1zCt08fPbFhJN4r0yWdfKLfMtlzoulgqLvJT67lAZP9uR2Z
ikMwcBsTdcIsZqJAmHM3tNCPJrEPBwlPlSsx7JL5dkVLAD9WPodpQQXzGEj5taG4
YOCOd9CnnYTvxQ0Fwa/62nV8XDCRd/xTLEv9HHjBI5RBv3GwHzXR4xDVBVYS8A9P
KgZ+r/cJnkFm+ISa7t3UB47A5O9qQFwksFgY3vhu8AoaZsMq07sO4x03N64iN0tD
nErRiivbRnvR4sLX+u/3s+FpSwNuBd56sv4WTv75p2w6GfqGZHO9AfeFkhDat10s
gdJhzvSO7QpDD5CWnLSc0at6NWtI4OcxMQFiq6Qd84UocIp4uEiggAak1SHJz8iU
lNnPKlQhnOd7siNK02ZtX1YhVSnJ3ELKP60IhS+Io9Z8xXFNUzWEZFFyrAGA/TOV
+pTqyk/dOHrhtEvKJJRAtFtnd285p9dbkq0jAqbWSxUJI/oJJCR4trAqHyTOG+aD
9XyZRBm0TIFZDRZVLzWhOTXlDMBSYBg6OuxaY6efJfM7XnMPSKImJAieGjj0B4o5
LYWx06EOAKgFWihZpLr5eXc0K1t2kqJimbiF2NSnL/FM6bETHItKtZs19dP1F2Re
LRJXlijSWKUonxdTYEUmgWF4hPSmcwdOBIQkhaKeNLEh6aIW1dWM6O4J1DnSCQjr
A7JdrDJ1y8XI35/9ooBZmzXIrggjeIhJo/m2/yY1hnzsRabK/mj1WRwvyW28K0ZA
URQcYRVqrxD7DBuaouYOcOvwFfiSYE4yEDm2PjOjqib1LkA6V4ZEjriqAREqscpW
eF03aXxKpo230JdzZNtPQsU3wBK9tzN98L7IDg2KkKlAbIE9jWX2Xuwnl1Cw8J/j
jiwD+gVhlyFdg5sw+omUSvEERSWxJwa2vQcoNh7v0hz/K1Sc//qr9K2wxKIsFnLG
u5AVp6GHYtm2MCoM36svJJ2nB3P0sk6/tLHdi+dDPmn0XZaNUCKj/cr0LGLrBMS7
TSCC38iRGFB2hMwHhsxUEKmjX2pxXluJdAZCvzuwXu2bL5oiAKYc16PmLq1mf5vc
Z7UXvcRNH21+viFjJIhX9D65WpsGY12/6J4BrW0Fujm87iPzoUhXlGNJ+xOmmYHD
fTqK5CQtJs/QnMj6ueLWp9RSSGA9QmcKIHDKgn8g5vQ6ZA0tMzNx52sF3suYsKk6
csmz8EUIWgpmWeX9ovk6pRNO5aIFR0z6/fpAYrmyY4xr1gJ9tIPenUEwvrmPcdu6
AGAPfzo/ut5umILn6nt+oG9gfg8+3ukxq4EtALq0woLrED+1zXGFlxlg3v8SBrU3
ZrneEJpkKlBduxcFhmJj49suwIqLzF6OSevPh7V65VjgURsXdInludrRvz1uZKzx
yfRAJS9yRQCCRyvromi+JtA5s9i9qdawoIknm6G4f03XLX3J9jxXutlD6NT4otUF
gKxEq5rIlZtEKbMJSQN+o8WvxdL3GmM3hAJCWRBraVR0rMsUTnB1b7AGeIH9r9x8
2V7gbdE6VYiAyDxarwzmO8KV34ozXLtPjoxORa8tZMz7oVZHmOCyinl2J0qXAKqz
9qF+ifb/eol5OmNCKel8xT8gYlS1JVJKRS6bPySY/TnX4hgR6MAqbQIuNTNzwtfy
gSqQVyySmkStQ7y7Ccvdyta7W5lx9Cig+ObtqkbIeo6Mh2fRDJyN5Z/+Hes7A41G
W4wfcu/ZwuBmL8ycZWgE9a/J7JLvxQMFd5Ef2PdHJWXZRArZPALUk2Ucl5lfAfbk
WOiy/7GSG3AXvQ0St6CRxtgzlSee2M2aWC4XSToGjVCm3m4fAqK1hG4+IOYfqZgL
Yrrs8knj9HREisWLseGLsgKO7XmnxRy9od7aYRaezfg+SASVQVKuoNaFsOB1V4Sv
OhlB06yiFH1S2ydqvgsxmIpYgab5n4niaSqtKAG42w1RgE37Q8/YuH9zVPwMfgZA
gJ0ffXcPUoJccY/lQ2wJgaIQiC0wjFJESzeJrwDoE6IhyCiPRGhCZHAIcbZpe988
WL35Hq6cukAIuju/6p1E8CjLJWjoPqQky9rgZAnYuvdFAwR1eqWESSOHpFdnx8OX
f8RjhP+8F8MIRMFTR4qZQ+qILRMcWmnoyw71wPA0HmoRt7zR5EERaEU7iiphg9/f
lbHs2dfLs1hrlJhe/mxGDIUIgT/7MM6DZlDXfjLCATjl7FwaofMwCKQNXzdhz7X2
UzWISiwRcScEaQimVws5XKm2XeOzKIHHV+ZxqhRiW2xQT51CpegELcw+g0WPYd/y
QYxmgxxtKiUg4DSXFquSVP1ugJSKnptechryEZilbqy1ceE0y7u60cF56nOcddX7
ZTzhJDlz8Cx+1YXy4DnszvL2wAiE2lepiw2vh1txP045eNo/Mh9J5ZzS93uZCJm6
DQJCTsHps2687ZZIxBWoFaOzTcIeYsYsZobQXyFqRKKeydXwCwVUahynoD2vBnvZ
emrI+4/F2t5j7DV8mFh5nqUedSzVbvqjXjXXCyphekcAIk5jH/FpMCl1zEB1GLL1
hcWzMWWQRE7AGdJJh9PbHPPSA97r+m/wLGeQ6lfynA/027ERSMEfRQEMNHI3zkd6
Njur7JmZuE4ZqIk0YDPWaNGRhDQiAG/kkM2aL27KbnheZ1+DZF287C2YhnthfdKB
oy4hQ3WB3hw663VAYWL5hNDgl/he2DT5vRTaImsgX0ZUYem1hIUSYWo8YKxikyB4
l3+6uBqewt7E1rC8A653UDmGjeQbM6s8/PR735jRC9wgkgGtI8WVU3HuOC2ShW7i
z6Smo4Ii8RGX4yGzdoMpe/RTnPqUVIFRDqS1PmI5E5EklTo8GbnJDx0C5/eT5hwn
yOBXJd3zKGHLNde6oUPpHzrvdv6jiRyP8yVJcIIlMJZaDU5tYUKxugTDx3G8WtDn
PoScUO7hlHq8Rb696mXkciz94y6i2upptuyLdfsCEXNPXgdHn9YFenksGpBPdU8Z
E4VJOmp/+Ud8lX3wucqmQN6eCRMoSaKSdqjhosRbV2uW1RJXJyeZ8uIGiYna7i6W
rv4S/gVI2HG8VgcatnW+iH1I+m/l53LnP6vDu3yUetEEBK+CahDhvtDQNCUwIuqz
PyLY7RwDvJIS4kQhp5/IHVEkAUTUBt7SCwmmZO0kqyQo7hTAiF7TU6d3ih6pjEdq
H6KKngkOazOaw7SnZO1RpSfdIknY5r7xeGIun64FfjGWQtyeGJYcknrylF29cJGK
7GmI67ikyBkIJLUnX2iCBv8Nxaljy3H5Mx1MHwhRQE7fos7CurqHl6IDiCxkUOoz
u1J11Y/gVN/Kco2zXySbw8w5UF+FR+gLOXk4e6Sk9TpLiDNHCj8mkAxwEkVIPJ2X
EKIvORkaHd6GdlFbmY68ETKA5sv5bv0OT0bqK4BxaiQbiPRv5pUx7cXLMb7jaa4B
cJdOOxG+Xc1HM2DprxvXsmR0Jd4vT9hlxZr+tENfZ46ZVrYXUUqoDA5+s7rh5Bv+
KZLwpsh4YyH9V0L+l8SS8xMpLvl5ZxUc8HpS9MSVTKFyKuHNnxUJkVVTHgTpM3la
461o74XYRfSh8Co2O/WrzrDOycQ0iUWJX7a/K9JTJjLX515NYCxA8DXAmoYRBc5P
tXurnA8u7L8Nv0RBnhE7gKzNk+HxdxxTro7exnVBikq+iXZ5VL32wfPUJ2MeStn3
gSC2ftNGgCkhVUA24e8rQwdGUhVsIC4567ztD/eFJGNMeOxDj99EGMq8X+JS6rOu
ox/bYhY0HO7QuyGNsNl9GlqQ4f5rebSUlO7lwwOkOvxsZ+dynKCrRI5bCkGetLSU
6j1oELLA8BXd+IbvalCz66GfkLYzcESfekg1doKCKP/SQxzqJAxTvX5CyEDiK6Dj
XyQTnppo4GOFX2oc5oKzdQx5t29KrrJ13juRAl0z7StUrCQKgbPXVxidW9NyZOu5
1urL9oG4FTZCUHYmTm66MQ3XNlWTdGttVKCQXKmY8EDaYU8i5E+V7lxy/0BSYfNN
S7q4b9WOBiIK2EnlTrXAqni5fjAnHUjKqO6zp962DhpR+p/eXzc2bmXUxFhZqjbI
W2yz4VoXW/hTCMWfDlH41d72UysaP0OGrdbyGi8GNdMivJuFVJ35/97pAlC/8gQc
P45wu0/7ztnstMC3fRyBP4Ah7nhh0gtdJyiat+xhm4WBwrr6S8OeDFEdBxOD8FYC
DeeUPREAXFA49p1fZgWjssOPTm01gAAGh65k18JKeof/LmLjZV/QjDsPHGUKO2Hl
ZGs3g0yKrRuaiLcB1dGtUqzcsRHDGh8TEfy40g7ZxPqIg7Sz5RgRHzyR8hnSvG5T
iixjnWOA7Hm3iaxmvk28x1YQBN/bsR2nbXgFAVSpaCyDaL1sBa1zbGZ/jq067G3d
othLIw0h+ShNKMeRsIkmspRsgWSQq0fvhmLlk+0O8fTCIBduuLDi9RvXJL7jNlju
KYZ6wNdVHiQlB3Nt3gLDhCx9x5aUeocoXeGSQleMqLtcf+pbTWW1pSrBxVmTr6Bq
SKpEajaW4JyV5dp5VRgQES17Bn1Da4PaKfSIJmBsecsS3HsSuyr1YEuXQJhFjKLr
lNIxJFuSf3RmPWKcPBNQvRWfybrIXxXnlTaNmpnubJ/6MstAk038b4AcQo5Dk2Kg
kz2ma4tCxjfstskMlaoA2alfzIjC+lE93UFAJ/2Z1JSf7ulPQSgw8kudfOx1v2uG
AmqpPvqhWv/0PRwzHgBT7sg/Z7uudui93PKz04TWjO/Lv7Gdg7Co+AdRkws+Ht4g
1pdlA6UzWGPc9SoRA+qzZ8htOD9spixknDds1NBhT+S+B+KzrftWraHevBXD4kLe
6tcybqAoRh3DqJ61XxfGvFJh4R5MfDQpAsUqJxedF1GIx7szxJkDJDGCLLzcf0J2
iCX3dPXsYmLC3zR4sWo1xF2cNawJFjpuA4GDYVzf80k6svYxe7feyv2N+QyaIQ6f
/mgLqYf9eCYCvla4WgeZ7dziWiZtbUKcS2/6qJMCZ88BNNOuC8BGyo+hva7Q2TFc
b/UTqJJ3/5m4Dy/B9wsSSPwywLF0KsUW+PeY+zbUkBDnC0wz03WY7LWuyGcEflit
md4uX1Y9wBsGNo3GEooKsYo/IhGuF5OaYyY2fZZlGvNStdrSSeTCD7OuS9KnoXDu
o0ZMzRWQNist5D/X9ANKe/uuhLYVpJqdtR6ZXxxUEG5NqAaBuHCPlDed7nWxu+vE
DIUPG/hRRUhb09wKgkUGMWGvcOcS6hA1yoWGb5iufYn+2yreTqHOE+GnPQBHWWCw
2QtwifFhoIRHWZjlAdrqnbAPm3stmfmWyJrzmT0wCdbEfg6tQZLH9Y8Qhgi9tKS0
gonEnS4IHoGZ+OZdYLiyOjqEpDkwYAuvN4cS091a+O1w65a78If4Rf10pEApTaFT
qmcr5bb/+Ag7yJilZzeNRYxvC28IC6m8JRgwoMd5usEsUkxy+ngwYsRZCcSUv/hP
R7OcrFvku9+OPhKlfrZ9LUonlZ5mbbu8zspvQPOIG7ZVE6UKtZ5rPUoqTHv9h06e
yGDlE24uB2xry9Y5RxrTFDqHyISLheg8jBZ+Ap6mD1hm50g73vCRZ34tLrHUjlHm
eU6AMB5PMyC9jSh6h+SeRobAukST8o8Nyoj67M/8FARcdiONqezZtB0HFxUW/4tY
Ov3Vy5uyByF+fCMXN7/WBziv+HJt/TmRjoZMkqCzjrQdbWYS3NHXkv/XW17Q6cHr
4fGHXqajY1CUlBOezmPVaXYaRz7n80U3F7xJ6g7GBuzlZjBD9UOby9k2CenHYwcc
EePEW2js5aJUtw+5t5KefvcgYkObKQ2fnYy74xcwkqlDe9fLysWPWwUEfFeRqHwi
wJG25d+N3L+0hCHTZYOwwym1UXndYDCjwEol97HLWkomVx1GBzg7RTGA5A7OhmQd
0ajWNnc3h9R9UbKEyYVyFPBu4fXdTutK9DYxNOdaVxnBMpac92+YXGhjPC9pM/mp
u5qQ3n1yjt/sWlQNh1D5btNyi3bApfmFftQEU+dPsyl2yVBzHPTK8W9qCAVWi7o9
w8dCMDbEZrnJw6izs7jz2xvB5eOLFyKPmt+8zKBZCLkWRn+saTNPMdw1jRkiXTWH
UQbBzjl4MnD2eBTEx1rXT7Bashec4aE2gYYl4ZM2qgG5rxQjC/7ewGJ0E0ebgDtv
4CI8QcMkN4UFiTS0xR5SeQdlnba0HiiMCqeMmbnc5LNWbVI6nTogUXKL1qBogx96
ILfRMTdrkXPBUImQhUKs2bWypvv4cWoJdwXTAE7JhAlVe5RJixip/3RB5umTA2NG
slZwGH9YE9EGG8d1r4+VYz1BT1/LTFwPowdrQSVRyy4EQLTdxjjG01BFt6UTxm83
UeLFZbKfINO82NXsRp1krWT4oP06fTPSVFsfs6FDIcripo8J/Ap/2Ebl4ZKcWuQ3
hHp+YBq5+dR5HSAg/HawA4shLiouWP/U68JXKiqQOOnagzt7FW/KpFuVO+mRnxMr
Ac6J1zco+tZC0u1zzQ5smKnuEsK86BccVq78eBptqhoOHB10QJ9KDs8Byjgv6lei
Zt4dbo467UamZrTTESQ9K/49H2bDy6ZcLaaT671SfeCxHPVwItoATWY7qe1eWbtN
CfB3gtecUTzGQcboxaHwW9TcBjO4k8nCFJkKGMJeJIHgCzZ2E9sNtsdhigJ4gtGP
RGtduD6WpzhvLFTtnUCHhUOsRUrIyAoPng4Yx3+k37soxk3Y0QEPmq34XU+HWaK7
HOuqTdKqj/L6yox/SsMc4b0EURww3tzfZevz65S5zzUra4M99ol0kTzfrPiSr3Sv
SAhxMUrTw7lSn81Rs8JSa+ek8cKYgASUQlBDbnsXKhPin5C3OIT5PFjFwRdJDle1
9pI6BBDgPwSe+hDHQOvopLBht28hF+VjpmVIovX1r7lJ5Uzinggr/eu6OmcpujZb
odNt7D3B9UcMmi9zkcEnpMN0wbI2HlbVHLDuw/h225C/hqxFJmvHdVJOBrEvyoMQ
Oven1Z/Ubf6Vy2l/BihcWHn9SXSEblN6q5JdvNXdUBC0QW5GOCKizAPmJ9M7flUB
3AvbdVvW9uTWrw89i+ZNc0JNL5RmFCcJedys5I9B90ZwcPebNE0SJwfWQ6Z2Uz3G
IpHRV7LGGMxa1CMXuCdZZULCoWEt0XFGNxeuOQa5w/F8z+er5i1fjY5A5qqQLuDy
slNN3fbNuXnt328yIj/UvkJa2lyBrP0C/BHxsGdAQc6hLxBNLzFXJmv4D7Jp4RxR
2ebyF6pc/tAy+UK14Fk1z2NH0i8rqoS2TXCtyS4za6J38ekO5o7fGomVm7DYGcTj
INzn0Z0qA4EtrU0yvGN235d1x6jcSGXaKOtTjX6XePn8KcPzu3LsMjEgTHs9IyZ8
+mglHMo+3j2OAwzUhEaaBLmWDYYfMVExd7Am7233ES407xPg+XH5tx7Y9TjrSpFn
ntYq68PGDLdoCXHR0UBlPBdBzyyDTwZEFX/QjmFn4NhddjXaURQUG0CWXwEAEiab
+kFnZ8aptPbJkYdWnEsCZOM0ImX/u+Dy6ykKIs+BD6fimDd3akZwgpoT6QlHw12k
lE2JhM+xaafCqL0GHUXayOcTm1PPY5gDsFaTAA2NE9HFfMUaXHpB9K0UZaDaQ8+W
pBKuYKMEgnJB3KSSFQSRSzmcjiejkaj8MvdHHawwRjSIMcLyPWAyGLV/gYRatZ5H
C9wFZFI8Us9VugTn3ZPRQp3Ww+TVMGfVPuSk9T1xQ3IHd7/hLvaU9i7F+8+sJFuv
+qHV/zzxhLjVkvBGwioCXDPQTbDwCZYk3x3raQWrv9bOK0Vnq8pelL/xQFnJq1DK
U+KBs5WDoilTKfqcK23eGvTHeIS6lfOqm//TkvBTazT0/PIUEBJNYaUpB3DOPbym
1P5vSWGGMngn8qt20l/HagTjaFYgeoKsBIktGtsPzw2LWjK+xYXc8+81aFhGSp0L
HgWx3hNhwI4rJ9+ZxNvMMDaysCdzmz+l6h75FTCmFcYXuDu+W6mWB7NpG4NyxFDr
AMAr7q3iRUR4EhMOpo52a4v69dEU9mlp8s7o9xzK6j/PCnec0oEq0T+1bDHmxqEJ
PBnIMHC3Mwf2mXHoBelTHz4AFEQTHb9cW/+ztv4LbFcC/aVjXlgxYDyQp2TtKPlq
TS2SNxc6rpjxPkqwwZ0UxyfjN8AXDoIQykXw/EcnYSXOr1o+GbVSb+emx9ZdCDf1
2i9EGvROlgdxWgCgBn2Ok0j0BnkMi8skPNhzPAvCIi3vyPXpofrUqUTK9ezxgi0P
4i2qqqJoFZoZKi0COegGUZQVeMbPEnhv3UHfztbJNGfA+krkGRaFxmXuINaUMC70
9i8tcpjDqZb42eNZ7Oiyp0hk0wY03BWKsv9Gr88W6kgyYO1kcmdkaXEhjpjqgcJo
KxzrF0xgpXqu0gQgbvdKot0UJ4EY5BJjAgObQKmyEPzH3VnWMixF2G2rRvuWQ33a
hnxa0DDC0VPhgSbd0lfDI6l4XVHrzmmTkk49iq5RPbgDFl204DSMkhhvH6+Av6nJ
7wIe2LY4yyf5yiI/z9vc/zSww+yuTS2YyNM4XrOKNGGVUZkHqqTW61COjoanQNxT
xoh9Q2ORqyNVB6atXBWtTYJVsf8MZg3wVRUN0rpNoyThnRs+uL7PjiUWCIXWPms0
1+lPk4s+Z/4O8VXE9D4c6Uy5qNWceaQdPjZGC58ekJdRgHnLgQK5D7vXTfD04+iM
bm4zh2wKYGcLRhb5Nh+MJr7uqYVP/a2koExek8RgzeHQGxFCRhUt2CZTmehNHQ+g
ykV7QI/QcQsAfrV44OXB/fmE+ah3w+6WgQYEONeYZhPjljcZIawHl5yjG9vhSWve
cvgx5wIU1P6ncC04UedVqsUpgxH0DZfv0YY+rnI8tydyDDMqJ6DjiuI5YPApAEDE
q1j09uafYJHvE5Itla3HNfqbmo2+JCAikXtkp26QD5isqbmU12QgBznegGjlJrro
L0bl856/92eUawl5j8evpGYYSXKUDuEcGtfiAf1mUN+f7PJO3Lqg6oA+jC/nHBfw
fhwrhtvAHZBtNFjPoxsYKPMP/S2S5v3ta8X29J5zPbKB2s8r+WK+bECCV32RzY0n
PYsxpZ3uI1cXxkpoAjGh2UyS74lzlsZIyB1vhD2FtFjyIkiAIhhs1XgtED27mvzY
4iAn9D4qdf3ZUW3C30YyDBlpmxxbwbZ/KZI5pUHmHAQusAl2IUTKc3a4T5SXY1vq
XN1D4YNyDlcuYcsgjqW59HSSfySZHHbuDvTejiLsKy7yaSFV+qC7vBDDhPFF71h9
83gH8UaL2xs3zN3zPeUHavac/iFRt6WPzXnXlUEBwr0ej0DrapxLBGBYDkGjReCQ
qig4Z5elpwl1zyOWL1ibnN/tVEFkoQo4VKM3JfArOa5tOX3Z6Gc8j5hd4HeSuMOW
tDbqQfYyC06VSALUvyKIgT/E6rn+4ESYsYak6XzV51YoyoWKDA/Ue3+2rCAlvjLA
3/Q14CKKyJxBLo9vyv7YBUZTxJ5Up5i/TqHpcHHzlNtYURqcYSq6lZ0O9c2qWWN4
EHMGEAg6ekEoOeGsfZiZg1gAoaU7r84yl97DAT0arNj5MlHAfif1gGqYA0vjm2oL
Ml7GAtFDH5TFV8B4NrU8piHSIQPbAZzvkadYgsspMpoZ30JL+PGJIuNF7iO8Hus/
Cw97eS5f7FcQWR35KDB7UdHDuGfEhz9geR0nXGRAVyY0jQK+hhaZSOfZJkrd2dSk
65asKw3Y8QUQcUkrJ5mOncibCJm2FsrI8GfGyE+pUSpH5ml2llLS/6k6lT2e89i8
1u9xJI8Xv2vY4OFs2BIXGsMJ2/5bXO7TAOtRbcGFBMYkD2EOLJhsTqZhoZClnfK+
/ElFBLyKunITAaWxAlIs/Bu/cyiWNKwezBDTahMnGZyPep3IQiPZUKI0YVxFRtiq
Fo/LxlpRaqver3xZvN3Bv4usoTtPOkAzeflFQtDTKU0M1f5uSU3L8rfE3IDYt/MQ
43iP8WAi69q4WrcAG/qlmSBAXmbhRu4T4gmMIc/D7wKBijtM2gGT3u6ZXDq2kcyF
1G7I2XPBd4MO9IVyRUoRR2mtXUEQ+gS+XneedZSHL7NjtANFKaCdV7hB7Nx4h4uf
g9j351UqLamOLiks+eQaHVfxOL8IeAFn3nMFsqF091axCq/4reqVRRxA99Ow5b45
v5i9SrV0KC1ER04plyJZCXXX5kzVdW2P9hu92vs4EFO/KlAsB/bl0U1pJ/3XweZb
Buz6UUl4zVrjSV8Tl5++hhgELmAAiimUtEcQFUYKoJvILBgOPi1TrGb3uh57b5O0
DpHVt+tA8lvulPN40Kgd6RGbwwRx4VsdZHPLRwzO+hWZl1wxuCOfgfAbxNEu6dkL
1TRQMDNfVAdXtENe2MtlHhQ85Uz+Q2EDE8VzlbXITj8xxb5PbmC84SQlKChpoFfA
mn9bjIL86c2D4tRHnOTrMcsmC9DmRjLmbttUjcQPgUNgJoZiy5tNA6ol3xfsF/Mm
wKSDfwQak7yKeFRf31Eftsa+veJGbIoJscJUgbC6vNN5xWmVVhjg6/jeSX8ljkA1
HkRYtt8fsP+8XVpa8OtOjWephsP9wV9WJ3Hx3JhA9MfcmFZAu+g30zSvKya67q97
8+l5EwXYto9olqSr6/VM6RCZs0XohOOqEGUD52BGWfgs6IJNuWugIM8pSq1O78Vb
X8/vM0lTUNdY6/nNQD8hvSI6k0xsOWEoF9+v/nGKXt9dskVRwTGS0X+zPveVAy5H
BIFT0Z4j1c97lUnfDIiq3ctYRgSxnypivkizYF6WI779Eq0ZfWxMHHLAYy049wrn
F7J/dz+EFXPcRYxb1LhBRQU5Wfh5DmeDR4vleDJ0GX7iarqf8ih5ktGY3uZr3s2O
t5Gv7e5pSRCZ0eRg9QkG3bq0uVuYMUQvEd8TU9jPMaJXt78pSLjhsU2rVM6s6gic
TTWELqeBKMd+KCxOX8SXvXpruyjNzYAkXVAKWvs3LVoG/W4MFmxUyYP2HdkpLQWe
s9lvQhD7Bi2GV+s/8z8i0luZPEFeVcXCz81Q25Zi1QrOfZGBEIGmVJ0+ljKqtHdL
J8Du8vb5ocBKk9eKBgf3r5CkeS2XDty1xarbTiS+t1ZnJ62uMw0iRmt0hlKhbhOZ
mc+Hq8T2qroA9FYHCRjrkpd64FXTMIT3YqGmUn18g51hb+niEFwYc5F/XJ2V+1Un
m60v5Fnl54dL+tdR2+y8+vtl/nH/9Zn0RsSyxzV1oriAKKCO/iPqpfiKggqoO6+a
Vyw+HpsSDRoXsNVxnYM6hTwB15IRJyT4zxV5Q0YZACjvVK/Axixr6lm92Z4x/ld3
LZluoN77zFOLEX9qYEO/3hcqZKNfVNTeq0ECmxKEu9a1XurOoPIkNN/6jbARPpQS
E3B3uIbsKw1i/G1khfHoL+PJmqGPP/zG7u+hFfeJtKrIVrFBRnbSuxxIzFuPVqAW
OfTdLQstoOo74Ii4w93MKca53g5DP1HoyMKIjB5JEOPOLmn+czajB2fcWkLWl7vT
F3i0KoZErSIUMAkY8k4yeJU34Dy0j0uQtla0Tj3nYuYcTV52nXAUWONMFCvq1wuH
9CqaLdZXs4eU29wuug3jBqA/maWjnhbq2aqiBjUj7QRy7hgMrAPsGkAKCJTTO+Kd
Nu5NQSsuJq3glePMnY1+QWuofnTPMNoyNnNaylrfloN3p+4yxj5rTrUVFjCo/Ej5
3Ts9fOD0x3KLL5Dv+GtenFHSe82XiaFPDUZv0iF2FRveqkSnaP0vI/kkMweACOO9
WFpTT7ao34IGtcMprvfRd+SOYsmnrjJeN2sQx2WmPenzaYrziHQNyqEROxsHh8gU
2jApFfOE5N4vC58fwCEohte0zSfXl0njvcfYjsuwR926eOY2SkDKEPVL7v1Ja/AD
UfqvOf06v+wXSR6+OxHspBF4HykbEe0YHaeoCe17B2jKeDaCtXvQe9Kn53eBn/0d
EeUuopKpWkPnsGzumlyJd+vLAmV6MVvgqKXD7vO1MoNMilLgxIYKtW+TkEiTjLKb
HucteScru6V9QxNwrInybuqZRN6FTtRRP4zedOC78P+wThyPJpI+sGUziRNPIxO1
0GrzSwZIl/QGw9zSuOwpFcOntSp2i5O109rkuZ4zRqCE6IZoJ+QokbNK0CzK6Nka
hGGf2nw0BmKw/5v8vj7c798aqn0qKhtltx+gK/17WEb+pJsAeacPfAJew+TaMS68
Nvrro0N3O+U71laUoJH1bQTPOG3cIAbcn83lHzaEmrY7dZmp+42oHCHeQOGsdeXa
X3cmM0dpBH9ceOELsFUA1V81WAQpOnqGcxI0DrqQ0QYqMdrp2e1F6B/3G2TU//Y/
G1/dQXffCK+AkJaZfZkSXj2S/ka7+Ke/r13ADL/Q/lpgAuS43veClUlenAPgkCw9
6eO7EUAf84i4TN17BGDIE8reSNmR1D3l9FJS5exgoTFjwa2XijXOg49fTIg7r7vL
3/Y44/4ySwfHIL5bLtGbVuVEK9JR5BApMepcnprjnIUcErz7VZx4fOV+bNyjrPsM
Hll6UtesNJWroHSEXzPOtNaU2v79K+YnjlHmcyiWNu1iotSRBOQkMKgKR0AYB+by
wK8MBST9qT/MFB8WzC/+Ytgsi1khe7Nb0HvnNVMMPqPM4Z9QxX6pxDhPVlof6mia
1XRUmWXQSU2kCYBot79XCa5oJURP2KK4ZCVOmfWgy+/RK/tZ/+sevPQCfxXg8Loe
slBYGK4SxzEJzN4eXrIlSq1h3gSiGTLwve9+H7B/LQKPLT3SnBHEVJgjuH8CdbuQ
ruKGFouzR8l9pqa6Tp+XdkkjJ9GAbVnjPZ94serLASK4V3nRD6XtAi1HRLFJ0lLn
fljzcvK4sUv4xyFHfFcxiYaMMhMaDiMeKZxEu+1Ma3bz70ZA1nb6CFyK0IyAaorR
wbpPXAif1VNjuM28gEDtn+ZOmjzXrHA/AjEUqiDQTDmPce5mILWo/izxmEzp/6X5
cqTbw9cN4JNyAMsGpsstDY/b/pXjTko7p5TUC/kBs45KzY0ngePwMYV2Gpsl7BO8
tM2P4zMtzR3pYq1Yk9d6/TFhP2Bsu1NkEhGExeyqW/XQ9rmF/xzTucD+QkYiwnOE
By/Wu7w/ZMF2d2FE1wq0P7bFyatDFstc3BCegasSjawP1ODqaBLW4p2koDL6SZEx
NMXCjK+3arjuTwb1ao7vQj/SRUr/P/0TkloLXML8+6JVafVbZMsjDLQgLQMp4oCv
d4rvOAgoTXruPibfJKfOAuEqVcdSK0biuTY23Osn1qSlsTXP8d77GH51NXPYcFo/
imygHRWNtQTf9+jBHMQIfQe7GBwL1D/+mFaey6f08KuCl0CbNg1F3ATmuvDd4aUs
TdPBGUEtQUhfusVDT/8hY28aHwLQXFhbxTyhBTFlKcgcpbWB1MFmNJ/DYasQ8aGG
Ix0evsbR/q0zFCXvRRFb9PXsME0TX8DyzW6mV3LcmMbVyUXrugu5vNJBc37PIWnJ
ZvmeQu5ePzZpfqtCqSgQyvlXB2KsxVNVbr1IpRrB4Qap6H9KvxANA3m36BKXm/Hr
R++ABXM/0GfwVbQkaa+e2EofvVNWAyVXJSiTK5BmZCoTTAFGmScQ3dgAlO7/Dj09
MqbnujRmPN5uPJgYeo3XS4sMBnLzobRf8C/7MLnjFanks5oy5WnG9z1c88+Wgeo7
Q/Z7vXFMFa9vTmDylYukMMmehX6DOE1egPe9rO2mLbdjfZc8voYDHQ6QA1tDDGBA
6BpZkPmt0iCObSnECS2+TVZawwVlCf1HcgdH2O7pTluIaaLx9I2mvYV+0U1n3i7y
4vFyqa93OKCe0qqWFRb9tGIXJs8BTyR6HSzNZJhWi2uZ9zJ4urWjVdHq6MZURewm
DV98+yGcS+VSNvnnPzQQETHxuN6ROmY5CuPvti1jZmvfE29Rn9eeGnQ/F3QbxUzU
y0eGW/aUSswQ7E7CrtE0rOx8E4cmFziaMXDnvkcKR6DVzX9QsIn7nllMSGJ8dB+U
2KqZtz1UK82zbU3QCdfo6a/FmU5iO2KB6ESb97spM6XGa3Q+ZC34klCZezzizM1C
Lc3wRQi/r8UGCTqCpTV9aiCpRkeAS2j0ChDb7YjcLtfHQI2zfZ9hxLb59gq06Xgk
oWcMVDapjXRtNkMcYYABYpzkJLW3Dn8CetCDEHXcOIQXw27mwnLW+J2WTOP74MnN
GhZK1qQUC3GQkulg6NferqvmhoawCkFIMQ11oLYfCacMum8loj5jxqvgWVFLAPi/
Ui2t5TTtz5VByTeJh3BULA5X2w6YZm3qAKukmiQjZLVRzdjH2c27cl5tlRYqxk53
zyBllCCkE9YUnOetbHOZ0Qzu+z036QcsF6IKS3TyzvHMG/G6Jk6xfcjdov7QArRD
nPjnfMboSBiNevBHIpYUQ4HsrHqmZdKaadndEV+DcZo6ZdeVeGwSTEEUVwAvOw95
+56kgSroyXPpPpaRNqjEtTmTYV/lf1Irj8ODzyMourrozOtA7N2s54+ZCF3wmjHA
MLzdWk0VzLWpL6NTERUCIq0GqqkEvO9FEsSrhfWcaCw7nDju27Ow6GsMrRIS32f/
B+TZtm9HISA/iom9Lpgz9d0Sx3QD5t7q/4kqXE3tBZ4ppwYbvvk91F/+7mhH4Qed
illD6+1GVAwHAZpu5nqNIemWNglq+fbN0SQTs7w4FgRGHgqKalIzSndGkNKsP3iL
e37NQOVBRgkZvwTQjuCxIm7BcOVjCY2PwicC4qyYP3eCo+myM1ar3YYKxqK2ytOE
1uBwQRN40xQnX1lZjSK33LeaQuvIV/BoaIS91ju4NA2pbRbu7Kkyh9fcMMUg/5rk
Xj5fGlmiS74Tx7rI3qB0ZrE0FIGQ/q/pq9Y/hn3k31t9YDQhvGaZteMsO91BaOWG
nF4H2N6kAuT7e72c15PMZhhonSCzFd7q6OgRbvlwgYJT1APH63CZnAHvK2WatV7X
LxX6UkrN1BRL/ng72oxHn0r1TgsPTENFLGx5RKmlXlAiJIqyKFCvPlFrOVzPPn7R
GbtkqnL6w+qQIh/RfMxJUOvYLM6IeiF0NURkK/Z2MEtp4Wz2+8FyxxxdqNrEv7Dw
P21EC19hE99ZxLGUvcplcN5R4qoDr/9vwayDGDSCXdK6LI6BI5o0w5RT3chhH0xP
7Co99LURL+2+/gCAV+LKiwcd/5OFMJwwBmWnk4ewdxP+WeJF789nu/9ulMl091Fh
gTfiih7ks5z/Ymt/yITjdEKL26BqZrvV+xwH57uhXZmo+Ytc++BiujWl8tImiau+
CvfOhTkYzwsCLUi9RHprjSr6wcYS4tSFgIyAvnJEsmg1voZAqCpmh1fcfcMtHV7H
4vy3uPLrOjGEdhghxpwAID5P1Ylbe6aCnRwKPSKlMClJ50aqIWotlO0532yUQIwB
c7ayCEWOG244REhvJRjXeP7Zlnr/vUItBlTOKI1mLM8BURQyx6Mgl+8gdWR/PbbY
qqV5F8Cl/HmXRrcnwE44cjiV8VVnY0SMtrJZ0MpNmJPCtgXz4u5Os4tzx0/1SsoL
JnHUNc9nqFZpU09s8FYWcSECdrITAgLbIC0BsGodFkNZLfGTfcF9MrbfeDup9TKL
4aGaseX3tdP09fiTRtxYGFH0+UmbpWjrEbm3O3QK1k946OSZZGTlnrj/8VnVXvIG
C2Lg1t4r9U38RqTeNmhOrMOVViTR2nP1EYvVwh+tHRTVKhEKuphKsBqNpKKB6jM7
HzVEjVhOgJRNwXU5YuhhQMp88TM7jwAM6GY1WqWMUk7yQIDTY6Dsr/BP/X12rjDK
zpiDHVp2eXLRg3Sv4cB16pQ9mEKvbqWVOjY98aKYO5xMmP1QwzqCoAyLnXgBXoE2
H+zBuw/+ux4Jr3zD6eib/2rtvwZ/N2e/Bdl6N89e9zdQFCHCF/h8bJ7iXZ4DDuOb
wDgdakweL3WpWVyRXrGkKg6OjmmXAB7ThiUI+JWqLLe+ldq8UgxcJCKp3Rh8XQpj
YgLYz65I6bh0nr5gQFNZ3L7OE7v2VxJ7R1tA5G1L60+uxEMjnKIBfXrJZgUWw/EN
glpDQvPnCT0MKWu6zHoulRm/svapLX4hRLX2t5SygmbASf1ChsJ7tdPkzYz4rtRV
eM5p8lwH4IGnuOBANmQ8UBM1KATD4uwgmHKZNYeL1Tk8ZfhfZYTsrQBtisYDosML
7KCe8ny2NvfTf+7TFuyyN+hmsUEwn9BvYVablfmd+xgxhhOQwYP6X88eOP31VWzE
dYtJnuwnwADfhnTqsK/np3/DBjBVNRPEXLJCrn5M+PVdfhClSv1l8Om5zun45PBt
Rx2xbHGNbdK4QvM8CvfqSCT/KfBZav71k3gC+DUAEaofbadc8nZmcu/zBiYq0VPZ
M+5iPDKUUr9fkpURX70iFWP8BiRYSMB8P/Dy1IflxIpYbRopBSEpe0QPffBtHYD/
m2LKSeHyeiWi4k4Kj8LDo7an7NL8+RNf+tPJIsjA/6PX0vWDBBdEmqivtRHwRH01
FJ0wllq9mJ3KoN7ZI4FWFVf8cTGZ8wF6Th66UemLMTBjSMzSsJCDRlLsWXVY24/j
HSH3oreOnncMmk681OZFF+PPEec1avjpioJ43Hh1LkoqSHEwlgbwy/9abERdUW6E
dH0k2DnS0PdFdm1tG+nNgyCFCtcwhDIlxlfzZhPZV0VUBYSzt7e3WlND+3sYFgac
4oazWn9cLXbFnXStJRXAUY/fWfHUid4Wt8PAdKSlv2Ew6gtSea+gVwqU6ltgLrzp
yRwJNgh0DDnRBkPXreRaDOQ39PUGO9VRMBO0bV10uU7KUJmzG0xKklBMRSBY36c9
0LFIUoWuHKPleoHzZMqg5xS86SDvnch02xSfbcToJjVro8LFvGvIFeQ8rV1Ci+G9
UgqrvlGkhzRE5T7/ZWCTpXf5FVLEujp+2EaNdegKA/Yvo0jLMWuXZjSVBvM7kEt9
OFKSX/rVcUAl8arzZiumUlSz/BAS4ABANnrYJHPMb86HiddYSCaOk7Q4LZJAFUeT
ArxzjQJjbjFZqlDJ4QC+elGI3cVQB6O71xlFaOy7UwNCOGfoQC/Ztf8mrf8fUGDT
RrBBRMsT5aJ9aXvEIiQJl7CHfruWk6MARUQaG6nqwofYUQvh2PDfJVPmSQiuYXnx
Tarse6Dbz0Dlv2jw1PO8zgeSJx0gs2Wp///Fl1MTsrs8RuGqR7Hg5s2OxL4qNrDC
vA6Vrya56gpjz129Tujhv8nVtsVSDxwio5c6qpeq2XoO3X5cqZTYTyHByzYn7iID
PEsVP/wxa2hRdKFrU4c/EQou7fozrHjMoQdIsYEYaBBlkqvxOCmUKR2/fzMcgXby
Y0yxvj1uCDsUUlNZumoE7ozy9H/jPZZ1mEPb1VhAgK741RMXY1c6Zv5cTH1u0noz
FiCQTaMo4WnlmaU0UgUhQ2UOxFbme6opCD5JvwDaxIy8cqxSqjlYgvn9KSp+ukGj
irCDv8J5cvgIFZqjq1Zf9XORw9cCju99eg0izUEdI+OvA5BwFHcKqqYUALiyvmfX
QfLQvD0sWOCtLlCtLWPNOSFC4sJ3EVr2sOOBN4NYGuYfjLLFBAlN7ikQ+zKzw3Ib
PhTftZ8uYqyW5+epozySN+Yz0wnCCTSww3nhvPHeGZHr5U+vIF3q1Vi723W8EHiv
mYA9V8s7+QHq8BFisu+qgjhvWdLP3bbsGhMeRAKqa9TAXbaQDfmj3hyLBx6osLHs
ZcBKhCew0ZXywU6rkST0TvQgrzINGwQX9/QnRy+1nI9+bhi3o+Se4S+uYx2IHoxQ
P2c8k01jPkxhX6Sw9ipMsm+sO9sxyjZ2/ZxnnUi9adfkIjOZ+vOSBo3EaxBBkcro
7GAZKwa83qvcirMv4C2SWrXFK4CBh9XadZRPEXcrOQ7YLJ7kD4R3AWyb0IZLRwnC
H6E+qGlkDrVfqLoBpdAI0qIu3KKyJ/Bpx2l8P75cokQr8XwoEjqVwEURq1XtclFP
Vh5mQrAFv7eL3EBB9z+1VBV0Z0GrLHMk8Td3mpCjtCgvtwwD4Iux5GiltwG1k4MM
wx0LWoW4UoZeMhhd0Aj7jSxqKxsYN4yq9IhZK6Wllz52QRKRpzKPZvK/jjKGLq2c
C4S9tyxLDqjWKpFTbdEA7LoYFeaGXOHTmFdkBga9O6p8B7Gp8ADeDjd0nd5yf48p
aSSochG69mUh+9jhkfN21lQlC2K2MiCsLepATMIMbYW5RCunP5FDgwbANf0w6NPw
8QFWMY8qGOyuBIweakU+nEFsfKJo0MCvZHCA7bUdOEVjo7RHQBcFOeJZN2Vy4e+9
/aXY/WR+E6iHF1+ZABtdfsh//hz86+vrBFz89Qoowfl4WTw96ARKTCl9LQCyGIvQ
7dSIgnkIIqasOauCyHdKm6RlBp1EbajxwQgnRM1LQ7Q3Cz7VGGCK0dmInlyS9nhk
sBdTo2ovUz78w3r2N1R3ZTMdh6cZb8861RpPjg0Xl3ccb9skvNnNuPJXICXA6aPO
/6BGH4xek51X8KCf3FNg0f1kGeuTrTKpWl5813bNFKzYz1C3sXOO6X7F0JhZyk9E
/67lp42F/hMrXUyieV3MU1nOW1glQfvLbSa+vrLdlWMnv8E34W5oWeAHqLV6ZEKO
GbQHZFsi8ZxbqKFw2MYKLKk+BGjidtw3LPve+kI1QnJdXrhjfRo0p1vNetDoSa1k
4/X0Fr/F/uRCGGKTdwk1Iv+Mi6LQ3oREft+ykWDYVSNG8LAqhgiqSXw/dLQTNwyQ
XNo9swD0ohE3av7jX8whD+bgw2jS9Bldb2C8PdfY+JtRJQxmxO/d/LGUnxD3hb5u
uluieshK/XuPAbrmakbOFSCWty9lAaDstjbQNe9lGee3FATzcZ/4fNbtjTi+JFfH
T6/nwhRFlPpZ7E+vq1vHoxuihO79OM+klW8FSkqS5DU4ynI2OW9u59ECDU/JXGyk
NlbCyzms7XBo4jzp8QOcoJnZX9xxNWM9up+9tpw+5CUlElU3CGVurHO7/roNRJNx
V4mhHj2WxXYbc0xcs0dDFGE9KNIg8ZY5gTT1cPIpYpyrEy1UIqX96lWK0NwgFfcu
DO6nP0sbOze0bkLW3wTRZeRrHe9Bsc3rov8NU/zYhOqmBLC8D5/WI1XctAzievoE
y5DetHLUzYW3CMusdOZsgJj0usQoQR5lzmGlml5ghkifaec5luiYEg/U62ObByTi
RpU3+Exf+0j17ASTLSeGbnnjy5oe0Bq6lbVC4WtsZPl7/Olc/bFoJ0CCe/3pgKdW
oxb6nYBAJLJDdAFqImrVOvW5HWnVNh5ECjjM9ErE7K6XfVSSETWSgje/KZJyAJlP
wPP2TrbXLP5qvPWyOEdaayZlZz++cxraxeDBBzunQYn1YZ++se7ilAomyuhbSFD7
qTZjxG85yh+wzsizXIGkEs0nIoaIRR+J4qu2Zk2P0+jXl8msKwB3NALx1g7NlN2q
it22D0bGsTyS5JH513ejo4I67oOMjCaC1TQziZe/l+8cU2O6YDDBScGS2qYArtQG
cgNjtzI4Ol5IFQcgIgXXlY8sraFie4H7E+wlRJ5mXqadiN2m61xKHCcFrTjL5dIq
PVrG1dGi/D+Kx4LGUTVArrSeVHl5PAwj2GXweY5heZAZb7OisTR2CaA5BU422hOC
11pBoHxWturnM7oqKyaGa7IqGAEMJRMmq5ZvilZlt0Z4UYJyekIp8b+yL6I0GvCd
je3SdjlMtz2WsNvu1fUAsgwZkGPyRocyFuleuEx5d9Q1xJYNksCAVsnX/kEE8ZZF
VO3YEg7fcKdIlYjsKxcCAJs+h6wP6paXUUJHvGWkIA6kRwi+KR00PkuHxF33iwOf
QsDedFe8kx9b8NN0YuQ7xnsuydsHR5cP5xj/S9Ta7bng1ZcSmyqtALg2pE5OgMSw
ThAK7cxNzBbTHcnAkttz/G3KGOvAUO96kY4LMgAFuGo9Ih78sYr71DTCr7eRQwcB
mGNi1s69S+GPA+kP2uwORS2IJWc7MQW2NN1CudNT/MCeLeNl2oOqk+lbyQFHCnPc
MBJVwUCmA1jEfwyFunj/CSmYvkVqm4em584Pe+E8dNHlSipvfusrrJAQGuaUS9cK
ic0EukxrY7KjrfsYRRtwLMM0+VyEOoh9H9kFkaBgBuuZZZbNO9nM4MGuLpSaaEs9
nmX9nNXT2IKTtM1IQVhuBo3CKA8wZKziBGTUexbmnSpp/DXJYIAoODRz+2g42280
8XfrKz/07wLURkeWz9TzPkQj8shcU7TXFY24sZYGN36MypdFlBqymFoEX0G0e8b5
8hHI3Ef6fI0Lw0vAZLc5swQ6sLhN02ZR/UK3gBMXzdE1g/Qq34wBXU5l22tV8E/8
FkkBwwTDBpCH8EmVnEdWUe7ZBZNC0j2BZgxEXgPl3iaMHg9uAUbGxg+m/2alHcBg
OSGu0drIKUM29auVOE/iC4/+IGoI1M3so3xsO89vKN2KsBnZizMFwgxxhJXS+vlp
5ibdo8vm8IoU/3N+zUUYhw98XGsks3HbIvfcZ0LwYEpmAFDDmo17Afd2i/SJq6gA
3dXSy3ZZHzOp9Mrz76Y3j/cVFYPg4diIKVptQC4aO3AXKcFKNm9l/pLldGL6w+6M
DVlvQzCZR4QkgEHZYomDYPLt4VNUkY0pjrHOWU/AcVsOpYsvFph/sETbIhMtuAYI
fjiBLEnMW6EZb4viKAIQf4gDArQQVGkAn625R/637kz1I9NmeYgTKbGAny5K3reF
boWDqlvFKz3g3aVdkQUG4wCfX/6yRugW3IHNe1Rna48D6V5UUcvMDanXAV9d1Jiz
ZMH5DsUDcpNrorKwGZHXexyyZtv4if0jvOiHwC+KVAjpIXdbmh6nZwhukb6Rx2Q8
2BfdtzmJTAhjmZu0xeIy51ptLP5EE1rilAdjjlHYvmFLIKlUU2dh3TDFKu6a2W80
OxalCgFGMYNW5J9XmDF1fF/D5XE5P0NKsRPSBmWnvnKug72Ku3d0tjl2G91KmGyO
A0E71EJDWCJTit8/ONGA0HuVxqPFB+Q6hteW95Cewo6b8hG9Wc8DmJb6Pn2m4fJl
taD5+X3qRRs6cpO2eOw64luhZBqyOGR8kiVm2keaOhuscTX/4RmUeJLvmKxEzKeC
WLa4/EYpqy8tFxss6cyswN8Tm70lJUpwcbE1rb6U55/WekvYPthxJE4QD3UI6sTY
8jLhTAPvaOpildeWaNb4iw3Fg6tDMIxHfqA7584ZzOV3nG43ihWcF7nE2sah0MnL
NLUl7z9NYemHIeOkDaLLIJRdG/UNNtjUOzQ6bHDu0iZzRplAME8nC8sMx0otss4M
XIuNO9Gf/cjWrPeziLP01QzAiUKzq1+gr0VkNCmcEdFEBZaJEW5MMpSAR5zkzEgY
VgEGsVc8jUGtBksVS5JIn9P+g6DT2n6/TlrIgLokrdvw0s8+MaktReqNiTRaw+09
Ig/wZT1ilxLm8Zvf3dQ3LafkybqHtrKgH6MMfqzy0PXO6wLmxiIdf1cR2OLtKs7f
S09L3oBA7fgBNGu0wGSs6Kf7O383qhVMp6w64FI5VG7VXf7lbaTrJpgjy22cFfeA
1tIke0hXqHkBG7QTHxaE517gmU0p0TfW7OOE4NxMJpQyogcfNCqpV5Mh0PCDocl0
7AE7MEXsLF2fFhf4+zKOC3hT44VLUCbZKe/14H1QekqjpLpG2EV2mQt2SZ2d2MAr
nfKzIlvlwqnTafOcMCFpCZ7edOpDDKZMffdDoDg7uYNdWCWMaG4zIaGrNZwl3cfd
BSU9hhsE8l2m2P34DhsB6l1i6VsgpmU3xPaAXcGb2OUBB7+G9EtoGbGN5d4rcTBw
FxytxSpjTqR6xBxPheje+SJJYVA3TrB/ZVtx8kSVtotPjt9f31Uuosvab8PxwaGL
Ug+CdqlJpqf78FYFP3vEm4BzMXfhoCCcHtyrfSu+1Ejh0qpK1TAR5fMQbKL9yxWy
gT7RDJhdfdsfu5Ji6cfpnWJPl5HgADcDkrwQAHk0WYBWGH2PUMgMWDRybmqPDYS1
yDBANoG1mepMUCCeWxFotFZc3K8kmlRC+agC+ub8FBGdCFLooq9Ce7QTuwMHYnnY
ZPsoMBtrZan1Hf5kZiwg+L40p8qZDwHep0mpPwN9ZCveIRh3jK8oBvKh/EBUP0SC
tDfw/sjB/oB9Zjmt3Gu4tlNdouniyeXEhwH40hAbl/ia2Wyshvpqx7vJVVyqZTK4
LFVIgYX4sFb+yJVvwrNl6rn9Y/0qR841gLF4nBMpOzTDhGQeohfFOdMiAkTKk11s
bkliaT+aiOi2p3fI7x74XXL0IsgwlL4v0fJmoTZvH2VspcoTcsE9hAm6BzprWd0G
2sjgbuoMbI45XmKSPtUW60ELdMVeOdnEkkv+bCaV3mhqdCjlcGOXqXzydOMtuG/X
ydx0gs56DkKqiCXlBw/djcNMGEGG+Bn/XPtVd+qrQqivQJqxJvHCb6X2SGeRwIY9
nQMatVHx+p3pvwl1hQxrzuJlFF/lDN6Z/jrxI6wHdrhM/V4j9lNPo0XmNeEbqYC3
0xHCPH9CyfKiwiqommO1YQx/KHRJKnWvBUVzNXyArfhzdqU52TlunKYNGdpjzHHy
es6ya5mSBMFwA05S23uo9PNHQFHZnDNJJ33vj3WqerswHlRk9Tq/5fgyNhGIPrk6
oFw36l9SG8FU1ZWnI4DW73vYRy7fYH9tlzwYV1hlyz/PjvU1Cx6XLFWzhA5akNg8
otHdd2dEJ4cuVscjZ5tGrLFGRaFxOhYqBopaiZwejS/KP/mcsmcnU/0hREzD/W5P
UrkwLAL8gbM7us7Q8RMuZuyS0P7AgisohnSafma2EEaZe+Anx29a29i00kL7T59S
vRXp1gXXrZczmruss0S+1oRoWDRHcMSfFRXuOOJAhpx143lESQ0cisSAjoU0YewV
erFPodq8bwIhzLZAyyqkwzz260Aplk1hhQMx+5aUNn0P1XHrROS8Phwq07RzG7IA
LmvhlTe4O07eYRnwKx4HtpiNDBPaFx2x5IoUB3M6+dUYNrHnslIjEa7D8dKjY9KP
eA/jqxoQ8siIaRUUFIT2zOPYcdRxfbDtd19zMEKaBXajW1D9LhHrlAQp6KaI1u09
w2pRhBJZBCWfpH1AnQ3+SNUrjRJZ87CzETCnmc1J2FR5jh0yaXUMyw9g7fyOsoIW
TM9LupCIX8pWbOUVvO/S8CaDQlRYSbpNhF9mu6rNviXMNg1ZbVU12Fpdz3mfGxNq
TlNR+TBOjoLWOxvY25jA8wG+O1DVXxhIn7H7mjlYN48sfy5efK9RIKdVWeKubM0P
+eIV5tK6RpPdx8r7LY69geONdCtwtF5LqJKI3jloGfVddt3cHgcTIC1Ii9mqtTyf
lMEEPxbJ3XCk4tsSi8wE8ruy4rKFixjAfVO7xpfHhu8nSxNI4tPlkBbOKH6Ax3RW
IWsn4qoqUyKTd+9S+wIolkLVCE2S+M+nEcyDMoDthT/W2dC2pQ074AVElHCuXBSQ
6QTXiyjNMmj0BzaJXgc28y+56CW5qaGhfRaBWfmclAY2QWgys8Uj16iWD5s+1/Rl
dMhwd2iqRPhbC2Iax9fbsto7GTbDRZqNMtevjE5yyZMrU0DJl2LLvIboMaK6GnnL
SoBSbKkZjjNj8Lmej1Jqkv55I9TRuwbrZxMqGTiW+B/PXzNfsYycO8O8j8Qm2ik+
WpfU4ICO/A7cCZVOBaRj4ym9pZ49ghlkQ1CXzgeXHCGfHFVCzeWNeRVRoPX4hTGu
QHDF12opUlu/er0UI7m6Ij0d7qqJcHEvYA1KdbORjWdykcccOHYJTHg7x66DSdph
+CSCHJDOTgCTdYI3LUB0070eHHzv/b7FdBGxEjcZGbRiOqCNuQNTH9hhbvwer+Ls
2WY/cTyUNYaORkMkRfSd0v0J/QpHCbN5tQthicFTeQ89lqxeBzVi7Ed4uAFwPDX6
8zoZvI3VxYADe9VJz4Ab5GwwNG4tK3ZJ6sAxX/WIUfv+y87Op2VV9lS7YjsuMTtu
QfyM2p3K3Aj7XUCoOsRYe7s1nFf/+iAozVOTPgboMiLGfhSSlY63E5MHgCdGzmim
SznzIwIdDcev2DEaaJ9IH8Oxo1QHMovl06xJMrRLCyfEGUHht2aqGPW0yaGL387b
XRi9sSF2O3NjbaI4f+lF3XJ6s2qsUJwXz0TISRrLQlgbx/vom0J30EsFoZLqplp4
ilgj/Tz7I44hHtnTgU6QZ31EDl0hQVBOYswGgUvWaq5VhHnXHd638ViG7/rh81JK
Fc3srOL1gwwHqqd+TOEQ+aYAoYx13ccTrhfYxRzCK/o/KCDy1E140VIZddBeoYSR
7Nk9wggl85mMQgdzMNIOswgVcZB4tW8GWtIz4uN0cgUE2TYRr7Nv7XNWfhE6ExGS
eQj0f+WMsRd3yNC85trsuYBF06ecqcs18w9HFapYkHFuEjVcmc5Llvca4Zqkkqyl
F3ynWfBfKHB4IJKLtXV/z8ydd05TNs0/pAtA7YtqeJCwHcZgycuUxpvY6P91PLGF
aHhLZaeLlDcHxxKk91skZ/7r+mKUZ2asaomsun7gZvOH3o3K197RlzMVielSyLJe
xHA4rHXBYT+xjPPrEhKEEzIzX5aP+lPkcxFcOotM6KacNnesdOwl06ri51U2mdnX
x+xjusD1qBWhTL56biZozZo6usK5SGg+t7VxZdlowBmunVU8jjhcdBrkwA8r7hyy
3Ap56MaKTqU5YKuw8w/ghGP0i1HkXlC9L7bHP/cXuPsmzREA5Vbc2XR9As7amIA3
rlpfYksTMUxn+rUjx5RUglRXYNSvztXJpwK5800Dx9dzCmrq1DaQdFDztjD8tIeZ
Iashu98qFS45ESyinrWPKeS4JkOc429Ujw81RB8W0qplgQ4g4nAr7jyi8ipjCpSx
El4wvHAKxPaTjH/0SlX3HwFCvxOfsnsMXeGfW/cU+xjdrp78TxmRpin014cZHHPf
w4FbBx2Si96r4ZuJDPDl696+DLNLpKqM4sLQ+WgERzcsEqtW/iVthdeRKDcWQ5g/
ewnKcF+jXA18oGdFV3QDh3S7FWSOP+9A+l4v6ppS6BpvIq1NVkKSoKVgPHxuXuIV
8EV6DcQGR/Qz4HuBqxWHzCgwmgxa4GfGnNtBu8z+aGKxEbBbNE0BsisHYef0XMwh
YRH4TcXcCXzg9wDIo2DMygHePtVKT/VOWTzvgmPc3i5dbEWI1nsjloQqBa0lbqZc
US8aTCZF+n+dYSzFaGLhiM2XslkXBx1qy+DcWPczRGufIVGh/I5i06urWTsm3aaE
L7559J8hg3S6U2pX3QAi8GH8hpwEj3Z2xNPP5VORaYL93rtcKzuhlWj2DoB4k/jC
BPIOYRdQAmzXC4JP2bGSNnXzbe9kX/1VZ+Gy1FfeZOhPDFVQNw8FSFirvVG+M/gd
l7LkbH7TrzQ9dvVCcxh8K1MxB6oGwfQEMkJDdd8SDa2xYfeOOvR2YHjbrokl5b8V
388V777M7sZ7BQ1oP+VsI3/z7gvqFpgl7OeGRZVrQVwCr5lLZCu2byE/DWbSQIW8
19A2NnHZyDSI0eOHA2DSR/21XG5S3MN0k61gxn9s1nrJ60BvGmHKvbMrAoJxAUKu
hQsZuKj6Tf2KUQ0edCfdN/z3+NjGBEo9OSdzwQfeCdB0ZQijk93nkKjd4eQe6BAf
F/+x3B0k8ydMqDx+A3bo1EZbRJbjdODkUHDvMrS3ojSKDFHi5NV/fFS1bFQ5dg6a
e4pVaiwOCIB7re/W+Tg+injo2TQLy7rKAY2gAYYW5peJHXaUH0rAqzeAJF7bG1/x
RL5wmOe9nAHD5SJBYxV8mL0mhWcmNY2ghrHiOtXWWgNLR+UKVye3V9pQ+Yqyba8C
PnYkGkUDlrJ2kTcR+jNCe9AQQ5XIgjFEE8Msz6X+V5aa1UuTAjuN+3LP0fSGN9PF
myYMnNiYViRVgDHtE5N1iktLDQL1Noq/OPQ4xOCcC2O8leGxbgDWos3E0KoFZkaM
gPJEOb1QWX+yAsVd3mQq4HrssfGagsgmQc1AJiy1v4xeqN6sIiUfOnWLGZq0//gv
gKFEhwvZqD99s4cEkCkPc5uCafxJ+pEv9A8ycEIVNlu+5X6oF3vQRL9/6hB9WreC
oJZDSxyY0HpIm/ZiUowwRBn5kJxfhVR1Vcui8yggaFlEhDp8GAOZJ+0uEh96yFbl
d7C6b9HZiCBo0bMl2SuUwPuAn3zJh7mO7Ddh6lfcsX/0qb/utZhngF1vLWzaCLFD
IowBIJ/c9lp8K5V5waXkIxfqvhYbBsICPZiRKT9hYbUxVilCJ8tiaPkxDc6Gz9Eg
QqQuz2ffSTSWtdVITCEmQLHlvmS6oPFUmKBq9gD5AGYQxFanNXcRQkueuOYxiIHh
7h6whTRKjUkxDJkmTqOaG3ORI2Rjhxt0kchJqPZNbmulCUCQ6IzY/EWi3donUKzi
A60q4WkyZY5lw5WejQmJ7J7PC+evMSzCu4HDWl+78LWzJRGbTbDW5/+4sJWnZVUG
1QHVNSHHXxAl8srpKYBmcM71Na1B6EUqPpkgMJTy9feYD6y9UwtM9nz7SjMSeVRo
3OzPnqEQO5cVdR8CFwPRyr1YzRBQQvMsmKKvOVkDM5+7+c4vo/AJkqQYJeV4mVKt
bRKLxYKZeN4m9nzOJOcH/LrUM+5KrgbugREoeee06rWmGPQdZqStbajhF5u6jhad
cbmrRJ4x1HaFNz5/Akk2ATTyS5PBmCTChEFBO8yuH3qzSZzJMUWzMLbAOf+QSQE+
8CuSjaeCXgwnsX2kObM/9Oil0hjMNU4m/+vXDlOKouDaXNF4PSU9DSx2C/tE4yeI
o1DvtGsmnbzEChbFl0qjGm/hGnD46GxzQzP4LX9sBAj8X6aYcBLPQVASVjT/JxXU
Mbr4foZ3a9gsRyBtFpUMWj5kcgq7/OxiWZnKg9sSJbWatPBiP0iO3Knym+jwrXeb
YSQA9oTHe8lqoFmaIuM4Gj53/UWK1ZS+DNZo4AzBKiLkh4cOZ+XkxEURv0IBHn1Y
xOu943XYigYneUqBp6WQmHCs7DWOyuJyuR6sLhJdehaYI8h7/rpiz2wV0M08x+I5
JR7t3zE/1vD3NC19Wae6Cf5dm/KmC4Jii42zfsFzsNB0qkYawa3JRD/rQL+OeCZL
etyWxekB0ugmFM9aMTs/ESUIWY8+YUR5JNTTVSs8mHK5Oxgx+3YKfSReGJ4hrzIr
vVpb5m54UcPhnxOuY6TOGKH8+oyo7RVFANP42DJlK9c4Z6wfLCt+zQ2s68KfOC9B
Ktjq5ILWUCHKkFDx3+PhSdvfcgcn4umI+YAFj/9wmSF184saCu78mJgydcofXFFa
gdL7Au9qwZHVe2jkQ6mekQEXgLQkNrCe9ikBbN/pP6MLPNCWX4sPESu5lM0YnR5x
UsRP7pGhxqTp3xmuVaMjavn66N2x63TXE5C1+5eeypvxXIV30JXQq0Tz5jOd5qZ7
EzT23JrKfSdtrUPATyTJ/1TXDpzhVYyuVILolFbwgMVPkeuZjQJmb9rg92tH76TJ
AMVHvgUhM0GYyv8ixMbBKIGch17qwlSdxFswkmTh9UYGlIOF7iJlREUM8A0qLNj8
QE52AbLuM7LLxrkaREBpiNXhx9oPj4nFEaeHwB6IvJYR1Q97o1EXNO0Kkh9COWiC
0bq6ErOfjJrA7HNefcn1MbZk0qfjZUCc3yn/Au2YAKOj3AedXb2JgCTuIst9ZvBQ
ThBFNjJWVND1YRtyY791Ph7qzLmFEl4mH6bCBsDDe0dYwJ8j3feZXhUNk8Otr3hg
D+RqBvVlRTNnA1OveNuiWsnHEeJu8S8V9Zf4lECRpgjtb+U1xQByAY2ZlminWr+r
BUlFhqq/+NCG34yM5zddv02GnSZ7b5RlNVkdqrHUvS1MbAfgEoTmG5V9nw1h8M4P
iSc5OM+e46vsUSqZBpBlSbwo2xUdV9H3B/O73my7vkJNzQ2hm/nPb6DnX1AFhnst
m8MiyI6S2jE4yXHy2E91ItjmtGocSiYBgLTppQp1EA4So/icJ1H9NRW0bodvXdoX
arJhM4bphavVO5xgM20+ONFWsOQy+CycurLFV1lWJEaCMC/ZrlCBHWILBAPT/gRv
KAlkjZWGdGE/IKafEO1Y6fBMBBX61Jb1UkfY8cPC+yFZzT9OprIhAbb60RwbMDJK
8CnwrpHrYH6sizBuLcghDttEoiJo/YGVMobuhzf2mmvnyfOulMW934SFDpzN1ga8
wcs40Ym63uP8O+6TCmm1fURciuPKNjnjkm4yB8Ij+Q/77qfXwbYqu3FhvVO/Jz0T
rNHwaqKvz/GniczhenqdQxaAizwpODtlpTP7TfD2Y3COEHnlNPTmOwmhsbxjptCQ
qqaGvLeDW8oPcV9aZuT8xGf8AZcAd+HgwecK2UY5nBjiMFh8tReNf1xTXD4zlAwF
hSwg1mRYwQ/ivV2HqRlgPqxH3nD/5nkL/L8YzKEMf131PDm0QI/T80udbZbMvME4
5kPMzlXlGUWez9zGmf3oLWXBy5krSQq4x+REzs51nspPWl40d7BQnxisV6tfLZG7
jYiMYajqcRP/Q3OmQ/ShztSqXnhFWv90SHDMq42ipIy1BQ9Q5hiI3+35U3ZtZw0b
FFBunrEBJRKkEaUMs4WB7ZDOa6NdoGYFOAP0Tb8HiaJ+pEKozzFqIoYfMQVQX7et
PLjiBYR+Ka6TFk4x4kMyxEs077m4ycC4vB+YN2YBwAosfvqcKXVg2yAo6JekaEQC
Mg98asuDs10BCdDe3DaT6DMCD7IDhmXyfpAdQbtCtkJeD92kizEGo3zQ6MIvjC1C
YCn/7Wqy0vy9A18ktF/LgP4UqVdKRip4yyuSuZvHuuTZ4MLiJ7e7LA+Q/q51MQ2y
30N09X4IPca/dNTDrIJkGaIsjpUTNUDwcn5gN+wScC2DPNP/ruMPudRE577Z5/DE
Wbsc9RcP5YyX4Qwcmf+4N1EpT1H39ekOh9r6A1koZbbdsn6MdcKnJPLSUYVwj5ML
1O7CfIckOFHxVVKrkwfuu1/BmJJ6/q/OfIw0l+eAQJBWVC9nlryDd0c+zX8JmvpY
bvK0SIGUScZI4Df25Z6lQkw1n1SyysyCedXHDvnZgv73QdyZCbfwqiN9AZ/sw4F/
fXsK7dWyCE6kvy9VEDcV32Cbd44ishJpGZOLcQCGlVqdWjQk+3X+I7j6+cGOzpLH
6D9i4g+NVe+XytWIUTPJV0v81wCtcL/8DOVbYjwiCljslK+6OCQmUya12UaCH1rv
tHF8L3lENEDtWxyAFF7eyEI0tIzNe9BJSOkLnDOhuN2c9VNelaOQZwcJVSf/cw0K
faSZzt7/kJ98o6Aid/OgR9eKhtTPCfPDN+1DwpfF4xN/hHve8Smba82JQWKTCEyp
HaF0J4RPoQ7XjUD4rmi/rSzQnAUGBkN6B0omuQzLZ//gzA+aMbTcrl0kBzFXrvWb
x6+ig6+sNhBq6e7wbwuO0nhHQQhTQDUnOK4DDeJ8aaY53Ikee1COy7h029sSAclP
ngVleNKSMg5MOy8Ru96NyCS/lOrI2890i4edWIuNfKDR+mKY+QM48RQn9qijr9CI
Zdtnw7uVsMrDG+9aovz+k8stmTWuulDr6hLhxVuwGPULjYgsTmBMg7WNyi2+za3/
hVr/D61/EPMUR7oHTRUeV/sKxxkk2FS1Tk8UKLgMhXzn2ec+e4EAXXJC8fymGu/L
FKQZvxJv+5MfsvwfyoUcpD5p2Sb699ST5j6NNstKQ+an2ABAJs+EGZ39p1I9eHxA
IYjha2/h0thlvkDNJWxiSmq7nYTlx6NpYC1AAgqyfF/tDWC7M65TAct2wPHAbl0X
GYW9BmURqmxdTzBmSK05InhkKCcSIlxpQ3uU0fwobYVGKBDDlqEYhHyf+4ssgGfu
s+5BLXS6AHhV9uJcftAW6UXB4TUVu9AyCEYxeXVtmVpUUtqVGGFdORryS3BAJ4/1
Vc5Jm66Y2ZDbx01bScfJtdjPeJCafmuewEZK85Qvr/9iZtWA0HENcbEJ84sUiCDZ
7wKZdu7tHBBzFgTjRohGd/SsTvRao4HKNl7oQZyCGJrkyQ0+LPGKGW/4tebRdKlZ
Wni9WJCYkqR5fUES3mJ3+Bx0JMQoWeZplMybTIpZ7uMlJHw5V+oVQY5tV2hrdJd3
1cRGhTHGGmHoD2rwWg0vSZl3+LhXjeTB9UqLRp+ACP6uCDTeTJxFJuq637lQN6pC
4fxxCzy8qHUP7ilq2FJ45yHcdiET5jl7/0v4OUxU2C+DM+akXt7maVd+lXrgIM0V
vY6KEvctViP0GWnG9OipywQafyLhab578FsNbKUhTKRw6h38P2KKmeckDFSnkvpT
B1hGWyYbFCZO/t5k2dB6w83tvs62XEOngXbdh+f3/4jG3LhA8Vx6vb76YeGWYvXB
cWpUuoQoHSLgDSLLUw4LRX8kO4qtYFhr0AgS7JmnUDTVNzd/ELJXEhpcz0KdlkVn
BtpR6WrsrkSbBmyb2nJjH5mtq0Z6ni+VzpFHduC04SSLgxsXKny/VTQ/wbyJeAx9
Gqb2a3YPzJH8R3jJQN+ATokzD7MTOrS0rCrqUzbp5ANXxF1f22CQjR09rCLNEPRy
pyhSwsPy1SqOMoqn9VjuwgG035lki86c4laL9PMocS/4MINnir7PaOMhQlNK6xFk
lBG7k6aCKKy72uCjtlXHBMD25rWeK+oYfuCZbddRm3EBlSwgH+TL/wIn1Fxmog0m
SXcMJvVa+vFSQPp5au6PdRT8m9NDO0kLCz8Y8Z7m7BUcL0bIDXOdmxDQ4rf9zvMs
`protect END_PROTECTED
