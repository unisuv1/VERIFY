`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DSX8vs4Zfz7usjkewmwQhlTZVYr2LmjeIG5aPXX64WB8zZ6QrYkn1+82FQuD56LA
lBR8QFNbwKZ0hopbjah2CEo2AjIVVQW2DY51jfOUj1DrPzlPaq6ZSEnM6FpTMVtM
nNLc5vI9+com3cSmvh3t4Cbilo7y6+SZ3W03ZrtOxfhy2AXVg+b4d5h3KlCBEOcX
1So7R/xhviIY+O0SW+dM6KQOfEDNsTRGmiHwY1RNR4/6JB1YN4QRk+ox7B3KOieJ
UOoan/fs4SYT+GTrYJAZKk71ry6pKnrpdo+M6q7i8YYSsZRWdb+pan1OnEcg58Ko
NdeN/dOAjWZa7GYUlJpzhvViTAKHVlYQRvZoqO2W/jD+QYy3K8LA6uIcOJfAe67U
FecX5S+QJPr+r7zMYb/6KHtwQdq9HohrNlYzbAI4ZCpUz+9ghOaDz9m4KqkqB1Bj
ZN7+U6vtsd8svn5ixkf79C1RetGFxSID9Dzji1J8IVvstS/MtXQgdJ+o8pieVGH7
RL5EX3fEImlLTG1UCsnpfholtRthk35F4rNRsDrrAQIE8fZ/mEzc23Ft/xaEWN5k
p3dnunj+wM01+pj/2YfgcH11NXYKFmAIqsHhk4ncfzL3mK5kszSZAeiwW/UZUgFt
/7S0kOTYtJMnrF9hd/vZWhvxLw0vB7NeaXvuumQ8asuN6DdjxLkizeiGUD1h5tFR
6yKPupVBDdy4hOdIVQlQazmGZzfGh/ylgjjEWp5zPc+gDY0TjA4w2OyVO/G/RuOJ
qUrIUlNRuZI3ZCuWGK5lfEEtxDiAZ2vjIpHHylA1Rl0/EiSDPLoVazdLl+wkg4X3
QIEUZbOQ6UsjrnzYu8eHkC8zSdkBRdcmCd78RDApic1h+4wP4/MSASQd7fejJLLS
/PTbygv3JLq37VR4HRtNAVfLBSZosQU4Ha5qIDoSWHBp+B3yB3cj5ZS6aC8qruyo
m4D5ENs0XCcx50BUUK/baLFn7SRAz1p8i726pe23mR1zTBYB249y7OCYFfdwWxPQ
5j2Rp7y7BLGf+cz9s9keWKk/VnspYAjEePcQJlb2DtKYnlk4mn2gQ9G9dDAzZkwk
MW+bVs+p5kcAs8J9tPzozfy4lXXQM4+nVfioF5MWCcB8WGplrpdhTsH+ET8971pZ
EM/3t8WDXUtch78U/E1gLIg3RPekyr96i9cqFLvYGUh7I2VTncu+ynI834a/FywQ
ZYZVebVsA9CG4m27jz5eRYU27r+xfk+TwzLTKixT/2orgw+FdRTeFI0NptMd3auO
ArjCTLB/5QvIaXMoBu6nduoN4LyZxrDqXDFX6NfzDpk/vLFyX3/cSS9WXbEPhcp8
wO0mdM5a1KID/4YMn8CTwxWe4HocVPa4naYB80gZIUB/qhit5AWk+bqTEowQqYF5
quYERhMw4oT5Inzr6wErdB8T0dbs39tlUQBeXvI2obM47d8tZYk7f99JL5vEUFjX
i3Rd+hWvk31ll3zVcxfwNT8oaJUlJ8q7gycminvMdO9Pe/rGuPlNpT3f5PfPZQMt
U2bpF0bJZVK5lURQBIySo7Lk9fSccqXt07Oe9w0e9a1kzPOmnZYuOsBiyGXLg+Wg
CqgoCgJuK9r3Sv6tJZG0FwmvE4aXzTFdlICh13mBmSZ0a+h5iJRMhtmPhFPwPpoj
tOd66habnKubBHhvyCF2wmra7puzerAwVVgLmJuKEWDGUjKV7qMqkh1JBQZt1wdJ
d8kBSDrlKy92sqwACv7VUyyvx7x//uIo+eTXeYY9JCHsYKIONgcuEdmDhGewFHeq
jOVr7eMO5dtPpMf44LIahHk9DXTvin51VfSAkFk5iRvaMTJRW/2oUX7I4CznnjBA
y6+7Zzd529Ru397luSDDjYC7TJZMsWmNgEVOUxCfPc2leuSIdsKuE6+jrHZitrCn
tosAEowj9sl84ITSKaZs2i+xnomOFakz7MP/knpIhzt+WfWaiodl2ohwjTkgJYVY
TS+7xOzJinYvzs2xTBbtd0lIGLclimtMpBVqKb/bTRomWSlrzm5t3V3CR8wSM6Ja
uGGWVi44zMEvkRIoaNRQmTP08GfWgvLUiVPaV1nT9gez+cMXOf8zueH3O89OIdq9
zNdYirhc0f0bWGxOLeszIKEm3Op/MynxLwsZwCkiWDHHq81qQSTX9T8XtdaBAm8R
PrKBsBRU8LNH5tqHIk5cGvj0vwlhvmHubCXtmcG6TrW/i1b3oDwwjknylIT2N3jV
m364swcGg1pb5ae9nxonqW10jT942QfwWNiZHtjekiiHKB71JrWbGsov8rXVWkR+
RQZKfyKn0+7Gt+upKG5DAwhVY4hHSNM0595QZ08ph2k0mbDkH+Gcj20GD6LXyA3o
su14zTTWafUil2e6DD8VCTo85ZbdWwUq9TQXTx87snhx/38t6qjw8d37vMBmGhfy
bHI51aupwiG9RwSqV4ozv3vR3JVJ+jkoVR7woZkZFGfRQjhRG8R7FLJm7FIhusFX
SnveUxynRb3X6hLweGfnVhAlbsW0LvFQk/XKrdNgau5WfgWypjmisSU2AO2ULUh8
VTm+a6taStB13wsS5hL4SJRG6pJxVODlo2JiRV/oQCCTeM0JNG1yibi1UDysj5zC
XHGWgFTDYXnnGfMYRRvd46IViazaY+DdM9c41aqE+qWIuKAvRIJ0UpFwlRxd4VnV
tf30Iil+U8kcVcbz5S5XluV9NYigshu7yJ6UiNDRoEwkOgFlYx4+AbaQtXtZ+2sY
P8M9BcJ10P9UnwrckY9Ll5cQM/xeT/OFX+Ar8Rle02NKGWGNCcH/PwuioS7b5ucZ
GL06J6xVHugKGq6DjihAwdzoNtyWStthg4Q4GoN0Bj9NdWpz51nn5Bv8gpB9XiED
bv8kzN6YLurog7Q1lkNKf4kE7Ne9HvTICBe8D8V6ZISfgPQdsZNiazXn1kfPWVvH
GgQwC0cCOvqm0L7fB0OZtpOMB7l58U7Zo1gQPkj2fZ5AOwi7I8M6AnlX6D1nNZTd
yNov9cPDQQOE+1nwt77Dwc+KpgGbGF9OD97Xa5/XQ1xISoIn1V/TNcadNkwocgui
W2z0GHnLyY3sTG40/F280NzBcP2/kifbKxcWckpLS0ChdtcTXBRndZx+b2qsVoDP
xRLmfz6NAgC/EXWld0/7pnYS0iQ6JWoYNXtBfoCw0pqJVsho3gT0kCWnN2OMcu3p
pMSzU5ErpL19FLTBgYnPviIpt9DIRa5ocuKdVGSZAlQ2buCbqq8aDhXcK0nzQWkQ
JOd1tHE+9xz14ODQu1c56bD1XF6AIFDn9W5pZ3ZfStsWLc6JK+hRX9p4gy0tig2v
L0p9hb5eZnmBf4ezM+koFn8kYCOU06S/k+Lnxb20o+DPtDvaW3J6YoaQ6mMP8V4O
8IUwikvOF1rFXwDMrgkHgl2JTd37Dt68pU+zomf8Q6ogemct+TLE0u5HsQW2uaAS
eCCOPGIXlGHawBuQU+L92MDAXEtFN1tE8eUHma4nEDLxJsitU9h9YF7hkK6fXRvd
myPzORKyO5T51TEWcdaT1MWCiUPCw+csFtaF+6FGlT9ahWfNfxc7keGhHys+g4Ka
K9VjKDfus5q+20YKsjAWg9hhc4s3GygI70GnBm+2n2bAy7gOU74+F9nsO2NXcdBb
29DpGMYAcGjDzisp8rd47J/MwSRqM0ZdmxeNIGWg70KAnREqFVgSv9aMC+rKwfUh
4GiGvh6qw9R1fUbtZtdD8JfOzeN19b93ehzpvyVqompRJi2qOLTcrW1Gmq309Oly
re+BfoL+KINJSaUS3fwk59TQfXyzYGCfNYU/2hZ+BMz+tV3ziym+X9U2Aht2Q5Ja
NlfLdbCmCA0jnKjaJUK1l2Y4drkZO0I11bBGv7aGG3P3tWkqGTTd6vHMXvLoll6r
1Gi5Jo0eo8lACCwAyDd26AFIT6BvWH3mJRCeWtcKgIVP1aNKb74xR5COrgHWybzO
BrSoln9ck0lK+Tdjq+zY5g4HlAkOXXe1y9WoojIyP/7HucsGhoz2uhKUo8oTxWAv
3fA1SOgm0u47arFWqFT5CajZRnn4WNaVBpjnhTz9y6XD8kJnvvCLwKtMMIf97fah
R/SHHKbRd/3uOzWKnuzewSCUiXNTX5sgu40GR1yQl8r3Kqmx/XRaZ8aoCBQROAES
qT/0PLSsFVH0iho8GA41l+tiPLLqCwY2Gjeb2x46KCAS58yz+ZLjn1T1jZj/bS/4
PPzO2/hhswi+KE+8/oyZ2vzJaTOCL1eUaKVLcglE2hMIVvhjHNN4QHUPSm8aG27W
qrpoQGZ72ZJJ97YEWEfVin246JgMRuxMOh2Tn42bWjiKn9H4tsDOHxjWce3nHSiX
8yCCqsVpQZbG4eEx6muDVndvk7Pj93CHLSBTNXDP+fQ65QyCKxIpX/wb+wZKf2GM
Pbmozk2ynT3/UCKpIYnLgyus9jqKrFYJ++UbD4HN4T4mPMRpoxjptu9uxaPLna4l
bC15TER+9dozASGH3oFPqVoFS6sVjQ6dlaO7KYF4xj6n3uvi/qzSUA84953Tagdw
IbSMq8Wucm5qaJvlCqd+1bRb6hsKe5k3SZBPrhhpwqSs3NNYTqIyvJH/mf/i5IMe
dbV+/aZe7U7HYKQEN2qDcuUMKeqcUPElR26I0+H6g9dOStvBb0U80CIAjPkHXUEw
D4REdbNPBNZytDeYlHDC8xIlA7iNZlx5EUitkGuy8GhnyG0mIsiieaqA2nJhJC5D
wxgZA/YfLNWzMDd17PNz7QRgYTCQq/ZXkCysp1UTrRPOsd5HLxQXqOllyxAPRPFG
ec99ClSTUIAhE3a0XB6n8HNl4eP9XLtkfRtUUyxAzm5igScj+USpdY2bDfu+cj/R
JU1igR6DOWhi86VuQfoy7pUP1AZsAEsPxTecody3+tYcxiPNbKGVOMiD6LLKXCYP
1i8njbT1CIp47oWoNd7QOmEXu8Hwg0Ci4mSZL5cFl0L+diiu2a/JuMSBY9vD77rG
AHueUh7jnhprjNVBS4cfA7tFVIKdfSt3OTdA90SKFhmXESW218Ce9D9HJ4ErjICa
6TQf4FC1/drt8zgoyohQHRe9ukdazYf4ziqIvlGoBo0cbCaKssINCR/fVwpH9Ohv
GFDwlm5W348X3GmCSV4ZUDRmI9m5HIwBmV0zyo9JrG//wa3hGz27sQDUk2VhW5Vj
uw8z+4+RJfcqdeQnwKknN2orVYQs+i2EJJPF9gpojEWfTdjxUc0Hh4V4wlm7NyE3
n11+VihoT9AR/vpQLFmgnJVkHGneXt4V7qJfoE9uANpwvepM6bRZZ99ox0Pve7Ff
J4gQpeV7ulz6MI6dsQxzIFv9xN604fgj97F7ZRpRIvJ/7sN2tAskpLdVeO6zIIR7
Sy7eDk/kDAxTiHDjPomiyOiePnG/cxa9b9TI6M5S4CoVWfXjQWE8Kg9cRzkCYsPV
gtZT/cc6VQZ6xKa+n1W9PPTUIRpArU00hMt9EDY0EGur9yRXnQxrBMy8KBkjdSrD
2QPGK5HiHhVsQ8ooSIc/Usy2kGt5H/zgxw3Ad1bfM3/n7BPsj8bCNLSkGHKMeTL5
dFLizAgtixiH+MwSC+Q6ChzZLqNb/WRJWzr3c1JFGHZQlpsqhNmnBRLMaJYnKdSl
sEEAgN67qJGWUuXIvVNnDZHOKXpXXM4TpwgeNNRtdZZM3cJXeyctyMQgNhCCfN9V
2Zuo3PO+lPbiOobP980KvXDfEMPKpyd+oTchVoKXx1iIuZkGzEeeAHVVgwzhs6Ng
TAxiBtDt8hS+OnQdnege3eCVBnSl2LWE4QtX6X3B6KJyeh2OJazC6T5qnCuWoss9
yHxViWwqLuNiFMAfCYsXwofr99xIYFz14lnXcienNnMn8/KXz5ZLf0VEE+JGzMFe
IFUYeWDID7Wt+SDN5xlT1LPB5KCSNyr3yNXkzJjrsBKoT563WpT26T3cxH0Lw+xo
HOn5Xf55Aipt9IGoSDXlPA==
`protect END_PROTECTED
