`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
z/BD21nubAkp/W+j/ZglTfOygt123fzIRqSPSwX+aI8aAZ/QfzYVm7AGpWXEjYfX
aXYRA3ll5u7mee+eRgy2tjkir6d9/Nj8GeSoTosnaSBnEpYY34GPpXGSOQgFWzyh
84wG0f4aySmncxv1kX/AbH3id4SIXIes1/eF/podDGkxJbIIlhU0ERLOEmI58MI8
gsxaeSvH2NbHdzshxL6dVGx/hIOQGZKDlVacUGLGZX4JJjm+uV1xbGRwWhqtsiRI
GcUs6+0hFg2TWAqIDwX1rfFYBu8brYTKh45gepK0XS8czCEuzZqyOqwkywpdO2fZ
3Hrsjat7yaEBAZcq+rjs2Irj9EBAcTLEtsiMeuOZQJ0GypR3lAto9ls7G/3STrlQ
86NpbuKlchbTQ83aXFn3vA2HDz4zzUD4V9m1HTL+xE9aTuV+E8aHgtAPtgYFAez2
iiuYlYVR71mvys3GxEE6Ht4Icjmz0MnwoXuIBqGQ8T2L6F+XPSY+xK3UVFQWoiG0
Fopwd3daCa/H6h+/Ub6QkffZj00FqeIf6tZm4PFzbv6cw+pRv6mYuDOEPyG2PL3e
W8uIPLDDIITJmZ/06T4s/F3IaA/o0jy8kPTeRtRGUb5L7Hjkknz39pHmrdp/gzLG
nw78SVcC+wCA86yPiy1KZZXJwcAA/DUbHIxW6Ol9foTWf/astpibapJp8Ox7ZMcm
yFfwb4tBJJt7govwb0WZF0XC6WlfLaXVC+Ko74U3dzs1nj3I9woP1IweN49Sw+pZ
n4eUi/A2Av9XerxkTMD7l9ee36j9hcBliCg8WoiZPQ1iRFA1/UTVRDE4t/dWvq9G
5x6bTvHDawi/iA6JQ1Tv1BP1rFnCwqwR/fWYzd7ge09wqeqWMTr2Ic7VRkVh65NV
XMcu+yQ3M0aYV12kJgI4N/65zxp0YAX1rYkyRPFZ+kTvipWo7CuWmlTSQ/CnlPZ3
w1JkJzy7jqfKU1Fqb1OimHjc/t2d3YYkFvEo2vP1KHv3zx/8uNJcodT3ENJH7Efm
/B+BJy02PofiHvmFFpv/L0WzbujYE2T4WB06fRlApQRsUddOTE5YJUNGWXSfAxnK
J/jqQBTT7yNu4lQpUF/vroVdMEi4iB8lhViQnBNCBR4OEaoDCep1Tm+jiDN0f6tU
Axab2Zgeg+df08Wsri7y2t2nvgZ8Nz0hbL66dcf/QFj693P2DoHRoYrN9dtJGfOb
cQB0M3+Bpo3Qqglzsy3lBO9q0Hl6WrhFWf1pNfp/z1sUi88MIpSIONtDZCyfGjde
chzvURkRCPVY3YcGiE/J0RC4zpADv7BnxrnSThQLjq35P1ZGQqspwwigofuAEd2d
V7hfyTZqJvVQSbwu5+Fp1Ie20DdDwaewRW9ttstL2ALUzH9MpR8aq5HZHag0zbQZ
5Pb1aE4Y1G3keSFrmUDS2VClcioCHGFKq2XafoyK60wfxlh9vVzi5TCUTAhNF/zA
LDEM5IPaSF/WM8rqe3xE1A0hK9rpFzvDtVmNme+iIjVnKeRsIT70gZD9/zxOisXW
rYQTOQXX/vOQm3Hq0gNRm+pVOMwdC620bnfP8NajcjNdS1qnT7Ip1GaAbdtQclWs
NiLmch+EBBmO6Ded+5/oo7xwtiJoTs1hPo5fsbtEKENo6FnO/XPWi6blBhYGlvxp
qZCU3iT6R08mcv17hQoGvfY8EOprJ6Pk3T+brjeaGELZOCbP/MnrmPMugdH7VmcF
xw01StgQdeAWYo2o6QPSfgKaFjROUk/alg2GVt/I4NLnLPlOc+IVo5gTL41GDkJd
gQzW5x9ZL2D9KKIl+0lt8m0Defkfvp+eWs4MoL/adrndOQTbjuOiz7laszthh/uL
0AmdF/GD1GRDqci1BeghSMt83bU0xvlNDzBcNV0EghPQoj4QTo5b/9/AGg/PNLkQ
oFSllKRT2oWa15d8PTPpLSsk0OSEHOAwtQskmeLoMjteUjGHmXvcL8ZmKrnupRWC
pdhVFn/Rnm1qvTECdyaLGsM0nEK4Gsu4vsBxesgumJ0lHMVJ6kPuhqKeC0cMtawQ
qQrJfdT+XNvC/2lHHx9rxPbuXnS7Z4TqOLzoYxruAMaiWvZdqEn6Xf5hFmHy3IPX
Eo2ZtdjS9ktMOGhEG1SJZ9hV0fZctPnPwakMOgWGr1AjBtlLuejUgCfljs/wvOww
uJs0BsfTKdLJGFUVfK+mNIKYPHtNJj+f8VDu0W5GBiwCgUwYFXPYJeDCoVzbxAoM
CMIU3CUkepNPfZZiOutBYBLnSA1svasiic+Z8ye4HrfLknHr2nyYyz10Yrf8/x5h
nLt//0SRux5juSXseblpWxM9b58Y03y6xPlbWyC0Mi6N2wOQAYmmoFjufGu0BFsU
oNJotdsHaULwctMn//qPhEm5nO6hBKQxijrMlfxAHVwp5aPGj8J50+i92ZIDP0Lr
3wD9YY/Q+mBe7DiV1D3m3x4vftOIZBL/V8afxMbSIcxIljNoo8Ri8WIx0IgMLFU6
FVlxH+y8Fq30G5nStApNK/FJi4QXN7p2PEtEnBL/iLYkf8I06Qgow2XXNIrhcuPT
7c584OcNFx1ySuHJqE85MzYnzhrflGKv+N1g1S4Kc8t/cNfBD4tvzUPHGP1S3CJi
lYMSLnJntlyeabwMGLs2N4XNdr0uIFVDQlVwfWBpM/keUVLQjG9kW3MzcBxS671c
e4nqJr2XAXtJWwtjBPOnK1oe4Ym4UQPm5mnJ5fuCduKKFBKsIjs87D3zEvaYg10D
JMC4wPLmTnJn63p/8UVQ0L0EVjE+1R+OEA49qSZCwDQs8uiUI2fvuFd+/dR6lgqn
1pMplbTK9dPqzsNV46BsXKVH8dL2kawloGceBdCf8eHyKA4It/GgTgFvKy4hqRMv
xick7qwAJ05dz7WnqnV3Y/9OoF/A0P7r34XU2StpSWen7/AELLa0XvknOBc/THHy
7H+tjEiZB3IeiKgDzaf7wEIUinVuoqywKLdJJxNfsVGxydM50XZzwuqe4UFt67z4
k4ksX/LQIxoxQGcyIQbfP9i5mSYe7bZw7QsdzQUd3VmNgRWdqZMCIUTfOLigUlQL
K41/wcWXtQUlar+gj6mfthssmTQgmPgi59RVzyjJspJbPzEUHGWLHsqlO/8J+lZY
TJNUK5c+VFofhQXkhxNNbY2BDSORacfDlok9/SxuzAMddvA49Dp5t5WxP3dFnkSH
bbSP3yAjKs7G2VI+3PE9C7czmOFleCdCBYmBH56CAhr6eC6BKkWdqgMxu6dT9W6B
LTg8iDg3O2DWGprFoDzn+/xdRtf9CbNem6WjgEYv7cEIzQwVzctMe0Z/Meutgacm
OX+KEwOfSTx/dGPzqPzzXMl/Hg9xjjsUyNK0cqctKYiMMFt8Hf4Vielhib+rX9FH
QoDZVyZ8noKREMRpJH3JQE4w3iFOmNqcc6CWy/GofKuT1IBV3ntBE9vcYRD5H49f
7xLC/2JgFv5MgcWJMTgSMT8GdTU6i5G+QoAVfwLc3ORjzNqNP0dwzzOaFzaV8SQa
9BZjZ9hOsT1ryt+3ShmjHnBO2Cp+JjGtmsyR1lYX4AOcA0W86thzQ7pMhUNw/ArM
Y5ikejkkKGF+x0InI0Gh9l3yjxV3R5oHYgAz61EihgNR7DqA0t+Fkbjx54PIzTcM
El3MU9zM4u5k/MWGtuLwXQYQMpcjNHtif2CvFeEjrO078LnzAISTLtzYZ7PX0k1s
bwi9eQZ2ATeMj1gduXd3NIsYsKex+fx5GXcGr+yRm/i0iAjsEERVsA/X9N5l2cLG
J9r2B6OGkYs3BgcCqEd2esQheXVZFbGQXsJBPOqZFwHCcqcWToTgIQY3GMfARvVD
EL14LUEFeHXUZcbZMuvFCqq3piXFMEsdX5LKXMX5dpiA1kTry/aDqVCnBHhaR1lD
LRowbDcVvMIqcJ8/Y7JhtTxPaOAxf3CGXoTpxW1FtffQMyVH7UN4uZwNB89DAiK6
eHdoCOXurfeqrYpiE3vpusfT93XHotSZf7QeO6B8rHVVNMX8FloAjNnhiQKO6/fA
+Csd79dpwbxcDRTfzKnXIPZErbo6lFwSnD5bxnl7opuSlEV/0A057DiUF44kkPVJ
skQMocaV4+ts9TmZHUSrkr6kl0JgWkbXhFEYEuilaraGa9JJLXPER5jzxMIqQ0X7
KXrvrXY4by93M0e7FfoX+cyZbjQQ3Y/0KYjRcO8X6oxZqliXN+8mtZ7hZA4vqw7Y
Z2yox8lo5E5emjrTQnjoXYejR01WFC6L4nlH6CPOoSafsRwoASOmqZQDYuzZpqc7
cJiYc+Tt5/MZHqdjRKVWxOf6ssEsTVgwuZiZS0h/6qLcqoNstH2uNK9/oviyqo4E
StRbU+r5h9pXo6tK9iKG9XYyHQGKBPDRP8if4EsQhYAWKhZ3c/R8RmJvEuuhi/TM
2Im/aPMRAEQf6uj7WX6fO24eQX5UdLcKbVeYs6iTsjUIuL6/+evAaUnp1qyRyDOo
1VnJPa8FRVtZF6IZwR2gEOB2Af7UNj/5pB26ER3g5mMvMt30a9lNfvVXk+Z4hidX
cEXEQlPYh7EG2idIWM6SHdpR7ngzKWLr3e+hpiHgGsIdhD4rD4F+PAVwW56cUzdv
fcfwnfz+YckUGj9d6WUqaJ1UrkEXZtB192Kz1PEad1TtrwX1VoCKLEuJoGXNQPec
HpYGYwpHLp49qoMG1ZGulV9mA1evlCAGPJ3Vs7Duo+QwsGTrFmiPGgIVHFJwF7mA
32Z4cKWOxkvH8WwMgCvyN01L1k7TP8N7SGei7mXSPViLeDDxsBHWFmzS0DMWdSBo
Zfk5wKJfwv/ikcp7ow1Tp82ZC8EP3tEc1dY6qSsX9i32qY5ad8jvKD69EcUT/jD+
Srtk8lPwBWWvHLlc0WfRFbdh8mBKNOf2mYamAALTNPDouasohci9NkdGiyOS8EGO
Ji6MXygbuqFy6nlnUUQAARvlTY2JJd0/OEIZMRNvxOkOztl9vl27bC6wy4m/dN4y
wcFz6Ep63CW7hBrQEIn6uLR+vmJ0WLJZoE3wKlwIXQyCsI3lZCO6+IjzW9Ov+/pC
L1cSxCHCL5zDPykPbapZdL/3+ew4dcL7HzEafYx2MZgCeueLsXCpLRuNyrfWwqtp
sLEUKoAO08s41n737aoDTi8geWu8h+QcZouFOPoIz4yN4wAq43G+u5U94JDr8FRT
WsSc9YqWI6s8R6ZLkvBGgwVhfokFf+ZG2FZiPBApsa+ar1qWCaV2e1pGTmu/wHHx
hfKcKCepA71qFiGHkOQcvprwWXCG9ufL5f72RjoejWKvguUhpz+LqKMf7Sk0X4rl
XlSwX21AM1KQFI7ScDHP7mrCVAcJ1/69303HDC4p0i42k7qYrtsJwUUXe510GJxg
KzBV3yJNv3wI8WegWUQs4piUrv/xKtTHymO/k0ju+FydxWYrokiPkPndGgEF/j4q
0wpGq5l4Kq5+F6zXsshL/3XhisiKZWw+Tlfg0YIVKhc3LWUVQy+eDVmU7M0lwoGz
n+7LhB18kFRpTGOGBxgAcWwFfzI5vj6bl414wLhbgPeN1Wat5dE6IwC18meAANfS
NXxDO1zbmREyWktzUWJc9UF2KR+Hdp8bRoijZHmQIj6Yj0BYlNSruKMiyJEk7kkB
ux1DRiVZLYckp2XGhdozigc6uH1ukGD8CO8bmp8ky3W0B/OCdV3hzv8HN8L4zopy
z5stU471q+YfP1VbSfbSLSAB2L2Mk8LwWAxNV+i4DPyw7lxfuqJ41YdAjKOC3YNl
VEr1TO0aS6OW9IkGUuCf1nfxvJLY76M0yK2G15WggxfJQ1QO1GPkcpp1zg0uLrX7
LwTMUHGvxdIVyjFslHivmzdIhadIQRZmCzKnzkQdC+Hvmn0f5qhBHpER1WhAFapl
Q71MXA11IzPHD//9m6xCpeNwlymv+MLYl+plMq/wpx7hfuijJ9f/DmFdawoiI3vv
X8L8O3RcDAJUZGEUdCAXwc44T2I4LnXFjXsVijvQB2smETu7bzZXOOtEUNmNZJwz
fI2IbLpFwWlVwNNEUbE2tWsoO173OR802EkHc9fBJy8H8hciSUTvvTKJ261AADux
vKmLwXzivH3M8fQxOaU2Ze/mqAlzFhqkzxOJD1tYnnCMaW/NeONk/HojZ6yJn5UN
u+CzsoAWMhWhK6EhLtrNEoyuakXiK5tremfR3EXicF0mk3yx4EKk1i9xNaGyDCYM
r+bJBRzXFAnlWcnqWhgXprBXXetyQPfVlgrB2H/jrDmk2j/xKBx/dOawYwOHn65R
FAYBMBh5sbNseyHZ4OIBWW90mDi0k3hKyonlvoitYyXu9vvhE/yQ8aR7rJm63P8F
hhE8fMrt1KWXHwiXJkpY1z0JcxnlxRkTbAY65tyIvoUBB64qPAaa4xY61u3unPyM
YZoLq4aF38j85jFQ5NXWnFkjP8c1O2FOpokMxcpTjaqmpDLk/yCi+nofXQpAucB/
KRCpOdi746JlMJd0Irg1rWxHQOnmKtNA/mK6Ns7w43AjpWRzORxGHj46ZwtJBKcc
oKlK92Q26/09zhQbv9JXYlwdA1rWNIY8Nhvr5/oViw7js96W30lxToJTUAZhgaHw
wrtpYVY4f84ahJTtSLtCaB/jx88ih+r1KimLLQi0GtWJAj45fCoiHnY+UrvvJnoc
6Hc+X/Z1SxXVpLF+xVVV/M/5jDcvPGsmONRp+E84ypRALFcRUed6FZ6pOFtOiAoo
6o46IAL4wigLdnFHpOJb5lNzM0s5dAQM5sY0cLKzY17R/HjQHQNXmQtCMOvacMjG
WL456S0UUP/wnlx0Rb35QqYgBGBouR/pcafh0MkzmoGPmanuEsXUHLwB9kdmn8ae
dqwxDtaz0LfxrADTOF+h1gL0MiXLoBPiX0etP32g+Q+UtqpKpKZ0tHLPQtVavags
DH+FMv1Na9/+3OLK9BNtv8ERjoSVcseOB+SQHmNi+Tscs03pnwId2WVUQwZt2LC9
9ZTOJZxuKar4dbwYxIMrrIcP/ZTPLek1hFOjrgNurXr/ncJvW1Fcr+N2s01k4dmd
qOWUOf7zdi6dKenE7UiGZVpIpkp1IDdzANZvz+PKUDXSUL0wluodvWEe1ETvTL6i
t9YsMd/TySArK4xGxTf8r0AMTRWkaif8LvYXB6bEUIb88TnRihR92Sl31yqvrdTY
uuvVc+k+mRnLLAN30V35iW6/68ao9QzF3I/49gV6PqZmkyfRPb0Xk33BAEU0KK92
EikxWBh28zTTS0gz+WtLeav9mctZwm+8IzlGoXwWNhQwL23J3FzXje77YTYhcZOC
Zk8RxoG/RmGyREarF/DZ7V9BkTHqKuCCfJXNn89z0hh1w7f7BKRuHcmSwSvSkB+j
MlYq0J4pWZ+M3r0jgpnMMjLf7chpWVYiogpqH/EKaWcVsnNiDimRqHqsDXB6r5xM
2y65WE8o3SX7RV0cwGyZyaa9gE8Lhb5pqV9LZmK8eq7Qrc1oi69Wz4lseE1/60eK
9n/29+2WbQpnefvj4xOrFWH15UAVe7sxYxFNR4jgSxxtMkfevWHqbislURATsCub
tv9qf08rtGEelJD4JB0p1IPafiAU0imxFDMxTF6jQKZfxV3+zpXS52QdAm2ZjLuS
mTb1dTirSZJ0Mp9i5p57zM7MzRBXQLjngwElsZFRLogLLyY7N1Ua5bFOnYjSktP4
bfNDIjVzoxlUDWr7TgDs97Yt0yg8PBAQiH74cYq6ucwyn7qLwGVv1SezG9TGyt06
yVztGei8pjlhtvz6WsAI2kceHSqZC6r0NNLqO3I2ELLhEwfUPdVVoF5mK66FQVKv
xOEsXDuipRGyqrilwCXK7OPqRUI2LESetqRK+vtwk6bHg3VO4HkIjJYcYCgZzKTV
qqqj/A/jeQb6NglM3JHRCdFzgLiQMsjPm6+oaia0OsrmENfPIet1E/gUE/FHWI/Q
ihwq+PM0uvgWYdL6bSS3WpOVsDA0ZN21Ww3k/M5D1g75mfkCY0RfIKlt0mXqbZ9g
7mVougY2emE2Z2vxPNGZrdKOMLZp8eT635ZrakrnK8EtFzguxxFs8hXghpcjE7Ak
SRAZpwKn5aAkJOhcaqVu5DChTX9sAWajEvQTJ0kQQhvA1Pccq2KrkV7omRg+rzqG
WCnZX/dEJ+K+nTPumSFKjn0tD8FZUSVDOcr1Bkc1u43t2kV5cK+GdltHgGbqF19A
FLUa/j7g1+kicKGOphXv/xzb/Vo4PFgR8OW9qyllvLt+gHapJZAZs5r50+0aw51j
y9FQ0nreDpfH6kqluo1Zl1lwaCsO5vhcJN9+bcuO5qU7AEgSjAiYuw8vwpEoerTg
Y7kd1d+9S8jvW2LXPo/iUPrgIPWwL3Da+/wZNL6G11iW3feybED1tngGvhhMyoiQ
j0/CTx494DVfESSv66L4LyHQrrg/MeJ5Ydi2ZgNISoFR1pSGwxwsqWcKeK6Rk/1w
NsolIXPM3BEWakgmbj6lL+QtvEimPLazJhDDy7axCALMs0BEfEpio+nrFcgVTBVL
WaBMb5KqLPu4EBDE1hG2/ubO+ALkTYA1boAPER9itc+SadJTpZqQ2AsT0FdLHLq1
sBW78MfuDEd1fwg6axEDHsmYhQfb2HLj59jMDFFRnGJyYiDr51SrZFPq8KhWPnWs
aKRcYPYOaLeyfJuSgOaTbzuCSHbKzMxBVyIsXue5908fi9V5U5fOzs2HQ+fA8sg9
V+41gaMO+AzIbTzGu5re8cQZVtV6sv9uwgHZy8xQ9PGhKiwcRDnm5mq1xzGBkSYo
hlEDlHLID0pEAUpvkhT1eqriXQyjYvsVjb9fvCbYI80+pMqXLpHfMaTlaYb6Vtkq
qK4YPW+gIUTRy/6EFkCkb9HpRSzU7imevOr63NT7/m+XGONkQtYAeTl8y//1Pjh3
xd2/QTRu4ZqIByWr8IKT75Q5A/Mbcyp3Mo3UCvFMmrsG/6wT9cv54B6VL95n95BE
1wskNeF5bM5HYh2FoFjko+kjFzCXRC2+iw7KyzJRGyumKJiqTRItKo4F3srD5E+y
ezsxQOLF6GJBCdNoLwsWOeKpvbmDtvG7ifVgS7kLVMHMZqbgobOJRsDisTmtVGWv
C4Kl8JvOK3cP+1Qu3i6V0IcdyoRoNGQC7YkFm7u2Ers1uTyT1IgubWrtTzdjKGWW
7BgO8FEhTwe2BL112lYVVq36LwTvaPuQazrsJ1HTWAf64r7Nz6WG6+tJvm7VYoWG
DG16RVdfb7zcjTGE9cnjQCh6JRgazSDcB6nFu/FJB8aWPjHBGNnUUZfLh2Wo/vqu
hQlyv85S2XfcZFop08T07CRwvpnDCPZG0CPvDC3i//SLJbGtooSItER3GYUA+9OT
N6jRJcfYUDITcAKrX3/y8SpZpBKvlJrGL7XUNKeM06LE4NjbpWsagBRnY67BQB+N
0+8Zwb3NTEbgTzpKwKUa6/U0j/XS/HAf2sKfyAoE9dJKU/tr41K6z8fFlmtsHT8k
80qS+l/Uof/ODEUZIE24Lb3zo/Qd80wUUAwvuxPj3nKbGhpc5BUyiLqFsDzPQRiS
lJ9obdKhedql9akdtsdtV/+h9qEzFGmiLFGJFcSXLEuA9gthlqWqGQ6E3XLHaxSB
PQXNRDX8hzvS0hfC2r1zEIqkvxbV6lVOSmZPWqj8nxUDA3CIRmMVnfMGDczHQShz
sK4i81w0obJ/sq8LMG8FvGQj+N5THrlBV7ZbYFXqIQtXWI6pHGcLHfx/1u6BuM6x
R277cNDNGwBgaDagGsdgwj8Fd2cFWyqJiHoNsfLAwT3dBjRbWsGpXk1ROmJWFhDS
DXFUHYBjhq3Hxrh3UgePBiX3Qkl+hkFLB+drGBDcc7ReeG/HKKE7mswXpWYS4lCw
NDQxjhzntO63QCdTc1c6IDKOLC1ZeOKeAquU1LYoa2pPOpLSxhhveflgc4wMAmXB
RAMBP+GXwh44uOouwE9XDFbQVJ3kF9HDZ5Re2A9SaCjZVoAbtSxe4Q8iqEaKoyea
h9KGHEkqF8S4+PiVNUqzYgvqUpql8YsRyc+xSHZpBh5ephQqNTjOekPFJ5VmmXq4
doclS20wzSFtAFiMXm1RqaYOpO/JAqDSXym0B2aTWxYVuU5xIZI0hhX6SS2+H/1E
WaKpVKvMHKlKreH5MKZldbtfbF72yE8RubEAU9tAOhQ3KRKta3SpzgirNuuSKnhg
lDtpDdyEptAuUNPWr3GwViC8r4fNoFjfdYvz+BuJeFgHGyvxFoB0GHsNgOjbf6vr
L6zf6kJceR7MFLb39pgxmv208+KqTbBif2oJabdSbGcAfpSOpeXfOmADfGN65AzU
QptsYr89fA8RWzbXmbsMvlYZNgUHGSUW3CJ++KrXuf0x2dQhEAnlelJpW6h9pMx5
9r8oNNdK/scrZmQKnhT7vVz7Mzt5Kk5RKxrnh2/vWVtTQ4rXhea8fxLfglI9DC2Q
ILydLdFPf+YwBtd1j8GMhTJlS4slDlr5YPOnk4tAqSch47FdWrYx3dfIcEGHuZ+c
3fo7yPI+5/HmijqhggxXHTb9giR4V5MMwbSXHZgqqW0lKUXFN71aD9mxSwGYB+G7
gksXta4impkcgAoAvkGLuPtyAkY/PmF8i3ycd27v8HS1RqDtH3bcsqIvsu0xkwo0
YXsTkyQdgGKS6SqemFf8CYBcnAHqpeVSd/5GtymbLX7OefwbRQDn8nleJvvH5NgE
2TVyRDX1SxJcn6IzMwMIwceTOTPO6se0SvJsIS+2cMwOdCCQfuUheey4k76B4YgE
vftdTcc2HibILRHuyt441tALLDSSthoMpvvCpUzIIKE0tRMk9C0aFbB2ATiW9oOS
fPkfG7St2+rSzUQuiQkeMspQKqFR6xop4hztchZod7yOzoh4qvpeOZQhQNox1asc
n+3HWfIXjvLKcerqPknpL1JyKaMIYQsg/w3xpHl1dIMmeLOXZ8d6qxDISBMjLS04
1Oal9jSY8L/3r66zmjd9xVpukRjEkduOhHQ+Y99Uq1mZnuvJ5/YBM4ruDiNCPG1p
kw4ZfefpyxcFlybrzJB/vhRG4ajentPiaJcb/bHP6cL/6iedhERiwzT6m2ewWfUu
eTx4hWCEb+JCiSRax85ifsbvG/qJACKZNChyDHs+/aTd4TMQxMwEl7iBbPV6CHqC
wX5I5CBMhRvfZWlYnEO/aO79SyDSZ3GdWyI7ab9kzWSFOtb7t2nDDZ/cNw9yis1F
ElvUvk3DZw2DIsAUKOUX0OnPrEOApr/z6NY1Vqtfc5oVl3mwroD5ZBYTUk94WqtX
sVSd3YgDiYPSDLIo+5hQnhRmOhNVBcrtFT4gF50oivnT2PBci/FuEZ+iAdZB856e
Dz4hGOAtIiISi4j9PTWBzAspwBbpVlm3qw4SD2JALWDIemdKf3otmsCz5NdC8WBe
AQ+MgUztF+GfFq5iNQh2aAlVfdNgiFk91YZi94goSVl6GvilMmO65JchffQWupd5
D8ZilsV+9dMIhBXZimLV+TNPyGcb6D7uG9pLWadg41cW2SNgz3ipORF7PmYJaRD1
zp6o4RlFJNn+G0wWobW0b2neMC6ZljDhbEqI7g5UONtcZ4+T5N/GKuNrDXUbLViv
7cjhsNZRdcFbzpSUSikl5xoywlQmqpJGe0KZZmv+b/tGfpI+UPRzFheyk35+PQ6Y
1qOdEdIvYlh+1mQLew9nx1jpPhrPvgBSntiRchg/jFici/mNNmO4aqLpwr2mUI2R
bTlKZa0vgfZRpxWU2vznIKTzdjrbk7277ZzjDp8F1umupQ5hOCi3ZSmlOFkLnKsd
4g+QXgYJf2AfpwTpSOGC/PS07a1XzheT39Z1g04jMjRwUajq1lyeKK9cO+z5BIMi
uTeXEmOk2aRkNcdzEvr1cgi8SHRK0FV2a/YHl5PFlRI2Y2nMGa/UoaENO1ahH1dy
xTZB9PxphYmi1PTrNsYlBUE2VCM2GMMTNPOhCT6zWclxHk1thHzvu4qnYM76pMxD
k7VQG+CraxAAMS50G1xaKgbNzGDWkByJyogVXkgVdDVhrZJf1Iqodd5GJrG9++iI
2JICEMyKenYbpG7Oa/nOAAYtCX39fkmh67zZnauLkLSJy5uptgNjIjJkJKZJMpbg
RVbecLa+VHtZUO2IM8L+ufqxoI+nhej0uR2/Ax8J1ryuVjzJYla6/aCwwkevx9a4
wRoJ1r1G6Bq9kOYTMlM2bM7juGA5IAevsuF3yXJUJWIoM3hN9icBP8t9dNMaWlvs
2MdhJLuCEbHYF156xUo4LnZjLPMavNec7txEcTVJm529bm5nNpRe93/Fl8P2ys/L
UDqvAwxBNjOSRLPpNMuyyF1m2uI5mKyUCeGYYT7CP/KVosphDk+tecr+isOp97Ip
PY+DRRNF4q5F3uKglorhDAPfufwjrVbk7MwMA2lhlN7+9qOlzAC54obKSgkrMW6j
mSITegSZ7wYbGcZ1oFJXNumUiN2/EuCgX6TOfG4SQZLjeMcdojwMHH0VJbDV2tA8
PP9Jug4jZCsK4B4A/zsvZm/5Q5OlElqDZh75Bz9QVesbZuKoAir+8tBIL6MWYjPU
9mu/SYdUCIEeSYXUzLOdCL0GN5rjCqs4lHkvvn5myNdyV0pGFAJzqC9sIFERbcOp
b/yIp9lI8iaIsqp2q5J1NcnwlVpStIRVdUGB6GNQFCRaPDQ5InNC/QAihZQr+/Qo
qZEKmrBTEyF8ErsTurQJu/46riYdE0s6lkyqd3o6DiSJEciA4nQiZOokhqof49dx
aCRSy4UhXYzZFakWLCsA9LTXJTk2Ysxu98DY2a6BrRz6PGEumMw2ZImsOyLGXfjU
zNISiU6Xuq+63vRfOJyS6LPcz6wdTcHqV9DGwBD+QXkJ0RNp8RRpdtkfuREDNPqX
J/1Pb7yYh2jeW/zvwmSDO9eZXSKb8Adb6zpnm9eDRxy9Kl4sWVgTSt8LM8fP7Uza
bSjO5XSt7q9bNNTft/oxF5nix4t57F8HBrqE5WLFzCBsUYkGsHki+nllrBGHBSUQ
D8/b+JUpq/Qrsp6xV1w2D0qOWW2esw8rO+GFE0WwZjREeeCULfSVSeIAThc87eu+
FKDhKsR/NCScc5Qt0sb9R5hiG54yOpznDWvBJqBo9VWqO3XsyqM6eUxop6Yd1yzZ
eBzwjKuMJXLmgbBudf2bQlG8wKUy5TUiSORu1RgKLLmXQaLrX/H2OOjEskYf70eW
lPWH2r1PvPiD6aZIqj9elLplEWGKGkCayfAthYXcfX9bdD7EUN6shkp6VRelIwLp
wbFyMhMjXEagWqBo2s89lepHelamE7GCGw8gQcttCll5NFBs/U+ov1k5oyNplaZ6
14+JdVOdSZsJMVnXpdlpL+Cy+SZQzM5GCN4Dglo+qLltPRx/dG/vE1B1tWm7SZWL
TM226XTjAlZAIMce6vzaA5rCZR5XePHqZ58/bZsb139shH6pUCebQ6VmF5rFbpo4
sYYI1703FXDYhbNXaHiyrlyLDa8kJSZ7QZDA+jGHWslfVMYEmmRob+i4Qsa1+++7
vkMNDSitcH6qYxQtlGkXBRn74PyzpzK0+qh86Ii/prUXBIBTlYvvFOsKvmfv3n8f
WY+J4Gz6fathmnpke6dqX+vqC9VGPfoUfbhmpvvBYFVwIM9pJXRCqsZTf+psJaUk
B/ozynQfEaFpgjUHw1kmUpGDDPBMcrxbIaOrWfr5NmF+MTyJLMCL4uAvIGMGWWYQ
qAQUSeAlnsVBhkjzACPNdMo1ZaNKPJaruOkE/h/hOZFKixW6twToCXJv+brcHoi+
r4S66BUyTnf4UXjviy9SWlcJ6lWZwL93A4e3+fEm5+22sAnP9nQiKzdhhJXbQYyA
YbWqoHd/oYlIr7j6s3He4hJahiFSy5bvWScSyIp5Ir/0O2rtLMh8qxCtwG1jDh01
zUVOCAMqKDFedjfmVlL+8OX2w8PbHN1Jd8nR7U6T9dfAZin1JbxKwWCahp98LRsF
FqgPEeIMGhZpjYFTFORpnCIbYveFqGmw4K874CyLgDDjF6mQaZAjrvCFR03mqdFd
HhaULvhD1CUUsyOWrqJaI7OjU6GUDUhBHWfSAGD2RGfh9fHrRGR+LobUX5GhAqZX
4xEljnoHFrU1nVC3lT73qColdCrS513fAcvmcR1NoeA1PjZyl2rIU/xvda97nkGH
UwwL8kpbGIg4hvS83MBnWtr1OcRhv9HRe3UHQh9mGC+7jXiHpB+1oQ6Ph5N2W+8Z
JoZKVJiSlD2n0qm4GLzqnf7g4fp4LNPMgmK0Klp2CCV7rPGs6sue2KFLwitYGw3v
aRbnV4Ain+sKjwC/7kJbhyW33RDYybrLUmC4IyGDPHHfkMlCP+PuK/7fTuXuRgYQ
nJiZYHzQTj5hBcs2bMadTaWYlN6h835gMHXA5YJ9bSnLmudeh4UWcjhMCKcTU3hS
M8xdY33asNvLpDa9OBPe6BGsfrXFPcPqKOya50lTpEvuBNAQ6jqXe9rWaY9MCPui
Ikt+plpEN4EXwqscSM4sxxjtQB06zVO2CP0ZWe1NJ4zr59d0qG4aZ9HBoaG2ssyY
sHxpFwwhsiHDBaWCOOyrCOsXktZBet7Nx3CzWl/hGHUzdVEd1A+Yw/4F3Lw0PzJp
JB8HZeaVUGzaW9mgd6UbCjXWDEFFDVIK+0nDgg5ACf6GdeWQU0MhuVeRMtlKXJb1
bbS0KOyfYj5XUZIOcmAJXhYhJAlNEF2jA1zDB2m7D/4t9U0gPiz8k2glq7odeTOq
A/Q5GXRwKwDSChWPtYhiG/pPekdwuB6xBx5xo3/dpxGPf/XpmWLmBcpfqE/eSvpP
FuUy56+mEEnPQkaC6BxRhVuQ+VdjH5tEziPjrzEkM4tFyhS9JDKOJNoagC2NKV3l
TYUOTLCKsMz3b/Y7lNaAtgimiZRf1eaCx4XPOdCcFOY8UMWUTDWVrzoK0CWpwc4d
VXrb9Y2RlyknahKmU8vnB5xebFqrb0AjWXnXN7OtBE+cmbvHED9ZFWAAkH5WE6+j
TOQ6IBNkWDM9AowNrlIQqwXPRlMk27+RAvs95EzODoolzwHCKAGG9blwwyLOfbbT
f7ZaX4a1bng3go7ba/BQi6fZsQiBthVsdtgMqiSVEX/g3KYhQpxJZFkstRFJqAHR
CdELIpehjFt9J4/vXVHCxKXWVA921jbl6BiFiD70siOuGiDplxeLqBN0D+6OvG5K
ewrwwToFyhORqDBWayyJ1HoWf+8vWIdMrdLjJPhtwnY0jQoLwuZ7JYsvC7Ueus9I
AK9TRoiXhRZAgCjq7PUNEeP1WcUjpvmPPRlu+GfNnni+CGZMeu4lVB3S8isxWS9W
an83HnGGi16/S7qiC23Cm3W9iwJCoeEpuATwcZZ2W5QSnZtoB8OlVYylnf6GLDn6
KOO4DpZV/eIVjMkO1N8VjCAeYB8JBli6ELwAeqve1UeQDlHmo7P4yMZ55vwKk2mb
hjj3T7zolns2Ai2zNk1v0891C10nuW6PG9lhP8zsBDG6BhzI6+6Oeozua0uxF9B9
V2W9mBflEal8lRMCFLnQ9SQijTyer1w/ZLb7b5rW8QH7BInKQFF+ak8mghcCa2+n
n2/TJ6WP918s8R45XzWyTNQffsn27vDMlAtJHRXv/CnrIoWVFC2VpvVG+VNjg5Lb
GxZFrfcDGHjJTRsTh4M9cpGW6fYYVNkOQ9rYhnD+krmOlrNVHl/keJlzbGj6amrC
RpdVGgciDpFHyoOjwCtz+J0R2u/drg/5Xdj3ALu8N3qcZdiD9eXaeERmiS2XORFD
ZlUQqpf2c+jMVQmnRfNl4F9Y9cfHMA0gbxP5sEqQq/1bDxAw0s8OqJz5AUoDxIJO
XWIEbJVqMpVyfFrnd8+2zzSNo3nPRb1bn33rSz8TmM2mRwvnmLiAcq6Yz+xZI6Nf
eeiQZk8lxLszlUCWFsBuJFHcdP7SnqpYXQBnRWX3PIhJ2t/VEK50XVCJ0PFvtz3G
oJ2TDlrDLgjtJtjLqh0iWWtDtH5QUKRc67u+7aNT3IJkq/GmReTVXpufjvN6LAd4
VMGOZ7qZwgpY8Qd9coPtYWzd46JRz+cHaMKKd3JT67S/Wh6tN6a1IJs2C+XmNlSQ
K+t1xJujuCzLIhOkgd8wWaByoHDHD3jd1xtAbA3yDxFeicLdoG/e/2V7D4IoB1dY
gi1/7joQ2LzPTTH0/E9aRHgTtpTge4D0442WK8vQ0CJs/1rpPmBLBnDCe1wGCshM
Bm4kcMUq8cuZ6p0bhmGxmlZnl4/QRieMGM39Qi6imNsLBGH3G4KQBjkPrDC+VXQE
kpwmnAkNmbOqGwjUaRxElcB4jzjPq9HQvDXRXLOOzlV18nh1c8USMTa2uOdFuqvK
gsTC/JWbnZVcoJJf8JU+qnZ6CKF7AP0iiYKY7D4pVNXjCNZWJNX+vFo4NVtmqQp/
5L1HjRmqSu99Qg/TPwLY6pHvqP+KJmN7kX/8ZD1UACPk4OTUXbAQr+zMagP2ncG+
4egW0BZOZmCBGGczp6Tnzn+C8gSXVOeB64u/ISRzrBus3E0turjCd34qhupF7n6d
MPVRAMoQVAmEf/YgPxHCXqtVKxf6JSuN9cRjCFgTjLMcLUeG9MoKYw0JxyBFNpY5
y3WEZs8all8TZEa6/ICMd/13ZHJIDQZTdy3E5lRIk3jSOjSCqT/4hAjKvsb7Fnlx
YrwHkzWikYixxyvaRsjd/VlaBmhEl74fo3MYDWEEx58gtK/63r3/w0aJfFgw95WM
l4AGoI7ZaVSQD2Di9Tg1NiROCO1h0M15F9i+j5l2A1xdtisAuiPVDTB1QyyUC4pC
JLHlHFqPZZbmRUv0Ef5iyTM1y4rzuJZYdwiS4aI7qUCis/BIt9JBUjrjDpVf4yWp
74eAmw7oVT5aUGsCFrF5lPjvFUh53AXsAQLnBMtXEDxgciaPFUxKrEtLjmvXnZ5j
JQTCDz7coU4HEoAD2/DdUrmREOGL2dGN5UmFDGEwfbSic31XTVnt76qZBZ88Mo+Y
HzXxrc6MoGjET/7A9V/iSBzw95lnnlPPg2/eEMQ1lClv4RLeEQief94uMFBQgsRf
xE2NyqAMA5eXPw6pXqlZMRSJMszlts7H7UbCANi2VbKZc8ABu/wcOB8hE+aS2Mal
xb3v5yh6nXJe6KrPoN5VcyE4Bzo0PqHddQty+HoYiKuQjfjYvgcAu15SQoWsu9EG
HrD5H8bWhD70p9raUxAWLO8GsQW2moPnRkWoPj9xyXaQUAs7BVczSRkdYKTdjdbK
Y1bzivQt0XsZRrI9mrZmGmoAE5sr28jmNKKWs4SNJ7Qu0eON2t1Wd8V2OMR2dvfD
1fUG4+Iw/CjNAyI8PTPRq3/Bmy8Zf8H4BqOnQ+YnMJSHALv/NfFUk4F0tsFjIbI8
djZh9dHE6CcgfOOGnf39tL9Do1tnUwlk6lMl63UaqGySQrUdq7Ss5Km8Ys0W2wkq
WiGV8hfZNPs63EUbOflVLf+ZiobOmQpgE75kkbILmKmnUPUsGy8OvvRx8RpQKJOl
y42tjjc9xMnsML0Ofwd8tIe4c890rMpEm67YqywRji1CuMVFKQcU5nT3/PuBGSrM
XE2lwa2V7Vnlj7NGeriJmOvNfT1h6YAx9eVBjuPxqMFNZuCAT+jSRUSnp0p3pvLA
QIVjCxGnsmbF36V+aM+N/FCOnKZrKBjtA0z5Qo/EVuc36bWiLCA0/Tt+QjeT36mG
ad/9GtUDS4o7NRssla+9KdB7OlCfupVwFl4abrIGwuCAgoJOsBrEv3/yfhWUmAhL
MzJPdVbz1hBldXxU8+ztUXhBi/Yh00qGJio082kKWmPxyzzrfu98hSculiMrzEex
U3jD0hKQVz/myUS8Go3sFhRpkqFimkTHdtl5FBoOZW2OnCXeE1lJKTgrs+mavkFU
6qiyj00CvsbrMp3TyuWfz+PIlEbGemnI7EDb37Lp0wyWnXoL5l0urhbuh8UV5ZG5
h1JicLcHVOXAq/RVdti8SukfJfsXVhZbEcsyvN89t1Ck1u40mZYCEEXt/rzQr9wC
+qkpK0p1E0UVgdnkhzDqgvbhCdjkYGx/BCelH729gpCJBzDg/bjgVkmh4xC/zeuV
Ftrj1tsGsKGTe4xHhnQVa477+l2IyBbZHbHvZIW+OWPodKoHVk6a8GpmoX7Wxqrk
XaoD6le+YtmKpQipPNdzRaKEoqKtBDnU6hC+ZjVipIPs7tvmUh0d/Y7hqMNSqc0+
igpdGSMbzxPly6caBla0Bki3ggmcHhQvTRkdsIMrmugpW3HjbA1CJ06CZoagLUzk
Ttd7mJtlMxFb/s/p2Y2sM2zIOFSK2O4uzLVRSVN2mFFUUo5Uu579cGGh7lxiVxv0
RXV6Ew7aOgjq2ldipgr8FJ3Cjf2OOOZh1bn4s3cmHPY4fGCpR4dFBAgr3cc1+zvx
Wg5ZAUvSEpOeO8Hk1K8kEuh/QAeLUt3z4oL35cna/6no6MagWLL7OoZTBUeRBcd4
uilfz/kII+EPUhKX+yftnDgplnm+4Uwk/MvAXKATR0DD0WWUMzIU/kyljB4asUkl
ws0Q1KK3fp8pXo7hpF72yGC+JcqGtm5RBy5oDTucO514qmaUHC492NGzqrc8Kwyi
v1jYMf4Z+CeVtU3q1p+ixblvzShKOB955FTCl/dmHlQFeF25lMz8Xtu45KyRrrYb
nvmgyQiGwlpsJdKp01mfJJf+h9fquHIhabJ/c5LFXvrb06qGuoVYx/gPVooSyTRR
1UXJDLNPDLaV3EQVMfOQcZ8UkVfRryCpUvJ2CtNTQp1AX9vy7aCPM7sVIAjllps3
d3PIquipkUyJX8IUP/MedynRkANo0LVe+Mp8fpbAiO7g3PHiggPra7sn4FsxRzO1
DyeiVibBNcWgoIfqH881KAl2YtU9+LrlKAjD/OHkvH9nTxidy1pIlT8n0+6ptWcU
pvAu+mbf7cZEYNTjeP+5fUOkMfE6zo9dNfTK3DyVYnyyZuw0Z8u8n6EElmLUHy94
3WJTH9++kqwokRS421oC+XRIOocljjsz1Ujd52tj32pQSYsrTMMdbzWJipoxyj/j
eTvLjRIC3a8FrZwGZiYjE28Mpc9K7Xtu4dAAgfcrh0Xiso/e+zXJffhO6lc4wJCH
kHAQOwdWvqyWUr/lZgK4jUOP0YLpl7wtu2qBINT19WbOobwwpDAacASqiRE5ccrJ
nu2fu7Izxhpjy0tAfBY7isrWw4AA4tHWRMTT6iG2YFmQ29yacTMDpZwuOYQKw1wW
mpZfcSngDgIf7ZIQ1eb7kVG/7TzY1sNu/SrEvmGiyLeEYHW1kQMxGXBiCnk5Tave
MvVgMHGci+msC/ZPoWB/qT9yMcTBttp+oSCHWvFjd+LAUvm3YLJwXc3D5HSM5Wmm
j7rHAlUeBnqOPqSQO72vMoaHPsjQHf4drdDqYT7rDG83nV511up79ykWAr9YjPot
7Pa7dmT279rmDYaspabj4vG4Ime+QrwXT5Ywl8umu6dJIO9paS/RROXfyEhFVorQ
0HS/9+8i6JkwdFOjaMwCUo7r8KKYHZ6LTjQod34cKL+183taQ23l7eXnCTjlezKi
q8BxLeAQ0UYUsMFBzmlhlTyE8CoAtliFFCgLo6NnYh5nltA1HxyKYmq/hl+RjUaZ
kZDS9arQxtHUS5Iqq1VeINAUhCy0Eb2pC1HqR/c9qek58mi6Uoe8hVpk4yRNZZqZ
5tAFY1Ta1bCQewzJP0SWkY6l1RPe4bj6hI1p5H2bxAqXUpgevCLsZbSZyqrlsPGb
NVft3gSYiR1JNxkcPDp5kZvXltFKVXZ8s3kT3m/c4vkj2gsYjUD6Omv6m6mRRSXR
dfBgcnUSZzvv+nPdCyV99OdjveiGxs7E5ZhjVSKChs8WMVo3i5JgUSR0yAfdJ2u6
w+Jy/Gj6Um7CbmnN/toxihT3pINOL7ulsJRVDM85ES+Ld+Cnu86epBjLn3LpOXZx
MtH2YCMkp8C6guQx/FjEWxthUUNIDAOdo/tgE+KeNTkaLsGbFL6+Oqt1moIapBJ9
o+ZDAlrHiodiioT2x9UB5ehflO9ljzk+b6zMN2ZP3XaHYRI2V+PUV2LBXcLNGv8i
kztKJFdQhsfUTacTD62tR98jH9kjS2r1wY+KTyYWQUYwrypzaY9FYVHoUAtm6v8/
3ZMIqHqQSFeM2h9D/HYsut9Tv1hiX1wUGLQxnG2gw5IV7ZQLuDG+I0+yB5mekBar
cYX95CuZYfw0FGehhbgKTt4uGRx7LzBRvMqUlRXCQkFIEPYTfN0YidZHnggoiJBS
ys3g/tP5rhr9yGyPnRl0cD6yLCMOj6rngu1+4/E7XjZocFKtsOvepgJDbgEuMrjL
PEyLtATP1xk/hEJLRUul5g+XlJclvI0WMHk+n/+n2zLZdM6aEpDLrauk0wpEosin
XvtUrWk617/PnjN8WtO4kVmAFtPbbAvjCqz3JGWT9MUVNgdVYsAHHiEl9WQ9Rghu
cqA9a7aa0ga1Zd2f0hGXBb/9hkjhKN3jHCeS4vFeuAh/ASIE54EawOUJzftwC7EL
K1AJwC4DW7RL0Uzdl2htzF8FbIfgeu2WH+WKD+GsA7JXaIG+uRf1Dp0f2Afd+A9Q
vDon5U4xQc2CYC6QfsN0NV8a/I2ZMlvm3NPVdcq/dL4YSL5604XatZvqKsXywRLq
NLrUdDUAZaYmS6yvj4OvZi68tAY2utGW4QMgDMhFwizitDdkttG5S3cQAju8lmGd
Czyz1As3ii0anXm7mIfrV7BPVMvatZpcOTR3uMZnfD2qi+reApMe4WmbJfsxSnle
b4VzNDNR41dTmPuPFr8RdVzjtReGgGwBZpEDRm6KFJaRBVISU2YmoF5gCNMsKxpn
WhcnKCufVRtAip+lsXe4WuPykjSpycqoyIIsxnLQUZGD+NlcEXngwCK1fKu8DdKm
wRVbBXmZZdKIA1ZiL5xNk5hfiVyx0mSh28UUtQ4szW/PSWDxVTvYAXUCQ+emXGrS
mvPy+cl/LqJQr94lX3H61hOy/Tu1RawsogiCa/58VPROyDuSBgr2rkyaX+DWxVAM
St9y/pGI2VyE/qxhi4g9OcC+XmSrc2aZzzGau2MZrf1anejyrYWXLB25XOhRxpPA
HN69gcPtkv7WaL41V9v+CzQ5v7xiP+XLw9V9198win+h8QIMpwSRdz+4hNEy+YKo
pbEfy9YkhgB+U4fgXeLWIrpSA2RLi7s3VGrDu6tSB1uoI/n/T2J21118oXJ0CK9V
mH/d/KTBYpQNC+mHihoSu7KxbYvdudDHg87McIdOwQTk5RhmxhAx3cTdPvBRbMaK
TrSNRewQOV/ysqgEvJ3OMCg14h58caCUaj0A0e6IKzAQwFvMyXiXA5XsKaZRXMSw
uK3SaY5NEYMJgA+hP8FyiBNauMdqfRUNvnPKCTuFx2zj1eDQWjo5MMkSCnx+NPLq
T3w9ogCFpFMLU9pYOI3RLM2K31rlGcI3n+xbT50AKIHZeMZsRkaEBhFi9jd915BI
t1KuKmOU80Mux6NQmMLU6QAXdkQ9iNmt3rYbIDwmaDEQZ47fLzaOVfJafAT7xzln
aDpUT9ajD1GZNapuma4C9AoPN5SNbCFHhZZgWVAyhOfizBopmar7PBKyCNB2zcIZ
dn/kxqQZgjmP0xuycUFSon8TceKtvcRi9O6sKlfZu8VCDa3vLt3RImXt5RPaDIJ4
mY+ihiMKMhuHWlIiVgiYOfUM++qVqFBN7CSBALevWKqRMpJTfvwXpfgx4/YDFCe4
fDZyuCSEzAhdnLuImnOmy1f5E8kME5hlzYQ4LZFydYjInzyzt/ipYvvpPX47kvm7
iucjmtRif+96LKNIJIznEYUJv9Lt0xWMkjx6bZqaOUCwuy39VP7WBA059g2ERDdR
bP39xvF8Ko9F8j6fwnB4Z6vR4WapD0TbH1Rq6PqqacGewkfda41G9MwGofNOl4Yu
HePgF1XdNS0SsG/MBA75ztHVBXtMeQfQqZWvrV7tiX9d+7UTyErS6KfpNTuITpEf
r3vr6uNnMogNAAoqZngFkr5BxJYOjiibEbPPGE0g5bNkcp0GR0rP++gmV78UlQNV
QjnkAnfUOcDjAOLZLalTLSxHbFyGGymkYqCeWPuQD7ssg3GSHPDETy+n+ODmgJYt
HMMpRwVRkOTnIpANeTwuZqqFpSxVYJxaaSNgnxH+DopdBszH9bAB79sdvwsKPH7B
tYADutxvFNK+nHCtcJ7JlzZbvSiQF/EY5QGXPceqSCJ6gqVMlO/I/STCrsSO1yyM
b0sIWIEEp1/lt1/zDd+t+JXWG26OsUTk0hefkLZiqpv/8E+zzGs14EiV36mUVAFF
RSZ2Um2UdWjcySWRy/Yi35RQaomqjWJMVBAx/sGHQpJCzHILDKTAnr1mPQjSqDc0
d0NxFrb+Jy9mydvBF+3LknltVZZDKslVprYuYav7ipEPrQxkXging4nICT+04u1W
Sovb+e3zGmbkDhoHRb2yE6kJhsePTos/QmZJmBymvlkqicd+AiCfe7tklEBl41/N
RHUuvOf4LIEKdm7YZEXyb/0ZwT2N8/R1PAyo9+Uq+2sObc9Q4RwLe4otp7ET/Ltj
HO4QD+Sc1aXZf1oKDIccqeE3H3zySqP1Vyl/RqTy047kfwEF0BkTTqau4vbq/VPl
jFWkQXo2TwRB4lLS/ytEXVacMYsF1QX9en/ZMOUDor2QildQXJs0EjioHoSNB2wM
EFVfPKI8vL/r510vr0p+N/bTUD6GP+t/FrIOSQVTIwSc4GWBNIW2bM2n3BPfqaB+
URWKM6507C6jPXOJR4gDqPmqBbUWzqopZSd2VHy1CiP6xnpGoNue75wnE8YFKMDi
Gl0C09jFZ2cMxoATDYVYkYr+A92VLKpf6imA9fI1TVebYFq5DMxil/L8anK9UoWp
X6AnEL6hF4HEEhB16oqyuZXgAS3dyPMcSJA8laTPMkFjfs35w0vB9i3yymimXZEz
4jnNUhloagpkzPwdHq8Lm9n2J6vUMO4IWid1G92dCi07DXQwY1bjis13+AsjzaqK
7kJBX3r6W9YZBMHxyd8Xj+px2Ixd287AnjmUATkH8gDYeQUZRFB5Ho98AU9yM5fR
SQOH1f8F0gNfeh4eG8GhnQtEBrN/oXgn6qsDw+QEnMgd9PbJ++6S2ptYHd2IJOkr
L/5WFWBxrytFh47ky151Mx2S0zQECFlJfRVAhdwCCSU4w9Xbadj7oMEsgf8hQVXF
5HxJx0OqywfTIrtfJZehCNDyKtVcOSpDpO2c8roe4omO30nYdj5QwiQvGaC1MaNB
NWxxa2OPRVNRs5MnTCKIctQXQqZ0m7losa9ZtVvU4iZ+AdvaoO5Mwnw/0q/Vw86j
9V2YczT3wV1bxaDztcWR9dXQ/2ZQhgcOeITsNOFmKjZexeA/2geJWJED1RbsiYwB
VBe8fE5VcJWiBKv4PJGdww5ULO2kvppZ4c1cCbM+kKBJHCAxMcxRf65RdS0mCO0q
7Yp8TsUAq52EMHogYHn2R7dD1xl1rl5SQsIbYw9tuTT+sRBurg8jmicCMSS6s1ov
s2UEsN39VITDAt/wKLq7WbKsMecEMp7ru/ma6O2+SK8HMxGmtUzdm/Iy8dDCbwqe
lftJe/gBuR4MUda7BQIMzO8CVEZW2DS+bDpcbcLXOJEEH+3gqn41TvLKUjBPwLsy
UIgtZWn8rHAYJ2BlQPYSRysUwQ4AZxF/Rl/eATZF2fqDgNOddwhon1Q9S4Eh5gFy
GjkvFnqWTNyRK+zrd6S4YboHXA+I/lcpK7FIfZ2SRjfu++zjqHYA9fztjdmY9D3H
QSZIl1hg9/HD7HJJJntZFr8aZdt06IIGtYor/R/1u4EzLOXcbfxteWWd1xbG9tHS
24kJvw96IhAnQM6RPk0xf965cG7eB6KW6gizbaXfdsHPQvlPyeYjANbAK5Vb42jo
cFESKdwYhqdYW0Bht6L16950MA7Zem0PttO9bVutJo3kWKccXpC0WmaRbA7ZXbZi
X6kvnyLgHyKnKXe6KVQ2Uvl5K0XBXp0fIhedpTfoydiB+5BvTCrNwAwQxFIh/Fcv
o3ABJkyxE6Crf6MCKWlDTQoufndBjXzoJgcc7Ezfw2PiGLd2eMrXRCQXZ1VpWMGw
OYToDTVj+MoXgohEKEDXaRvn1hGrLg7axNk4OAs5MW3zfEyQ8xv69PwYMxuef8js
n/xfzNdFdJ2iCqBtIRlVolpXTdOl3b36vs4M44xu0GlGxEdh5LysfWhhaMgWoUAn
tjPy7xB6Ohe3OuXgESgHIcST/i3CPDFsV6xRIX/bJeIHZYdjkx5mVqVRfV6xePXq
n3CzigkWPBO78oTfmbTA05bvoVi41Rec3U8SN1OI+J1WDyWB3Kg96zb8PPEE2LvF
1XNszMnaZ4QHuLGh31b4yJqOb+ErJJgEKV6UCNmGzI/2xEAOxRO1B5UBf3KezyCX
QjzhdetqJW2eNNb6wTpSE3P/v8I4IEdhtOsdtkt/6BQ3a8q0ClM1qUfgt300PRIS
tbMYpOxezNpsd/LMSUhm5iJwv3RtsMcdh5P925YMq5DS84CT8nX6wQP3SIr441m+
2dLqcRabpZCgAN2PGfjwww0Xbhlvjt/U3x5uLI/J4kHxh0CoW+D114241wlWiMUP
mu2nrgKekG1LQzazraeBe1tgFWn7alfdj8/rblonQXwwSylJ5U0K/n+LOa8EfpLv
aodcO2RuIL/wu6d/ytXI9nuxsFv1OM+HTkpjJkXR81L/Pp8TyFmtkp4TAtV7mSKT
d7us4BYjymbPmBfqPDcYb75nuRqzK0QmJxjo2C/PKFHnkplZunt/geJUCYLbbSq0
T8FafdjVxDVLorFySfAODceYsk1Sjn9V9m2EENfnv5eppjcEV1hDZ/frDcyjk//o
RYlbylWHk/kS670N55CKAxWhZmiZGSsdSXBpWYMutJiQZP47ivNC7PtLZbvCPM6H
e/8c0Qy6TSMp/rROrz9BC87FQW60vvknjJHcC1IlSS30YOuyGiEDor3675S6nWKi
g+GKU3RaHrY4S7egOmSR/gPPNjmlUDIFkniZCQ8Wesc9zkQjPkrvmpbX+wphwyHK
QY2eOEixGdewW71cghVoxQbq6QuhnXq+/InUX6LlGoR2q39jKPajFQgRuWQz02BH
Z7LJzqDZfKkSOKzZAUpZ1oGxqcQgIxx+b+UlzlBCUKta6f5LyWBeEhI2UQ1EAcw5
5BDAUKpvEG2ktXC7Y/hEijbBXKr7vNtSsgwPJ+ziTC4l5GjRRWnDq6GpJqHy9dyG
Zqwu48Yp+89l9wuEMwx6OHhWCVDZdCPV5t2WgBzwt8sR435OHKdBZ8lRnkwC6zZR
fdwR7QeYB9qPin3Lz8KnmbxGlfp4l+4E+9JPy3dOAN23cT165gsNCKolaTetKQ+X
DZzcHuhFbkxlMf6eoSh+iwXKVBW2NCD4pO/qqTN2CPbceLKoB2QYEsuswME6/9Q+
xGWbSwGIFYOXPqQADdff6nd7dffuyynUc9q2pvhByVylEiGzrpwzsoandPclYu+/
6O4Mot0ela8kCBvVJfiUcU7MAr70CjmX3CW9WsckJnzLddo/sRfUu3LuD/y5JpS0
ZIrzfQgkHHh+/Bbm49ceyjLbsrA2d0fiFXUvlYugjI3QDKdtSdJEmUo34HhwZqri
1tAiBenRNpWuP4t4e1bXm0fshzFcdPR7V2Jc8cQ1XUGIpmqnmKzBa6ON5o75v68/
xIAAk0sEHRyEjwrUktdNKmgCstbs/T/worFDxsQvU1OqaQN0dV4+WTDx0Hk1/foP
bdv85u9ylc6BhOSePSbU9LdImkESrFC4eVqVNk4OxhkMe4ZGBmeN1bC4K5iC2EQB
OAzRbhJmXg204u4oms5/IdMbsWxUXOG33VdiWw2zyUAyRMC1iMSpDPtTTi+ypOfj
YJIhHDBEffRvhBkjK05sOmRGhkuBDvRRVAiFQ4OF3PGnqSLvofbJV3SHcqyhnDrM
bjMieijB6e47v0MdO6iiEguf/NwSTNuqT9buvJJd4J/twcMrTZfydq8oroygtOj3
Z4xyMpLzmfCljyOvFeEJY52S7BfGhufDVwVNJBZ2WNplPxKRd3YVw19/JZ7/3Npl
Iqf49/S24u8J4sfscTOEZdg2/13bs5+RLd1NpAPv34XipFA30r2XUOSVdxuL8CxL
hWg9qY4DDpB4nMc+6ZuiCQ08g5kR62nK5QBJHK9tJE/jHSTf0sBo/LTbWc73uGfU
lOabrmbnWG88bUMl9fwKJ2DgBU0LoH8oEsuSZ8572QIcrjTAxTyVr1hvbuGxCca6
E9aOqM8Y4PMk+PNggOzD0gj9FWvSLmii6zgOQf+Y+tsz5LEvVNJSO4MfiQbPs+hB
brKjQNnwt48MTN/cUeWk1zpiXrUXgrnTvbB8jqXM7CmetttoAKqYi75EVr/ai9Uq
Jtl/xm0STQp62FHkhrHAokW6M+9HbVhBC4BIeZ266AWMGWyyllvD0468pb05ZDcV
SPRRSieoBVOzcZDOWznHKxuiygVdVN7helXnLiduKzHOumySgrFFTQuwIx/ac7Hm
iuoSiQevdRgfExcsW66uVGkM8ycc1eeZjnZnScwM65YCmaOoM36szbYM7MNgkAyU
Hhvk2ghW7LoSZA4XUOYxSw+Mdc0c73zkVhwSohTUkGA+L/qXsr9vohrSZPV1Vsma
hZg9SquiFf1XK7xWGAz8+j8XZZve9Jgw50BE0M242d5KPVfhblPMhTWV3s/qkYBJ
BXWi2xn8zaNaZKuUFQrGm1C5fY7RddMOpMHHUwwfx6E+twlRuD1ebpsSYxQ1oY5a
emQ8FsxE6eR33/HK9gAt87/NwJfiFHqyzOz98v9ceScAV1cpX8wzNGvFE4Q+tKGM
6GAUylrmakGMyHO2QlJEfRhJfv6Po4Ef3YGRbHKe8lorxQvIvT3Ls+17U02Ai06X
F2KsuDvxPPrfMp7309oxGvejTWryhyUph1SKVd1xk8/HSdDeXQdq6LbJwNPacZ9l
PdyuqaATCfrna9yh+7P6QACFu9ZZaUNY4w0UU2/LAeKYV7hzhkIi8qrNR+fsu9Db
rTNBtqsDBSAznTU45iFKEYeCpq/5ntsOjyZcwp4Xbbk4ISQkFcYms/K+TK1oIq4K
EZ/3KgPsA3ouaZ2gE7y1a0L4/3NqQazUqibTDmzIjobhMO6pVWlK7wS3rINysBOB
rDVKoTEwT7uy9x/oEljcS3KGlU5MTeU907gxiKxRNl4/iBUTT/dLsWAd0fKzn+2w
yAzxADcPI29yVDsz/zBiu9WBHbSfh+QQwWRKvao86SesqSclms5DdcgJVAZagGgl
5cZc2Rj/vvAGnEk1Ct0yNv+0UfZXU4H5ncR+UL/ZCX30m453JwgkyBelvfjNZL3M
EzOdtTBmtDzmaC8cRK02y1aMQcloC4m1yUuq4mX5SAAJCkY3ekHqtJiFUD2zqmYY
U3scRqmyg1EKahhWD+bxTrG8eH7XmThmQV6DZfe8AAX8/T/LKGMthS3/ERCm2Tu6
dj9jdn28pqqYhD0sGDh2F4xJDPkV0r/BCYCb65QbOsRRZ3wQ0DEIN8U229BBawR3
XS27XZj0GZNsK8xlA5pMoqfDJ8pC3cLXhAUodA5d4N9bGPMYbTXr1iCouK6nJOya
TIJONPAlUSnorN3+EfrGYRzjsT7T8TgCRTCiAnPbOlQ0wrra5o9p9H45zh0ANpQ6
fO4f0s2ljE72ctOsa2BBthy8x7A8jbOgbtfNABSwCB47psTgVb2dYn6H34w789sT
4ck7vsU7+tnZZ3B7IdP2/eiwUq8mdzwZcXCMnpmLIFSOmN/WWcRRyocOm6eDByRm
SCwAaM4biBoVS2voNLNH6AjDlA3jcVxV0hiToHPQP8p5pw1CsiA1JcLDh9mtA7cn
dsUxsTHgcKYNhPnqsqEr8PjFmozy8ksieqeFjiBOTOC8Vxf3KTji6xELvpD7T3js
liSQkCVT2gYGj/sOuVBhQkcVhAzutHtirN2rRN+d2g+I1pZCo/7l/IyX2goKIf1T
9vcLFTq6maHkzut5EZDPDTKlx5eGT+k92MtjIujGwWJd7EIct5FFF03W8OKOdlsR
5QrprgvbZm4BAsukPAqoKr3xuYnltdQPlANarXIzUyIjVlfaY3PNHewaU18EwrUO
ETZmCaxBeZxRy6BCNMWeAfKsTr6cJem0BfdDaAzVK+zO2H6rN5sbcbXBbN2zZ40R
EO9qVcIUYjtG8GZAOJ7BOB6vgwiF77GQSa2uNYHjDpVIU0slDOSWrNSPWuD29EnY
XdjqMoXBnLYgpd/mQB0COOPZimn2vvfNgwTmgecxiFp7xjamMvUPGwY7Exi59J1h
cY4lLcBJpysbR2eKJfBFk/k4ojWT3ooCn4fT7iQCtPOSLqe98iWpJNzinPZ9Gnxq
dumTxKU/9QJdj4O/kyeyEAwnMeVIQrMdUV0kxzUvb0SN2t0f338wJIbBfke/s2kE
99gTWNI51QAifBzPEOxEx9BWrZbO5JF6jBkMjWDA285mN+otniIiYMTbYOseYqxn
+UA8mRDwony9URc51/E1iNxuFj0OemyvlPRKIVu4zVKhxUvs62fq4sqC+CPbViuy
7jinB2/cEk7wV3RKK+4oKFMxruwfkXCX2r22Dy12FcMbFUCGPj6L/IKlUIsVIJeo
MIk7y9gHgE9TxNg9cr6P/PESs94VcwrPaGBEK6iK7SoGkeRC5dqi3zvt9fls4xVK
ItOLwXVMAZBKEjyoZhexJvNBVaCv7QR3oxjUfy6WUPaIHCLQw+tAQ3V6bcUNWBC9
+Eptoo86mG3M3KiVpQRqp22zW8QApLEPZaF/wbAOTUSKw7sIXbZef6Y8k5SL9PQe
9n6wpIa2buxeP78BXA5AocHvoPWrGI9hgVa+9rHuNhdwOVDr2n0k9N++SVhDjiy8
bjnRtikX0Sn8OP6RGrtGrJCb5H3J5/9FTerCHUkwpRpKuqwCWInambMuxqs0/+ob
2z0SksQI4XOcea6hS5ZAFEn3QQ7unLoMKire4DNgwJQsrh5uMjDvYuor4TlhXjj1
AhkGvStS/w4Ynzc2YvmkE+rWnu8RGqbJliyQfqb6aOoicAw4fl66J4hGbvLYLLci
F105jdmq8gAtXKYW5uSWr5Wl73c581ZpbxC78gCuBtMVxLhxajzrO9Uc6WMWlaq+
HVAFs5k3yeZ9jxKf6o618/yia3Tz+8o78T5EFuOtGvkn6Gslv+5oCNbjEvgF33/6
qL4+P+uc6jSbVmC2jCHSmtYGhQkGLlka7dstjvrmJ0SggZE9BRfMyz9AgZj40gQi
Zsfrf71LqCI7q/FLPypDTD5qYuGvwhreQs0+9GpGA29mOMmJGfcaa9QPMFkQ/hXj
IAiAFBtr1OrAPCtCa4CNpa6xkQAQBYEQ9rSA16iI372snTxI1KIKYfVZ073abUFY
PruV4sLBMT6HCbr8J0CoBY67FR3IYxZDrdrlluS9SR8s6Zvh9Q6Z+g7S+vVvKexh
G+4QEdAVRMknE2D05/iRluXVZdhH2KPsXaFvHMnBzTp1KYJQOYju9TouZZYXHu8p
LDqjxe6wfjPJ7zbxGUCsxCEAwJS7YZt66/zDQr3DvCWS/t93O/6Xgu9JhoJK/g2y
0h200OCcLlsjpHHg5ktEE3i81b2AKoXcT6zYCVA2R9ggIJ5S/rhiwqBTKx60Qfbj
bp8Qafg2sfHraQ7+EkSUs5t75PIhAA09GYWvq/byKiUkiHS3j2tkSIAca4dDlg5U
C1TiCgqCpsWn5kWU2LSiucn0/oYuLuqyy37HG1bLYxE8y7kRuPct9qkEv3I4X7jz
BqPQvfoRr76XalRfzfR840RCQGNWc4Kh8YXGRhqJJjRPD0764ijvYHVFZ/kzPogT
C5dV4T98yD59XOIemFGkvRU14jWSliLJNzCUg5jXHE0oOTuQ0Vakuf4JE4uir3Xn
8ws7kI3dzQ2VYsgAdmCRDApU3r87DhIWKpfrrr10EipQOHDveMWpn8VnQPMZ482c
n37oXX77w+yibQb9ERH8jNu7Xk7o7xrIuQu3StFmuwPuLm+x6pWjQKUibjG895Fy
YG6sdNL3KCcyO2Jtw7NN0fbeuZH+mSKXI7udZ/TkCCmr7fpGh56O7EX7dz+Xu2jI
9xFKO590hcdFD2xYl0ODsyJCy//ZrweZQ1EUP9YyqsjC7q0rOO2VKZv/y6/4mx0/
9l+I+fQIyvPG1GBFDcE+UBDnv7roMiLpwWsUOkI+/Pl5guj/V73YjjkNpYUcdS90
lj1q96TyZzC7Tuh3/T4pI4z9e/wzltKoel42tGEDjHik3gYMtOPciA6piF/MTu9Y
h/iTXERRNL8eClXTSWCVpP4Kd9zaDoniJgIo9SynL3PVhYVzLQtUykuIEZTja/oi
e0yJTvGEsyVRPopyTvdcmLcC8Z+f1FFdhNdLiIpSyAZBPFsuif+QdBQHmFu3oxR2
k+SibupwxvU+TAHq4dGI2b8u5Eu5ar31FJUNhrlZ4poUXwzebMg4d6gEdnq9kGTE
8/c0hMzt6Ab03KEhEBzz6UKYuvr0PsE/obndxafci+hTd2+fdivbIBw3XYZ5oeiC
DULktPBKDqXF0Fydr6UqEolARS9hCC3aPc3u9qEdywCbNL9ufr293SoQXSb0ngoQ
Ng5sLasrLCHrdIG2In7CvPvU/tr85Fy4vXd3wMZheg1KhuFG35fWbOd0cxgZkAkC
39CodE0Q+6+9/PVV3xgLy93guB4oMqKLzLiPKUKgkUQ/HjAIChIafccgYZykFpWZ
q7Sp0NQ4dUs+m/AqX/Sth7G+CJRzXEGuDxM2MevDxkyeuRXTD9iHUZ4PvvsnonZf
T/P1w1qNj+e1qByImXr46LH0+IOjA5OOdoxawMyw2XsBVsBiuQqOeRcGJZBKvB0a
8ABNwgLn83p8gF4v6WF24kEs/p5fHvS5IVzdQZN7ipt6exYYg03U9dQVTbKxEcFS
yvCCQGS8arp+L851TZHBbsWho+DxfVu2TSY+zr69QNvSiOuOOKomMB1giGBM4X/l
MgM7HRksbS3qS89RUOxF8qFckxGeBw5HX+e+U0kKIOna55kzYJ/5CtRs7/Xguw2i
CSYXfE2CFe77wtWasMI1VnZEo4P9cNVVJXG8Mg4RoRKGXONbr4TB+/gd3z1HOv4E
9ztbl18GGoE56l5pxyOchYPEzslL6SKdOyw7/8VIF8YLhgEGd0LiT8GF8+4YeUj7
RZ6zT9Q7KOHb3vj1M0DcF2ZxdSTAU7mQwsFqDMvWnff/DP69tM9doDuUM2eod+Ya
76CVyt3xhoeTr839JjAu+YrDistGWZtO1i2GxqCzcaxjNRFTDMwcLHgguc3GeOZq
7Q2Qr1um9ugZtiVAKHnhxSUTuNWdAu/PKb55i6K4JsxpXeCc0wsHhYZyI8Imvt7Z
XAPNoD9Y12svA1+vwYRaXqYO5bfB952/gOWjeWa0kute2yfaL2j7EWxUP9W3wEJ3
PDfZO1p/tNtxcWc/56BvkP2kdfaFOumESuSOBfpdip6sZpl6gkyo02KfjY/lRhSh
Wif27AZfFJ6deNoASIMeYPmPb8SNMPT+vC4etpplaUnYcizfe/30KrOV726QlwJG
1EZqraAAKrPcndwdgZrn8z97UMn1iQr867puWeS7Cufx73FqnNctlWGAdjAyXaBE
+naCKcCMeAnj8i1PyG2PrSxuUyfvPbNgKtxduRSPVw3z+DowYQqMctCXLxd46s3i
EPab+zN3PgaDF80vnLQqmqZ/MqdNROp6I7tf6C51EtoC+SHm1GkBWXOxf7zK9l80
Sa8d//ASPGGbnU+W9ZJ2jngdTWCejVxVAafPHKHto8SV4BBdYplpfw7SwM3iR/du
MS4fWfi5x6TvmVKxk0HwFeEzKdj8zUX8FGLsGGZyD90HYgBmOzYyguHfZoxTTnRY
MSzNg2vfjEL7ZJLtu8HwMAqdh06FKZJbWso+soiGqeKUQ4/LhhYwA++XoGNSHjmy
3KXFtuhDEidj4s+qdkqL0xnYi3QvbacAT+aCkEvi+4cI4E1/ABJqHpR7aZ7o+yWR
YiLE5tgF/KJbGgbA/bIG8kOh6+r/aZ8/BecsUgC6d8fiHSN9JM0eB31R5DE5dgwn
ELJ1jDnwyh6UIfb7x9jqvdcCG/vky1e7sDZrC9kHRTg8fg/G5SmDeKa0BaMXDmys
PcgLW21rbNaQEC9btJwU87QlT4whaO7rsIvTf/59L9QtYGl81zps0NKTuO1nEqeO
36fmtfjJP7W3yaBtokyWDyvvEwC122eGO+p4s2EwFgc9MIey4eOBJmescaOqj+T2
5rjnnGb2f53Jj4P5lERoHdHet8tezcUI340xnjSBLoPEchQNz9ud+t1ZgJRsggOr
42IV1QX+BzKarfaCXpsg8rKvJH/T8Cat3VUcFml1Cfk+eM+wNFcWnM00hxSNaVES
aWewb8IT3z69c+YRwYnzERk4VOGNRQdF6iILp/bTk8UoWIAUfcIyaxw3Ast4Mx51
HmyXwlVaghzD626eJVC/d/AMJ8IJEua51gNJDLnHCU1DLuWAGJurPqwD7rD9JuW1
tNND7AfYLyob+ODC+bI+eN9AfPkv1ajZruttj+K0KX7HzTspI04hEJ07OZDplsR9
IZzWD1YJMdwNprnDnskVYFpAawJifgJ0gE/rU1/lkqdyzLxWFjEQXG6wZyFdnN7U
SF7jXE6oFjGT6kVK5Ss6PfCg6wiYAR29622pPY4PoiRBl8d7aLmXmKMdiOMqzXhB
WrunVAtgRjDyZLZE8o1w1tCU5u2DSDsMvAodOyU6uBzdkSL/hSI3feeSijIx7+ow
MaWx2bwOueQImKXCQ7dZgfG4HSwcRzAx+JKM1wkQUD46wUiAAVuA/ptzemMWFCfb
/nMVSc3xB69LzcH5ZGoUrutcVwsumNZltE11mjvP8JfcZoDyUmNKPNbh6JETWVpJ
ORjRz0f/b7JscIjyjpmI4TJzDKKDaIe94eqbM/XAbP2KAY1z5IKy6uFGLUIu0n3/
J8g5GHoei78IHWhZtTmCdrcxvpPdK6WDtokDncf+lWDsOAD4EUzu266StCWXeYBf
tdKDPxtKrPTcVxbVUrMp6kZnSRtdPV8mXsa9KtyBTQsSny3IiysgtNgCOT3WaTel
RWHZtSrAQ7Mg34/7JlJwnk+lvm4PcKBmlayH6fcCga9hGgBI75yDnGbG9mZ6u2oW
EbLFr1YTswZiDlxzKuDOa3O2ytUT+f0Sk/o7Qi43a6ovaWTKUBegU6u7tGVUZIBf
1QGtavemQNqQ6e3BBryE7rSKJtnK5RKcgx9Em4tBvYhoBkdYUjZdglX87pAIFPV/
ujfxbBbk4PC1LWrxqE9IzjcM7MND6Sln/nBjV0oOXjhnor7ufnPRVpqopjUKR43i
XDW982uOvySRa/HjWtlzrWiCJqTUlqtzR08tMi5kEJ2yfWZXMcB8rpIGNUgCHnrF
uQaUxpPCqM6u7njyKkwqXIhN4A+Rrw36/wwRyNWgz5Y7YhViEJA7SceDnLuX6+Yh
IN5iO+ylWpwtxR6rGmjNxODykt5b2wxIbr2UlLmhh/hY6zrlbDI1Mg0njKNmODhf
kYPfp48Rkr3V5nLKFjCjXcg7KMvPULAThwHBPbHCQyeQ9nCl8cT2yuKcRgmOSm07
/KEubaUrBZ0s71lkgQsI/UOaWt7qY+kemEQ/0hysNoPUMQ9iUHodUNqbBnculIZe
Zmvph0Q72u8xYMsEWD4JA0Vq4EbXQjhzWRcvda+uWfl9SoKgWjvTx1T1fZTj1YA7
5Wyf0cxqRqLvaKQLCMuz720BAYyTdDKmLZoFtpaP+RWf9ZmOPP+92//n7MHvkLLY
N0mCKk2jo1U8uztNbGgsyiIam3qywkGiEzS89ho0TMLpTrl5SnubZ+RQEqMaYEiM
coWTp7n1Wx9tw+ylNfYGUeaiscrVB2ooIMn4Bnu1sTWPzVPxs/Fh8Cp4JEPZBwlW
n5adOoIetDWy3gM6GjzsFi8k1tx76vBPzuUkOF2/XTS9Pem1W8gvYIuhqVMcPIK8
/IAVBg/snUrWY8Zrk9hbR+faYSpd6YvetCQIVsEQIP502zB/8eK0w8BslJUFYVRJ
UMsvHvZI2BMvEEXClGR49JfHH44rpAaphPzy1h+VINV6qCVAdumjvtGY52ywU3Be
pfODtidJ5Ro4lR+37ejpeSaPt3xFimK/oyA83sSEjGk1xUzLhRvSy67+AbgqHMUU
+8U/RCchuhWVSIvhOZQmzYYXaP5SOCUYL7Agvs83EAprHOBsBfFGn8QJN3KY2pfm
qyr9pbskd0JYrTiskKQ6z/wXr/TsAvZm5vNz083f1zFH6Rp84glfDXLumX7vW4VQ
Dz27V0smB+zu1lYrTWQe5SrsgcCGKF02ZbP/tIbGdsaqUsGQjill18TA3lvjnyJX
TCBHwND8pfVyvO0SKUuoIy5QWGoNDTqSHsvYnLqOX1athKYMqHUjbqpDGFnrVD+u
AXoaG+MhOaKSAsOEt2bTekF3DCURhGR9Cgym6xb0WjuYfGBOZCDAJ6+dERQloMQx
OZVomqD5EiXa9XCIAU6zgmPLfjjWM0YevaAg8ZJ0yUgHlrvB/thXV2QHrHz8XMkD
cKPj7CmENPLU4ateIvkFpjedCm+JmTmPUmMeKh/gtH7/sbyOp00bep5ZQJxaGMd5
JmmAjkJ1xeTO/FUB8HlCLOxeXLHtTfWKgiryYf6zWLLDlbXtO91aPdcPNDp3PVQ4
7gPEAo8IxvwMxxHxfaZtWKCYVQCykoRRsXw+1S05DGRzVh4wLs29Oy5cshB3Rfop
6ZqR+m3ckBKa0QO29YJ3GyLgSBswmqvdieUnf2Mr3zSuYiBmHTNOSFWwiRQIRznG
3FsPYnNsGkSdijNGLwbty5e3i3eYNzTUF6Z6IZ1HuAujtgBex6FexaahoACHmfiq
9grkZwdM/nXO1Q4gjXduP76dyoPQp/4GP4TR+orjCQpd0cEA+1DlVOmTl33o5Izb
t+VDnUqQdltpgK1v42zdjmX6YEOOfP4rkjyEN4MoA93+MdpLF56UspC4zyvxUnrK
BuCXeQNXpYtpd1alQSaPGNsgLJ9dgbnUuEjFg3wjFH5/LV6mSPjMj+uiT81qe+TJ
sChU6KzsHmpndIXIp0aImXkN4aLf3iMzwgxBCInov2IkpKBkn7LltMIPBgTALeM5
o9sATo335b60lkFWrZwsLyECa+sdb0JW+7UUUK73DViKVnAWeU8s98EVcupVm9mp
ZR1Jityg1i0XHe4uosDZhb8BMueGI0Cv76vq8c1uvBxYG8YRF9eubaSk6gl+hQ+B
YukbVYLRnn+F5UYMkmqRQ5n1TNU+/cpAW/I80jqW8H+M415Ks1aJEcCea5NgbACv
nFX09qNC6uowQw9UmVtS0wrhBXE0qo9/J4C6ZDrFg8kjrHzgXPkdSi7RPn7c5HAn
TqC+n6b0AXuVUKaXy61z3lbnbiv/zXIoghQazfoY+ZTcDKkDCdrikej0Pdi8qm0p
u8IOkDtNrIZH21lfsAxkdEHygb7QJuG5aA3k0HVWK6yISESQJNvIHG5ygx+HMbt6
zKZWX6r4SUEOj2lMOTB6xlDsTTgM+MtmAjrZUBVv1IebBDCZ9hWV/lHYbai8kzDB
CdyXgzUkzcJUokYOAcX1VuvbQntPTd7PasCh59iSgoZPq1e4eRM+54g14THb2fKM
Vesx0VhShFyuy92TSLTjzaLlZs9RqPN4eRpt7FTBiQzOGngmco+fc5T+GXZqsL9l
M/jqaA6kQnTGRg8iUyrePtMLxY907p9ccW7tT5iRwu5UZnAQE+K7XnUazlknvuhB
pTx/K2SHUk46zitk4Wzw6CnqmKnd/MIwsGl4mbEwchcSNraC4XZqgpYu3f04FZKl
cGmEnwjKTb2YoneXSPXcyKd5M6bU1ii3zTi97+eHrRXS2LYso6qga5nOa0pO/P5T
GS/qtJJ3JiD67oR7kehstoJZpyUf2DP6WLnY8d6L/R7/V6i7cmMHjlw5jcF4k2gX
CSj02TaKfovQcxORFYsAnNefM+tTipUi67RQztRxY9AQ/4HjJKSIgQaHaZ6gOume
7ebEwt+dpaO0t3xuHvoIuCnNekCNeDZ4gI6P7AZdxbpg8FZavNIEWEFDRAF6Ufwe
lJDaX5d9/ybL4xqm/FlBjozDT3gwFZOWWRUFWLEOTT7E7ocKhYbeimiVh+nItJ6M
v60r21JmwD6cZr1S3g4i/wjV9A7bdUdpMEfk4DtrP2FneVhCjnv8zGmWsA4dL116
/7Ir6NHzH+44ku41y8dk/0ekE+AsKMjshs6aLpbUUQIXh0AJ276T4MeHxfgfkSzs
AYBzNUZUWGeFevouqcktvrXrysKxITOcDACwvtTdDuDvYHYGQ8bv61HHD5jLVqlk
Npjs0c9ekg7yYPvZ1UoxidGpBmPF3TLGvSjLDg/Q/bYNo3kjstRfnTrcD3DvvUoh
4n4KynEqlS+L82T6CZ0IJuymAP+QNcufrQGlaUuB4Oxc2Qg0B2LJPbk9EtqLfAey
mltflNk/ikplxHk3rMe/6zcH7zb8Io0bfgkjPBMIOvgHeBFiCOiQTFhSd6dAnyUO
BvoJ+20+Pr/LQKuolsYIOeVPOluuVL9YKnEXfNUuB8wkaGA+c3fCDNWLhS5CqDp/
xGAlAnQV+UT/eb71grye/ptq/R3MLKZ9uL+KrE3rzkAfPYRiXXUwCGHwOl8Zn3Es
nuByN0+L/+r5gmkOp8nMXQUex5GjaxekwHXIXBCvahVjYdyVIenK25WgFUqVvAaE
NBTwD9vh2BdIl/VAB7JndnUE6Q9NliazGO01LZYJAwPgQSFaTLnzuSCwKXZFT8e5
PgKjGY5xhGODHr7ahelMaLfYThqMCHHFQaSiTv5ZzafFKURWCmDU3okMkZqfO//Q
coIRDUpl7skUuYjKhxhRhdXbf4xHUktcAQ3VOr0iDNCxAv4MS/GHloaw91Ia+qCQ
V/ZLqvZSG8GQvUxUEHVqGp9JcgHqtoyCMoWK3jhP5KtH4rn3gIhgmMPBiwV4nvNO
WKy9kCmIzoRotb+blR4rbhygjkc6DiWbrY5uIVRQHrgOgxKAhlc6gmL9lN02OfEB
yMddhTTUgX1GYDNdVSsxctnao0xkdN/kyI1BMINQbUH6F41MTLK8APq2yXk1Cb9B
k78w6EZb065AqLDdeNodLhM52294w4r7NyOAHFMIwmI1e+GU6QjqRuxRscccWOg5
pe6L8snmEZbfj0KN3qllUxch8mbEMOrwuBLmENOGoItPsgRUtzXVQXTEvDI/LXtC
LDqZn7ZjqD6xEaKREkGFcRH7XE7FB2j2/4JdnUbgmzUq8yXWmitYRv2lg+KHkYEW
aUsUJaUwwQFzKKUY3Ww5eFBLCWpGFRQfYv9+MaCDChN87IUBYrL8HzsRO28pe9HY
VY4eAH6JhdWrGIDbN+3XRUkyNK6IQbJGpBpM9VlcrrAaF9abnCTcFW/9rei2zfay
7okU50a8JJ+2JcQI31SinROxek3Piu3o657opIr4rdIN9PYiC28mzywB1UWzasFV
0cKMQt//c4EIWoDgLHVsyxmTFNBzPAly9QGNp+dr5dPmMD4D1j/8rXO3GTCw2Udz
ZlxjGENOdqN/M5fWiEtx9Oa+A9tqaQAP9Afx+8/+rcYabwZvxLN9hUm1PTj/vQod
TB4IVJhd8lVPOnEXRjF0+xh6eFj0/a+XQW/IM/zk4Y8+f3PX48rqVmb7kwt+UIyv
nI6RRiNtQN+Rq5cutwLd2bTUAoYfnjB60MlnDJW9mHtiX417ertjvCWuKPnTpTrN
P3A0z50ieaOPYfunuqIVRoCl8F1NkwVusVsZ1dfyyl3zjHP/AA04pYQAQqcUseVY
54RORLBNMHKJT+uCSOIfNTXzShlx2NIymdGiF6oXsqVOHByF3Z6yoLStf55CbNj4
GJ7lzO1mgxKRg3rqTueXGwyYoBZSHdqL4L9ONvhS/NYyRIR2FHLrYE24BcRdKonU
eVFP3TGyvg/1groIn6wD0E09vpr3+cEki3dHsIAinyyu9UtgVWXIdWtJDtcX0B/E
RjJVO5p1qxBo0Uav3cHfN7RJmx9bjhoqoKAd5R+5a5XIedB8hDQ7wrOlBEXrYq1a
i+kpNwYJSHqDhVLnU0u8UHoeK2QM1urVRkt7s8FrF2dJUtt0aV8Nrlf7wzXlrQre
2VuqnFnME4++UJ8RkZaZdKRdARcZ93lSUNXb3wC0HRuypqyMpKUPo2Q3zTDahqqm
r3Nyo9Skt94rpdSl8G/+yBbRiYQC3FGbz4DBUXQR0UWMITYYVGG7IJukivnZ7os4
SqVKK7iYJzKCD2GET0wSjGDgk08GD1HZIsbgHAiTv65FJzlo3t7ZoxWKQJ6dpoDq
dsTrSglfpXrDm68fhmNbWHYrB5NIyamCpSM956HYGqadPzeEsAzn6M87JIRkSTP0
kNEln+XGH4hlKpTInD87Gs5S4WeXw28GX2a5cCHlTganSuIse1LqgNOc1+YWe7Hz
HDbcci+R04YCO8Lrpq+gYOudm76KT3tWVvQ3PALpmehTJdYRI+tv7zzy7n4Xv0Wh
Ea9l3aYnSlBKgz2bYqiMY8VpGh8xc+A4T0zD+EIIheweuM/+kYvT6U9lzDxW5i5G
Ucwokp9oZFciwUUfgLRH2DUfY/xoD1ISgSKxdmUW4us1SCuXpf+QDVH+w11cx2hF
odT3TxDHy5xlRJVXIzrUdI24WJqi5uPRlsuedaw7FMPAw62DSVkgpvpkLF3Et8ps
EsRW/j9bJw+WWpjw1hOLzAFZ2B8tTIl6U2Ze9ZHlsWOtA+ZreuPf+rSOkSrOm1G3
zFJTdoz/l83CUW5On2JD0AgfAqptVGmRfCJ16Bng2DuFY6j6B9JgnRTphkqfwQt/
vUYqWyoutYhKSSNe53KaX2euRzcz6YvEj4kP/pYrp4xQc13a+Im4ti3Z+Nxd2yBs
SAmS1j2K2Q6sfpPJ2XmSRpxpqd3iqQzV1KRfHBarA6iTX0ZttzD2EAlyrH+gRgGy
We0KWVS/codJRfUSNrAQvnEbr8QsYa8qeAc+3BZxmuTJG49TVDBllPzg1gfFpRGl
ivh4KNo/vs/7RN6lH6qS5wEvdrVEbCB1e6b7m+KsoaIl6g4yUucCLV5cYQRMti+P
1mtksmrPFNdTZAzorZcLMSV8AOScIDfTtNjI960qv/iKKyIEYduN58IS3PKG49Vh
shSL5hjwjeqzodclryFgMBTRGsHAvmp50ZcGrBt2zciVWdtzTnp6r2de/owKUSjt
xBkLakJLj5UUTJwALagFx+UEQhwsA0G98muCpNizm5avMdJmlzVNh3iLLzt9y35/
VSlaazflH5pVWJPqqBQ8leVgP9kKBCJ6QilC6VbyFmQ=
`protect END_PROTECTED
