`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wegshS6ibIMNo0rvvWPvJPFZb5WPcB7xlUvOTTdPuZmSm7eSuLAIshBhplb/K73s
XBKjB9CEoHypfrgiKQwsDFMGuGMlMbuHuUXDPASYBn+U2UT+OaA8a4USqGZcEbNv
SV+xSpDpcCHQONK0ZbxMZCvbTrVOBQugIXAkdxZcSNIugObYiorfFSXTj/47NFjp
0jRT2sBc66eVfOD+SFveXbpJK83HdRSc+fB5OASlcItUTA9f1nA4cdZlvT6FjE0b
UkCrXkGX9pm0Jr3sv0fRVIl2Z8c8OKNBN67GjSFa+gK6te1A8l33Z7Ad9c8rp4jK
W3pVep8tNunQKq/aQsGSnZzClm6eU80ff7FyJb3oc65KFMA0zrf/C0fweNQdEECf
/rsPiSVpzmvOUmGzLjU/bMxT5eQv/PvcO17hTdU8dh+jh3QBBNvwIyqp0dQd4ktJ
2nM43kWtriQPBQxiX5+xB3/OqTfeLvUq5u5UcnCdutl+U4EhIsdvz+ICRoThgetO
RskysTMs/vZJx2u+Xj5fWCipT32wqoTkg0qnpOPZRu0SXBvgnSZt4daCwqXjiiOl
SQaGFrO2aV639wB3sQp3420xVo3p8QxkBWiDd9FKt5zKesuzV0aEwneN6qBjH+g4
3rFwJZw0XxLAmcrY0oEy3pTBZFMw4OGA5ifI2b/UetFqMfcON0pXpvWlFSyf6WBb
YyvWJsTNzJ5sHtNfBrYrP8t7JADgcOJa4bhMgI6SPbKuv0IYGH6Thf/RcwaRBmCv
EKw30jGFEAyYIStc6+ZYYLwt1RZKhP99PnaTtjMWNfljCu0t1vBBwiQSnmkj+0If
eKqD7WnPLxNfoI+cPUG+jdaZ/a7oD/BgsdODsmJIBSOE8l2q8pMBF/VHtPJSl0ly
MVL4fCaXeHelEyaLgbRaMpqOCHt/Yyte+gF9Ni6cVLb3YfE2fgBqdomLiK7OBrO2
kRcoTAOQVdC2jkuavtz6EQXKRX6vN+ZPpx+EhIlEN9VwY4b8vlZS+qsPpWSeMiml
zfhxibuMfTI6y7CwbDoLQtAotNFZDGgb24aMf/XsKdcKOEqDSJWHodg6x/OGVfzg
QGXtUK2EzZCffJPkdMntJYDsA/KvzyTSUJinH3e7ghbfyCVzuRZf8FeQp6wV53lK
E2og800ejsMB9xjShxSXPATXXKXY1Q/o7LnxNAVQuNK2Jyv2Al+9AUDEoyyfTld4
ph43YjeM3jsPVCXUWk30BB4YaFCDMs4nSEKzJ1R3cQDxJ+O4puwMPpXrv1/jggxE
qWtRcZbBtepjkI8YchnrFxBqPcLDVn3H0JCwDnOVIDCtQKWr7b/muSfDdGY6QZq5
TTONzJsPSO92HBC99c7nLlUGL0BxHoRLdtaUBphbce+m/As9W815fp3ZOa8Z383P
SH4U78W1Zjqwheu8u7sCcVLWNM0IA9hwVXkTjjv2Rlr6Znnt+1DcHc9vQZmt1YYk
r3Iar3PXkYP68oatwJx4CpwT6tOtMRw70t2XcDULrWRkdu0n1gsJ5QMxyN1NxEkD
RTaYseA2OKoRSYS/OEE0DuLSircCSh5vdQirzshp9pR+Vv+3FBoYXpGHT77/zq4W
l0TasDRLtvbOVC6stcZWbinc3mcpLbuYMRlaJgczMzc6V0aduakAXkNr4JfKYsiV
bpYBiGPHmZDnt0CWmx/lHQaiyPov88wZ09MOcIZnbqkcfltrcjEqGYdmlfVC780B
QoTmVi7jlmHlWY+EmrH0EseQTk5MXSDDcCj/AfGdyilvUXizKcIq25eYJxWcoaD4
owDq3qDoQ4A3Ks9K6oEEL3me0BLVnKlfXsNVoNz4p3XfWmJui4TN0PKEpYJ5aEPT
/JLRgAsme/eN+DvcMCDj3E/BICuF8nVEUEwXbO5gS6cn3HO8HWjVIM6XKWjXerFv
iDcedmdsrh/ssVQUrbHwOwleaUaH7LGLhhHOLOtJtL1z1DpEzEUqZ+0YL4/gZaKk
o0/1PfHnmgMtbJlVHJllwOs6RMjfslnYfWsZmfv0m91FwOYlXpXTJpJckwzCv1Cb
ldTY7jo+RP/ZbOaeuKwe9j2orOKQgxEOfsLZ27uAqsCZWZ1BME8s4g+wPWHcJF88
gzqvTJP06kcNx0HlzoFRmMEV3qy+olGyjjFflJQdP7qklfhPuIy7Tnb56HJTHhOG
J4OeM63ytRRzH6E7yewASy8rO2OxGDSfUpAJTUFThNVGEAwE/qoUi8kavED7DdX1
UuMZY8di/uLxVIxwNVLecSHg7cWgWqYSiRhbcC2cKLYXSPJ3rI9lMZGfrHwDcSxi
OtkYfFu3udiD0TkL9CirIW6zhFr7R8yAkXOkPUyeRfRT/wbqWTXM40NQlBo8HxGx
SO9R4ok8v7x4mOuVcsTiuOQEVOsQUXGux73C2hQ4t6Vn1ieZDvjgIvRQhWVGOI6h
FceNy6fz7I9ytbHZN9PBO4USseGkMN+HF5k4zyGvrDKZ8zepNKCiiIej9sYWhVZr
LKl6PWU6sGwQGPQVwQ//4nlnyJAYq8Pjy3sZNXUGhifeOnP6P83Eis9fWl+njKRf
Ckx2807qzqP2jzD3j0QhSwZPldEB/MFxideOJtz/tAcK0SGsQXoMdmeS57Yw8dPt
iL5dx5fIvizeozTwLWeJOoxhT0KZo7QdyeBOaqElwZqTH909QjmQth39fngK71dd
NQQtBH9jyzuHFiZMo6OWD8ardnfg+DcUv9mFeQ4lbGwIGpJmc3UM2gahf6ywG/Ri
lSkf25bvtBikyQGqZqw4IQHZyxoa7Ua+H10L/haN8ivk654Bj6l2+BZewmWzT0Z5
6bp0WH5Co8gyuLHnmqeMUA6SLQkaRfxciodmw0Um9qVK6h2oSGpywKS5UE3HSU8c
2vmB2aA5mLAl8PSkrWWCKmDx1dl+KxQ0Pha22TbKKfvyJu3GI14dkGVcyCZzC34d
/Srg0tz8Z4Eoa/Jcot8638tCY0q7C5S/1DxnelH5CcDFoQREOaSGkfGygQjynNyy
PHj72JVW5DoHZ4m7qQB7bA7/H/Mpurcy2psRos7MBaM/iN61KBZJyfz1a03ZZZ2x
edIL8glgHbm4NHuH+k1qwNPPX/y41rkYv8wYpb31VMwjWaPFGdIcfIHK1qaZXtNO
y2/S3k3IRjKdUcZJLxMrZczhwEahGG7iqbzQCxFNVt2Zp6L+/M0YUlgaCqq46qcS
ZYkb7XthcRgCX4Ocr+mPGwxnmrhImvvT4Gh0HGq6OP6wpFuN1lAZGButi26xTtmD
6cw7VCCRB7fOqm7pBFwZHIzSNjQU7Oqjb0J65vZdx6Q0WKUZ/mAPR37to7Rh3MTQ
8ur07/3tmuX/HS54rSp/qPpJIGE55yFUu+QUGtNrHwowjMpWbs5vShOwCL6sSL1O
IgqyYAcq5Nd54AcGZeNhDInYlJHWVBIUQQ9KOVlvz+3CvvOh6Pj6/Iy9oeLjtz/O
pQkZfCk5H4uleCg4sgUl+ubpdqNEyuUSMq6QBk8NfEETHxhd/mxrHMR2q0LL5t05
m7pKrLyPZz/wVzmvlDbGSnOOn22Sw7xGHyTTCuu1yQjaZz9xEuqlF4qsMAu3/Epu
Tiz41VK03evJTN8A+rbmBR5qSZkzd25PSMnpfr1F8j4hxrG2LwQAsOz+8BIxzqXl
Eshi0NZNQg9wDzdlbIj27WRdu1Rf1DaLp6JOqE5OrL7DZRt2Scdo66nccftav4Lw
EI3ugqD9acdM/ncUVqGFbYB0u8H8jjLOIZHMjBjFArtNwqAFoxvRNB1pJXpSI9Zk
DLyFKFUy4ckK0l4LJQuuIFLfuUb3ya4NuzyrrVnN6TAeSxxGRLVo5wk7us7thWAx
RB1ZQCUXEqvuE2HiozYcE1HzXl11a3bJoQkZ1aXl7UfySKy44SsljDNrwH+eH+uq
2UKGYNnFGmJU+xPwkUCveYI/AXBxv1fsefHeSgcLcTPp7MjNFzK5v9ZEUD2BSte/
NQPGQgzF2H2PUC4tBuy1MXqbIs9wLU+Fk7qK26pc4kUu4JVz31W7Mwvr1zERWYXa
ftS/ZHccql6gQegCuXRMAcPR4RAkTzu3+YUQKM+FEkIZTrZzZK4E+LnT+QGzQ21L
+d/QhMl03xKlhaJ5Aj/3x1L8HRV64OGan/ucTF54kp9zem76flcuy75Av8MFer15
PJ+1XHHRH8M9nCqs+Hj7EwGU3owYTR6PZrrI+Jg4wQZPZZo1tjjvCWSebTvi2Ebq
GST9iZdbCwQUefkM2VnDTOhnuU79m17tQNderPCFyPtp7exoSEP9SoETv6UrjDJo
bKcAm54qiviHqbXoBr9DTHIsEwtAheXIBTStk3CjbB/2cf3nKAMmQu2dpokenC0B
4S3PbeQw0/R1thuzIy2c10gU7H8vAKNa9WjSL410Q+1E0Kzc1H2S6a7yzKU6ELkr
bJSymseNbYHGBPDAqNV1jcIEdRcGCzLJ8eCOdadwi9/Zb4xNtYCbTOX31Dcb5oiI
9VeCo6HQX7qe4josPRFHMAbD8b11v5D5d0GGujTr77rVH4YCVD/B0Je+NS3d45BG
XqjbzobzJ0W97KIjr1hJckAdTX3ipSF2PqVOAovSg8BH4z1r4HHbFzB6EJz1BQSK
ykKgtxMSwFuqWp5asBFLAZ4WIUUXGaWeEJ39zHu5QJGGQDDJW+Oac8703Uh3je9K
6PEcMFezhupXMJ3+wrcbVqKZZxpDW9pimz6rNGCp1MwG6SVNCl25dr1DyzxB+cFx
fME4oggflAsX1+XbXO16495Cm5JEWabCbB3rQtZZbOQOrVVTZ79KbCK9LeXNEwRe
pA3jZ5btzk9RtMEyRC0Wck9b7oI06a87D1zoJTE2GvcL5/KOiL03VyAfUh/mgbW7
fb0h7PwragZzI0qTeTruNG3grl2jOu3ayIlkknPBmkMjr2vv86nJFPtZwRMcGlNy
EZfCDAG27lozWV5vEEM5hGjZ2Qw0uueP38uXn3if//yls0a9sp0YqWbzvKOjI0iB
fWlTK40EgXu6M7E0rvIUCu+vslp1dNSXbT1bzZIaBKAHXPmn9+un5ApkFNOSXpx3
ePgGfi1MDmRHVox5cTZc93XOjKCD7Z5hcWOzITM9K4SQvAFLlwKfYW2j6cDbs2AP
czovOPd8RwOnMbaCMKD0Y65pvIda/6c6MggmYO71z3gZkoRvr1DBzzc9U1YMRBps
366De/bowTaXEN7t776pOAEMANKdsgZX31rx1SP2a3l/6BldqKtGE0T5RiXe1f6u
yJSnBsb1P/OIsoDWvcjcXjlgAsJKRfgw4mlyHhZpbv4WeLBZO0MMyhRZ2nu25DQC
aOvtR/ovIzRAbi5LRR1OlxqQRoFrlkexjC2kG0Ry01ET6lPgstPj4R2M+Mt1K92V
NrZsX3UKN+CY5GEsBbwHalRYu7BrhY52UoyFQorqXBc0JMJM4M/2wUIWXmodei/9
ym3kpWoEdgDShAeE9aTb8fZngeeuO+MaS0KhdWQ/GcsJoKFXkkDwSxOiLWvb9RHo
d8xCcWTp2eq/rvAyzJYFb6gVn/t7jHiHHKMXoP+mQd5TOAnWIrFlyKtUS0JVGcQl
7m4ajxK5HBqyPb147zPUkfbpnfeoCZ0wa1kODTP8Li6jptffmQB5fqYyui64r/Cy
XoTJN1r5pCbgSpMLiZEabSGfXbIDil9ZmLQVwAxqWyhmsaNCrXrXOJQZetHazgAJ
`protect END_PROTECTED
