`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tt1DsHVLDzZsKPI3cAayo5Dtzp2xolgopzwkyF4lVzmFOiiGdm8zsVLLyG2YuN5d
JBgH63gtApfHH9Q6V0O5tzlUYuU+dxVQCHfzvtymsoKtfV5MvfxyX0bG2/p7FXRC
eEJZobz+Sq+0V32yepBnIUPh3Rbta3UlF0RwMu8dYFLl+OJzEY+ZlC14p+6R3rDH
cz9LCKSjaOcAiJtA7qJyPhWq4ZNJWPGnvxAl/SkOvXhpyPXfvMRLlpRToHI1PCYv
6smZomoAso5Z6itpICWRonBnra31RMSEhvuh3B2uPIlwCvc6UbcpW4/NwublLqoF
XKdb6LKBKoSNX3AjhCAar2aEqjEe4vlHnlIdWs4aWdyt29uoOrYXUh1WgtC66qap
XCf3o3n7r2CmLo5zdzQmxIVSn7KkBZCBH+wA4Ade6AQ2d4AAnnjo7gC9RlCFm/pN
GXCooRbbsCoLmK6ftfKFp+AC9pBPYVG7sMaMmudaXKPBXLUoSdbenxdDkSgorAsL
oQJoIgKPI8/0nNjKE8wFASlfF4mSoDR0+bYQA6uTMU3rWUzmp1d8gSDemT77ixaw
9l9nSXwIvx6ZZj3zX1QZW4ete2HVGxEhkn3EbyRWEeDp+PN40eAKkuGOWraNDUy/
YpLVkb2DsgjmM4vttL2pOKVNNaJKAW/BgpjPoBIUWrFN2c4xosr6PrAr2+CB3Qj2
lA5jThjSN7VYhV/cVtO8qAzbe0UuMeUGR+B2WkyW3yRL1Nfig1nXhyoELzLvA2ZM
1Y4/56jVZK1gkHn6JY+dhh3qEHGigLDJJ/ufBisGi4CraZvxgAINNCeEjebGuh3j
0oj9CKzVrH22jA6GbydVWazqqhO/Yz/Ea5J6GCeA3dDTvMgwAX1D0YpwbYo0M7xh
o1AnZnMESI49uQFvA1Dh1nfjHSuzYeSmqQ4jqzwLcpsZFzB7Q6N8iBI4MA5/R4T8
R9bBqIalVUhilZxxMQQ9l0JG8niVZuQpaBiokrvLycR2h5IRfrvGdNZE4/+bhtou
SWdheOun4d6mr/Cp5HeuLyiCspr+qZisELPYbzqCblGBbW2W2l/MygEJdPk0fzuS
tRL7YaAHcknNaX3BwLmsnSttt2vsHwhbb0iCP3Ji7BENSwgqevzhBfLIo+jHGtoA
qj1xacVJ5cM8dewrF1OC8qXKQvB6+Y5ZETkTBddDu3fYHcs0UyDkQRDICTxv6c7H
6kVO2z1Vfcja4Y5HeLb1DFnITOrsESgVCOZzCMfINHpL1ZC2FvHGv3QMY3Y4WroI
DIKEQzP+OvtLMEPgllKERpa5tgDWpKWiaK+Px/GKuerHKNCXUHKw+m8so8wgB900
PM4Tf/U+3MrNY8w6Ji76GTTGesAlSVq75kC3VCAfFgJcuF03vPgmpqDwOTr17cF8
dJ4SOsCXWutqU4lLupFMFXYgDN0cDL06W32axB/2TJDF2WsY7Mj/L1PZY+8QafVM
G0G597KPOBR/Tc2rnbHYgAS2PGNvIOXgNnQOeQjLpLa/I4y8qcdBWuZXaVY0QDf6
ouJU+jTjpG5WKm7whpPOw31vVCL4d0gVtGJteYnDTfNXadvHW/NrG6YjS3c06seR
s/HVFHMbF7Tm4tpp7KbKmu97PAJGVuD7wca4uJvqzuxY/Z8rvlwMe3GLid18881g
Z9wzRuCxHK4AqEoTvvDocmMvt60WlTnMiFYsAfhW+b30n8nsb3uwz6UhIbZJVMQ4
wxfVkQ5V+QZwkhW/BctZTTwpCEWei63kTovMo8I/Swwgv8ardTiXeHmbFn0FXyAy
8aGh3j0FFyj3SKR7bLuoI4PIMy6kJOzJvPDpAFGAH40GEVUNVACPjQ0CPR06g8cv
9bcLN7YrCJGLEWtL3WGxWFaBHmufbkEL9AcGbIj5BoZwxNohmgmcy5kcqklBmVDf
fvgR/iCexzpfqCfG+yWEfQxshHx2O3i/3YANBoyUbPSz8Ey4L2+dTWL4w6ppuqRU
xWiehYzV7YKJXcHw7f+mKVrVxbraEz7Mf7owySpI0PAJ1m6T9sWtWKGKBViJ/eC1
f7/5yeIPmVo8uJulNR5wPe1vKWlK4vu6c4kRbD1z9Be/NHHnIeM+1JmuxXW+oZOq
CAdJdTfaknbhJ7YIAHTn6tiSwxCkMl/9qMb8pLWp6SXofgteWUzYwSRqNPZY0xXX
63vA2BaKNXA/4iG0aQ29LpMCNLR7p1TS8IywUVsrghm1E6dUl6hb12VzrcsT3TAn
BYOb2djBhLMxRWXyr8S9Javufn0UcwGeacoRnTYnUCWFN6A3R/fw9ATUUCfaNvLw
i5XDOKW1+UjjPRGMP0MOGg4C+5lewtuDXpV45iV8i4Tt+C6g9SKFxARjdnbIqp3d
ytH4rmeQV1zMYrKd8ipS5XygipYybaMxLsMpgl+r8ax3vn73eILXCDk75Hw3pGw3
SDDbKRSXVUurhwjkEYua8mQ4YLZqTVbVdC5NTfX22Y1kzSUf5c5w7I9VZcnxJfnP
IXToUzREl7R4oSz1q2ZuTnLjKR/Dl9usiqHOBzvF9piOMmW7tUSLRC5Rc6y3UnO3
q9oNqa4gyWo19wEwV0uIXoPgtASj2jE5VxTZrpOE8JThT8Y11OpoAOmsol34sEnd
ghOl88NcpPtxOaoo/KCkFx90ukguydgm36mlVmH12W3rb3XlOPnlvHGCLIaQhXN/
+1RWW7UjRdXvVB9EKlPiThJRgdLkhBOUPUoO2df8V8DPJC8yXaH3ptugUHAwpkOY
t+veepTv7sqZMdA51mWLj1fgTBUhfIFllwXr2/Iioq9QJSSBNfu06c4SU4RcEiDC
7aqqrX03nshqy/6WoJyvcIh9KlZ+N5vCxEyqZgctvMWZgXkdKu990Y9U+hNEmo6O
H3IrNGUztwLMNa2JJeaApfUfYDQBDl/TGJvMokUBx7X0IYPrMGBuyP9g4lCCVf+s
Xl44fT9gCrBla4jaweSRXCt6dWAxzdLVGKNkZ0kg7MXXAfNjI6xFvnLxdf5wUZ6A
DPaiItHhag3fi8JYhr3sGMxFO1XBtPfZPJNC0aGh6Xk/iKduuXPBPEav+OjYdeR1
6U3UsPWYLU/ky+sqdqfCRmbrtT12VeRt+br7HaWON3DWQpxgMADBwoJSGKcfI4H6
sNBSH8b10TjLPU0l47JMuM6jJwXYiDLxMRinOi/WwoFxK9P/LDwpBXpAJCKn5H9Y
Cox9vNtoqjyRDJkWoNnu7TPKZUwnxt+DCw44qg8qA92JFka2NoSx1Wwb8lA/67o1
8JqyN0X2YqW1q7xYRlDUi1hQS73U6rQYkl00EjGAlQguOnqwaNk7MzukrkqGS/lQ
YiVKv9SeJASSjLJPMrndXwG26RT3KLHekvA9xUqLclY/rd55qlMeBeWML2OKVT4Q
ULYNBmWYa3/hWbUJmIEmpu9fJf+1CpqS1jkGqdexuNbzTvu4IRAkNkqLDO+gkJXg
weXuSAQP888fPKPnr7PRIqKuCOVdAVmUwQS7kaRDWQKuWHo45VcGa+tiJeokSEYi
rHE1fpMuUtuGP9od2ZsLMdMDx7lPTvkF7Iq+f2Y4K8/EWHQC0g52F4ejYkt93bA8
vXVXboTEF3WI7JW2OUW50bJhjwRN+wZS18jTt9cUWIr8JTveAtyBMV1VkdikcE+M
2xDaRPRE/wfi1ZAbnVqa757O9DDvAK2QCNWUNRnhqY8+UhUmcadAgPWvjcfxSavQ
GEw0GoRAUi5mIwxRxdM2FrVF/srFEna13tYaH0i6LrVdzcCrus8V7waNl0dz3oY6
yt9C9V5brN1A4rj4YO/BT91OhftpRaiYFYlxsECpOI8Spd9q5kxbds3ZhSp8jk8F
EQMkroEH696INNRjw7oufR1PAUUBXMf02U8qZ9GKQc9blI66UCaRWgoA6u/sHoAh
rb2BtBV2yalufkyAQV9qe/O5HxEl5z3hsFrj1qmPhrFyilaOzKKi5VDy2jawUomf
ktLKrHFihxgSxrWsE4/rJ0yuqHdUwwQHmiRjlew+h/anUweT9d8QxqKvElzjJukN
Px78l1mSUwrZDoLKYe94+MUFfZT4K4hTKJZGIqDoHZQ13Y5rQp5v6iVLxceI0534
mGeULMhSjBf20es7K8PvlAd5I4tG3TdS1uVIQkRmJ/gTyd1eqoT5Ss+w7bx8fJ5R
K2rcuaGdSK080blDSH29KOpP59ybi7c/3dqLWOc8CBTX9094CoVYQ6opyCppgotk
M72wWlrNiTzHEKvGUqwBuBhKmxnDbLr/k1ArmfdDzGQse22wMdSseT2250pRPY72
xHD0d/Qngbzkq0AsQ6pSF/FvH5fAK5BhbwnrmWcqGbh0hpFZfXvyUhrKmzUuPfV8
iesrn4+3zYAX04NAItULam8BGjGZKHIByfODwZ2XQLlrkeE8xH14Vri6TaZ404TE
OnpzYXK3yleOKBklBgSvHdiKNJM3wX47hq4XX+o1D/+2U+uBN/gu+OCB3KuNDVY5
ZcbDz0eGiZXpjUFKEsyIVozNNFB6jTi6GQ5ivgwUtkqQm5u0fHuGPLvc0eH1tYCK
upulZ8RKP5iIIHBVUwdd62Oj6qmcf+bc238v6ipTAviIhxBuEciT/t12DWo6nZbX
iM5cceMHh28CDJbmIsmxCCwAFTWSzH/0/2vLl6jmUAjMltfiituxtyc/Ytm6YpPG
iXeGCeMmMwR91HamT4r/w2tzWTUWZHcic+jCrZcVWTq4fNY6J2Q6LjRFzz8IRvz8
EugkFI70oOVgycKCVxM65fse2WEUEBOjvOPHtWgfrS6GvGkaUhNpOf+elcejLfAq
uvvHkY7yLP+no/t9gQD+BWlXEk2V1pgbQQYIDvdYVY4eP4eOJCINEYc2yeOTit2c
8zayYwtSkxvsiSQgerkmZYDxyu6ygfVeeB1NTpeCxBQtUm1wYj5vY5wiSKteTWd4
6vADU5tTQjnfjqWPe6f6n7rPuxq1lqjHIcc6LWfJ22ceStQbRZGOj7aXCLjMIOXf
ijZcMeK/B1QOLQqTXTdajrqvjBugTPig6D9rM7A4nuKZEniaot0sc9/V0HB5HsF4
KnUmWwkez/KjOPeim74tPT/3GQ9LlM6GmVF72g8OeOLgj2/6CSR9zwFqAEgCrh2S
HiEki3O2BZPVsZePot767S6Do3wTCJkuKh5BDSz0Pmwys8WPo19l9+A00xRJF7g2
Kzorlq4jqZmNt99RtPWr6XXivkBwAZoRC7zxQ59z1qglFNRz5lZ0v6ypTpExz92r
FloI7cy/KL7cO+bpVjWDj4S6G/2l2ZYTBeNEj1rWu6CejEtT2qH5Xr1LPNUNECTJ
Ki2MYKHV8uGrO+2TKFfJNiysxft7rfQQcMkQTHxoPvvlZarTCMBzKqK7ojt8iHKj
tmb6LySYkXvHNfQOtqkqUYM4dNXzzRLNsOwwL3iKEjZT3cRKAZ8XdeUZ/Rrl2Sad
QL68beT0lg2jhgjpfrcm1G/qdJ+8IzKT4Rw9u+7BGsI7vSFGc2vxEs0Pgcch+Ch9
rXaekVeHCTFPA66YhsjEzxvN2uW1UlrLtS51LqbPhckvbD9HU+mtW22j+gpMGAWy
faIohb28D6e9+FuBv3u0wPU1v+n3J7da94B4Dovud91a4RScenjrc5CR8ysqH6In
dSDazVPt6aFJ6o97qCF2kOLw8ywW+bzTt6qc3BC4gaRCTTUhHmjXwRTnvf01WeX/
`protect END_PROTECTED
