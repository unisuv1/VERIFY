`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M3G5B1834BrrQ1PgLQ9z8e4HBOCz1uLrXYJfEgVIZ1EMyY2um6bDdsxxYvHq9J3J
j5fwvBjO87CGBSBdQIMJJh+CXbZJo2YlVxln5iXQ+6CWp31/L5Z9icA19Hka/lP7
7aez8XeeQVrOmj4ZWTF6X31tdAYZM4U04L/0XDslmeUWUqANpfZSczjiampn2U1l
Fg7RK+lPBK7rvvn2zSNodxW8Iq2hqsyQrrqu2xqyZ1qr+X1DT99MLhhGP0gpu6A+
eyk5GvypI+MxvyU68xDzltE5rYh24Q89LxKWzo9qfO1VAdLLQSJiiEYbVmJxLZ2w
Y7HbdJNLl15IKv0GAtNfVuJi6sxyQ7wxzQaDytvJgXKuZXld3gXivpyU7tK51OMF
Y77Pqs21hQKdee5AiUNfrGt0d5cbLpKN86+KVrdixd/iPIIdM4l3vGrP190Yk/rq
bJUAzSo89+TMjcu0ef941IMM7dxAup0VsslLayZATOiLqQXXthrWhO4pFbW7z/uC
8eKAIBNTCcp4s8Yj7eoVzMHwECVxkPNsQrp34Ocu95SkRjWJN/bmiQ2qH/w9OiB5
SRVCVSqaWIiR1zxbWpKQ80h2FH7VJte5NjSh44cnRl4uYiYsKxz8SHDEdPJGinEC
tnFCQwqOvJgXQmQ5qIcewoLVR1lhcHcTQldV90BPs9MsRmR71iT8bnFg5nKUg2dM
P+CUsLAHO2SoO+M7indcI3yXv/vxoaWcFxHKmjzauOwElSQUxECCwI0bP+eVzo5V
xa9XvMJyqT53BYgNmLTrFuMECGhtIE+TGvIE42rZBXDvNmhVLOw9J4fkxbckxXnp
8HqHaRaqEyj+/QP/11W/cf2fw9QxX/uiiv8Q0W9BPWk9iMXUVBH2KLICVT3hHb/k
JSL6mYSJIy788XDp0NgvxK+BLe1gofOKV/6cE3ly9a2l+7BeCXplmQ0TisFrSEIe
x6ekjRN7CPopP5uS+5rE/YafMI/Qaw2ETqzp3rv8A3Pbr3nppLVmxWEFKI7+omYX
evs7d84DBLMF6YCxFrwQ05azQxXJUg8yJ8/H5FVVfCL3olNc3CsxmwqlxWtk2HtX
Z/6sv0g0umLrzrRTIxRZiFSY1EKviBWxPYcj9lUTAo+BpyaMlqL8lWyJ21+1tbTf
/2oDCw5wpa7r00F20S5xXJfaDHatUAcHU10sB3A7+LVI2YCQPhr9DO398DUWmmct
2YAosDTUFzVPva3R1ZCiJ8wZ9gGIZKOGostUf63y/reMpSRRlaUMLKbDyXdf8CUr
cgy7tRN2BVO+j5iIny3QJ88uhV7kq6jujnfoXtEmgTJ6O43Jdrapg+Gtge7MmJia
1Yh72kZ+o/CXj012NHOHXc8aFtKfgTRJ0gv4cxHz2lAq/xaAASK+TeuIHYjQpk0C
99yqGcb54zzlR/iVtLoqCxhFqghLWYOU8B9sJ6nUmNItwdtRN0HrtA4GOPjeqLIy
W8fdvQEq1rIhSzxkR12/d6+Vvv9ECgmhTv+N1tQI7htSy1TOUBfehG/fQ5SRTV2G
gmpJLl4BIPwXuKOwSaRQfWuGAkk6BH/rtS9XGxsC5Iq9uVdGwe4rDoggmUpLrYuE
gznHdf+pKanYm04C3Aa2fgQ70VQ8AYWrtN3V0YD7EqhtRoq/n0QO5okZSXCoISgY
i/ssGgQwCOWdiagyRg/BYnAX+Gtx2ZmjowxmpSDOS3o4E/F3i4s2jiK9Z5AI/9Sk
brZUm3Ct3WjHy+PnLE2RR+Byf9yF1WxWFNhyDJzRMDCM8Hxrx47z//WNNcnTTai7
gt37ccC1+Az42g63DIHD6Pvt4Vh1VZe6lRupltW2Kfoqte1gVYnHEDA+47PUgDRp
T+pnPu4F7dALnnQIGulQWlCeXXyQBYlTaizlRSRE9Zuo8hU6ptIo/fkFv6tVIVpj
YKuX26V2jT9s1js57E8onW8V3P0gFWTauA3eV9l+B5eYk4YreWIc92g+UE2d6siY
9EFlPVOw3AePKiK1Uran8LYfHnYLsvAgl9fOjkgR5Fgbjw71IQNNYyZojIuW1PGb
s6PGQL/WoExbIYe5FoDsgn0v1q+2Be3bywP5S4FLjyzbvB5kBOQATeHpjlR4GFtY
XNtgSOoBDLEXVqy70I/U6y3TdDiYzsZ30DP4YcvDifbBZRRZ3/U6QuyiXBoG+hNZ
bUQ78aE5h5PZZ3y2ga6ZQqm5DyuqQk3b68+nTdw0Yxd5ksYffqdv66iwxiSQY0Tb
LWWgKW7QHI333OJZrr7E40SU509YO7OiOyfKfKQC1bQLsSKtwnF4kWeDFPmmVHQz
pZKO4Vcitd81/h31ZSamSitLBoYPjB9iJHOAG8sZi7CgOLvO8GfGjs6NTmhQCyjC
ZX/9gOyDYSVIFkof5uwo6zm0mEatpuTAwZHazhq9CrEOVbs/Gujk5m6bDc2Imq++
UPqXtBxMr9g68gZLVBO62KXah95uxVYk8kL3mAfEDJDUd6VdgG/cEquQ1QvqwyRW
9fPEQm5CyhIaN4hoKUp63c8v+BKgZ+wZqJUjH/9DNqkQsDlIJPD5UImBrnMftjh6
IdKWVYcNVOUjW6fWoqgylelW13GRAiWISSWrBO1Befl3swCkKUqlmwZUUowtGcVj
3w2z0KbfQwtOHWnHtx3XAsSebJxDS0dVTfpNoY65KuSTGD+vmoS80u66z26AXkfC
zN3NBrjHyi9C6uqOeBVB4Wsg8fm1uLePoEhGrWBepOIkr1eSWOMR3oDSc71XfOEW
zFslR19VBBXUYoOaXBwZcMgD/doUuwQA2P4+s1gCQZuykCf+O2rs8L8s8nrnT0gS
Y7nJCs0pzOJ7IJ+1YsHx0IX6Nx54dY6MVvElrm/Zjv5jYXUK+P5kuCQiscB3wu8H
DSlbQmg7iVH5L/zAFNjua/P0Z8vKLoOSpu2pEAtw9obCLeFGOyn5fBjalgFvPaCC
tgwRQ6R6q3xfjM5aLZfx3MjjW/Qfq6PR7fcnns1Z8Xp1g8CameW+935kSDU5B9QB
qDhuL1OusHhJ7uuKzL2yccGMD70shp405+hdFBwKCnlpz8HbMZryNlGNCQg7GnVC
kSxzK5v83aVXNa/W9CzdaSSmHdKbMHRDHwOTKgUQyseRtryn9bECQ1hMM6poAzwg
dKXDoKcfS/FIHdw/FNpv4S8OAC7qYtrN2U2J9FXkOB3qC598kISNvmAowyMokDnC
gsxjqEPts6sRkLLOR9obZyX1vciV0w8SRF6+PdiwnB9fmfXyucPCiwvbvW+JEEGf
g8+C/F1J99a1d22YEv2XxZfnSosa67/7XU0NlHB5M8Y+jRlBvrn8ebrScnsblRBf
Dw+LtJoX/KU3SmMROGztIwfkwcs4CTlcs3AIZqCWXFNhPBshHOLzI2Nv97P6nMT2
feBtgfmIhtFouKHdb2LJ7ldiza/YHmJxf4C1v/zQy29A1In0us4Su2bw8SnOWd09
4qiJ6bZONeYvDKt45OAH8Ug/Q9FD3xQqR8kqTvq5efrH5llGoK9wfCMMe8R5Ddqt
XWKOZbSOngkj6vig6FOTKlTo2jds/Rh7iskrVXC+SLV++9Ys8CjE/YMX/33sOd3B
wjWcHRr7fdc9K26CEUUNni9WrBmcc0EEks+9dois9ku3Bn62+UYTASQmzCB6CXMg
LFKog30tJh4oEQETU3hlPSwPfUrvj36Z+1Svco1K0Szb2Nf5FqVNuyd0aKLEZXG4
dGJmM9umH11QjZER0kKESp9tdR+biz20CShPelSyInP3rEKOIrAGGCwYHV7r49gk
R6MYcNw3KvlP6XluSeK70BSVy6aiK6j9uX64ajAjHtu+zYcIBUrFlUh1FYmu715E
8wB6pWXfPKOvmLOsrEiaFgjEl48Mb6VsHlLJb+c9IbX8tVRjSts1e+Kez1GAmzTZ
WaH0FzxIc95wTWEPUKAQDHVx75UbsBF3T+2TQ8jFX6XEUqhVAyQ5rhn+aloTjuEP
de53sHzOJDxIbcK3nDJoijTgyL9teQvFj+U2CUpmn3pER6+yDnPFQvAJCVImtOKw
Bj7q0yzhyCVXSUt8UwevCE1wtTh+R2g94JYgFF4XisGaKGKGNTz4ETlO/Rn7NMZg
kZZFG+EG5a4VDE8SS7sSCxOtRkbaF2lAk9nXiuiIpL2A3WtHbe+8OBf7lROqVA0X
9hYBD8rS+o8Vywuln5TOB9q7BiSxcQCXclV51pajG6BAa1uMyFIPyAqOuQ1kjZOC
iMx4+ZX/1AC8a4tp2G2bKLk7ABy2s/EQdjDOvGZAEUVhDpQmH0bPAw8lMbAO5ruQ
EkzaF5rZkV57FrYfAESMUwUOkBgwBCw6G5orQZCY3V8t/bjV6ZQc1IczfkLAv6Nz
73u9ym1Eqv1nmD4k9n5XC2zyhPEc+7iUeSBzSii4a5ItunMutWU3qf4HGrHIz4AB
OJm19E7vl1nbe+vqJHf5JBZHtAogR9b5P1D2I29S+D0f+o2J/7yxB2j6R603Jby4
iLGhxGGYrYqBBzUsJs6mZzBso1/wnlPzvOfukZxy3Dw/9+nI3w2Q84SngEnO236r
pIhfzcJpYSYat1PfY4KnkWilNXBzo0Rc283Wlh0+GLUwDxLQVB3+7gMK9s8WztgT
rBIYjHAZCoo6b4xkPl82ixw+1LfsM4E5z4umnJu5uFO5BcxwGeTHKaqqW5rTh2pT
fiNPqSxcuE7ia4ww2cvFUJzjDJcoLj1mFOvT0l1wyQy2lE0DsAJL8oEphBem0kKA
wabh5ivpDiiH8QXQm7AlMcaWjI42+tWV0fRmDwIahY7K49S+ZOk3fc+SLHDdkeGE
ZeVBATjG0dF1SCCv9D8ymPFG1BIkFVxNpnnJDDGyKo2N4EqrIMpk8wn/8JMBATki
AAvGYaQo1f2CowsOFmfPLFBZ9CUusi/xzrxbDhVQpNUm/OAErs4pWU0q3dZlHTKS
C3Smgxwg3Ht1wpz5ipm7vCYTbmjwl2Kx6ZepzcQAjV6O7dhFb7jjoEcRSm6np41Y
/2Mj3fexOap6NiBtIwyTauDLEvZwn8CprhGdYpSsXxpxoKEobcJVxZ4q/aTASI4u
IDtoMlpspb2GyKz79EzXep2fZxKjt1GepzP6vQ0KCcDnA6LLiKLqiyGcbPuRkGxv
IzlnyOBoD5D5uXM6P/mGc98mmsl6lHVDaVtpjXBFTGs/rWHkvGJVSSKDHct7/aeZ
K+PWRbOCdYDYzGpZqzf9IaF6wN0hDdKjNTlneaBWskFtaGkvAppr8QNIaEQqTMrJ
PwLD55Tqi1QmMMgeh78oY2ugodwa34KYM8+Fc5zy3zQ3cwX8I64BY5DECh9GNInL
`protect END_PROTECTED
