`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wxJREY/P77NLTCL9aI85T2K6q08A0akZBsqRL/p9+ZORs46SWtWWKJXoCysxXX1Z
NdenM6JvcfeSr0g6WXZDP6zJyHBkDYz3wJWT7HyDKngDSWt9ffHFvDSlfZRzP21o
S2kqrWIURGF4x+qP0ZwR+1U4GcBqwv2ljML3AY3DnAvhiyNnWylgg/IGhP/SOVi3
`protect END_PROTECTED
