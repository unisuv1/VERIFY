`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g7y4to93pUn9uPgFlypqzZpZ3AQyrHSbakCpM7H5y1b2FgcQBx5sHoFprEMRhi2F
WZv1jpK8dbkj74cMbJG6GHhr8g0ZnmU3+4klFfVMjff0DHCyxALAJmkJPmWKJ0vP
omi9SocrrOnPXvYoerqgT7hUOo7n1OFF4rXxkuSbms162HBsuNrhp0eDJ208TcFv
HYGJwF72sBDE9UFyg1kdiGhama+7CtxraZumetrwukGBIEjgcJduvHEAnVoAZfPF
Z2VNeeQl+aiqalcDEQIf8PuZ92IB7XuNvoFWhLrO3O/gU/iwmyaPxhl14AsdmO5u
1XbnlsEls1oltSVSRPqR09FGKKi50q+m2t1b+SpQAiSiWz5rZByD5O9+rQDhZjhb
P4AOJyQjLz6I3hfSHPDN4a6XJbUplhtboePrIS5IPAhvbGIOf1ttIpmPCyYw8HJA
9l2jtL+1Jg1EbayomubRV9YsMbFmSrMjjLvtYEFC1WnJRnvaUEvGFiClbVoZNmoZ
ZKNThRrZhCnE1uOdnB5uFYchvREsxfnyV3zbktfA8NeIKe5qIqAWubgo36qwhGFx
IDmU6DrqCQR5NuQM5M5w6uWnlW6LTo5tdcnhYameRkHw+eoqfrBIYQieH6rR9Hp5
VWlGQ1mXoJkBYt3xRVH47Pds9WDcfqWLutCDwm1MNdbmxTpXURhTerRTks9hrm/h
PHXTsv+P6VEkCVADTUPsdWt1Wt/DSD5bW/4QLi3WTdIjaiz7QYq9qRznWy1gy9Va
+DJGGE/S+JCo1pxVpBfhhLykYmUz7RvFr4j0rbEMrRLX1x4u+j28lbV4nUlQhg8F
y5GCguUi8M7cWiX1Ps5EdCXOJDxro3gADJAeLTaM6zRjnACveId4W1Hcsw4PQFX6
IsZ2YZ/0B8mWc1AyBgne3wVevq4g4DvucGZF/0KrA5KOJzjhlrA3fp48ybyxwaTi
Tfcoj/T7X2fqfZsSPZukJ27UGA9tyq2nYzSQlkMjJxWFqGEJaFPnPmTkFbnt3R+X
3NP9ApBz/2XdK+7e/6Tinolke1IN9HCU01W/ag+Q43v+FEWydTKpmwLcXDYnbpL9
Q3mJiLvQ53TGkM7u/3gHljb8evbsI9efDYLGt09ZY/ffufHsGlVMA+oJudsiEyIe
5ZVVxeJEgjHCe0eoIWA2LF8/z2BwLGelCTxMlEtwPs31+yFKbKQokuzJt2F7nRl9
+oC/LxI62yyJBj8lQc9IEytfoDI3oIP5tp6g8X8WBE7fQssJ0526xpzCRM5Cd0y/
zvyY1aReFLcoOrZOPmj8y2AgzIrt4nlNhmMj+skM/frJX2LIVgrKwlr/K6LDFKOL
i7aspKwG2EdM/CVjcMwLDNL0ouUycmTmambo+usSwITRrtgBYQZVTWIowLhRfHyq
PZTChnc3VXxgq7W5ii7FEJJJLbIHM6Iwm1XjuIx7OKYGitdG8Nm6632Ib06pR3V+
uav9Pi9rnUoSpGiykQ6XcJtIhVmrnNv8us50qxpYvDluSttusJon+EWwFgJYyoGb
lpZB6HD6xSQA88cbXknHApM6XRhB5VYgYrX5SlGFbFdwJFtOSgTtpGP239Bf2oYg
7yz5K/W5NxVvMokQQhdshTMgQlAKh0OeKIj6E2Hx3BgjkR3jrciYWA9ur5K4RLVd
CMPIVmN+VonYwWLyVXzMD+R8Cs6nwlv+7CqARojlT83wiayeaXy/ouKCdH16calW
5G72EwVm+vg0uUcHjDtZz8f8rUFP52u4OTSoV9WAxtg1Pbv5J2LsIf1x0DCe/4Ki
7v8Aog9Pc2hfDO6ufbfo7YKUMZnB2dOCZcluC8yyIFER6pUAeHvO9yVo5qnGgG7P
s0Eyi2Z+MD7k03KLkHkkz3egcjJfCwlf29kZEoQdx703zLPFiA1Ar5joe9PT29yQ
bwUrZJ3Kb1f858Dvmj3wYgJMoJaptiT5o0z5Mz40nAhpaAbtQqe28MvRbto74ZKk
oFyIZL1XK29UY04piMjULGd+t0W+X01vlE20lUJEZYQ+2frPtOs3jxxRRqaH+AY1
LnQh59JK4NTOr9IL2eO5i2OI4lz7STiPchXnIIVt2afUzkpA0Fbu4TlBI52GCX9s
7clHaw1j42ORKQaiRW6xQ1IekqclcR0tzlAeiY61GWllV9RE1CHMhJYTMMaQfVc0
u5xzDldhwpCQuMtL1cjH2UKDhWauoJnHwUCMQ9tswa6Txs9jB9l3VU13tVZU6p/E
kfOpQVJVki2s5EHobQYuFJ7dnGJ5xVfrNz8ttwXWneEllMhPD7nWpqMqQV3gN/kH
CXo+naezQqE0Py+GGlvsdnSu/UCZtPEjAsbBAtEP+TnoRb7yaTf5fqDTWHuqEOSp
5ehNMTTsE5KXd607fsi7rHACiVcrUwSt4bVmBCl1Dr7wTJGPGqmB6m3iw+xm0gg4
+Oa+5Gb3eSrnjlQsEHUrv0fZ08d1tJo8FeXI6FpG6lsdY+I0JogTlKnvv6K0bC8T
8yB/ESeqMl/d3VZoiDV7Phyaj47J9a7Yii65TbPN55j4/lWUUHCT1Aw/YXZ+QHYj
arpSEPlJvmpg+KgnNZxPE6iwRJsbLwVDKNRmP8XrRFQHp+L28TkkD+/PwZLrFwmx
yZD1ff5EeZznVo9lEO2MM9db/jSryYX+Urew+0DFQCQ1lpjKy9Grc7dOKaUEw4JA
j2PtToC3NSRfj+QtmIvLmFCZyFrxfi/donO37dEHWYwsujz/ReUTSYPxtSz7mAyW
A8bofacdYoTJguNY/G+9sW7OSA7kpGjgBHpMAmPjs9t4qZyOvVGW1CIZjOxk1AY3
K6iq2135rg1v6HCtNYAVXKfsVw7rvIQ2Z4Or5HSPfDaVeEfVdr97WXEygyiPYSu2
1iB4apNBbh3f4Hm/VxLWcwaRH+OqLNMqQvcozL2ifdVgrzwngQec8uiHzhFDhvsn
YRZvk7QDznLYX5jHXyfnGa+FUuhjJxLozwMQxQ0XV5xB7wS6+x0NOMHK9LATT7Yw
6tsKOuibwxYjUsqVI3ofvzeb2QrMdntXijaLSFoXhV5CuaYljTtERmyr4SJ8i1Ba
83SyFbr7lB0ZLQYYSKRY+oufgDv0Ktj7ALTuYsNK7zVIFV21Q0lEGv6D6qqh7GUF
m3ddWW50pe8R11L6Qj934crLOjD2FDWD48/2ldGDmNOi5YUH9bn+BIa0jzdplzsq
drC3yDlzKPM/yuTWefS5F/Nt+EKl9kPVoz7g+HMi1ZD7waCDlVIKArrKm1zYpzf/
TARPP/HlIrz2n/M9m+adsoTd54obYkX8z1DYTHKe/eS5sItcH+giGbqp//w++1Tg
8piWpoxwnM7N6Wd85UlFSAiuS/QJtsHmuvHiv3v5VQJjY/ZDgucDSHdbgEClGkl0
q2v7x7O4v/dQbbUX7Xw5qGZ3VB4gkzvATUG7W7ydDmBFEhrTaccbLERQrQtddYUN
o9Fz4VsA3ERipMnnIdiLyNO5x4iHot+3e0ln2TfULlxn4uwPweoSsA9O4N25etLw
tr/ceoFaHXGfPzoaHcIm3M5TJ3SUxRYa0prAbUPB/haf+JQ+Y5ohm3iCSj+X/8z/
G3Yb1qazDZgjhaPhU+Of9P0T7eqrIBjqpi7ZeRha310NzufeJATLt6MVS3bvmDl0
I4Dv7Wj/N8rQ/a2mcXeQO+vuHjJtdDKouYOVSwKEjyACG/3ycWUY1Pa4i9xqDq0Q
7Xr6Ar2yBky6jeCoxflu/w==
`protect END_PROTECTED
