`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
HxiDEuIW/bSED2DTh8gujiu8JGh4oQ35vkoHCeYte9Q2SEtLIWwCMcOdFksyrPuC
6X512y36RWAbsiKDQFMscTLePtdF7UiDDdsqsrsS5tck+HQT/Oj+kODUC2gx6UDM
FMe5qejQ0rbxkxNWYtrCwDvz4rA8GEiDpj3bKFohU0L3QTwUBk4q8chs7OmsEK0c
hngwEyknCDXaSbFDk9fRgBoppjy4WNjd+K6Ke/E2HSLHx0caVxsvWm7/rbgzWs1B
pggavf39Zt9lxrJF2XcEeLRyHmJTWcZoQBEL5Jqybye062bTBzKw5ablqPgAUeGU
WyViuTeCTj2ppX/b3zcpkfeE+BGja+LDyu9wamhuUztoM2QRnHr64vZbjXB9kVRT
pKn0aFP4EArtNuuUw4tAxdTpvw65aLd53+fDH6lIShy53W9QIZmgcDLQOcIVxemD
cuTXzjeqCCt7j6y98ACFdsXjqDVKO9Nzy+Cys4u0+HoWvAXiiInrbS/CBWaMWjtJ
rTNZiHvUxuCWqg3PJdgYhC2L4llXccvXzLsx8y6W5Tx4gqMy7qPn/yJHw3RBqK49
9YQdH854FtGLvNmgrL646qHmj73ZZYzkQuU8LoaBPV8r6QHcNtI159KZOuRYo0aX
MFRxhnT/QMcNEc7D81172ObthlRRjNKA4g6JCCSSwLnvPUWoYzFBU++crwRlrYgm
cp6gGPnZSiHqau3ybmBwjFQ5FBehLH8164b4ruLlsIA7wKka8X+LKH0NZng61jAA
RiEx9JpQ7ChV9Kfrm8ECq+egAj4dY150/MyiXMnEJdnC5eIOsuUWziDZfW7wVrnF
`protect END_PROTECTED
