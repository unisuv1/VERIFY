`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
7Bco1uOMY8v14/2/qg0Yl/X+yyzhGJCH8cX3ge1948nKRqtA1aMQeydlHn+qrStE
Y3Ajz3NSOcnK8ycT42NqezEIGah4rxSNi4+8umNdJsBITNhXDCac4k8mBm/+CJxE
UxxdOI5cNzx7VyvWoWOOMyy+yaHz3HbB4U5zjJ3NbPBVXPjK84F52JYHptI2Crph
0vCkvPt88LP3ZKD3IxBmQfNFnDEg5zaTF8wjVic1OxQjxorpIUdVhH5TgFxvsuyB
72Yge0jUVcXWh6S6F/ilMBS2o3bi+FcS4LHRMPvxU9WiqLVtUfNCnrk/KF+fefPw
knG+3/YDIBbuLqZ34LjMIzoPTlfwI3wc6ynkJja0du281c0VZ0l2lG+/7btEauCz
VnsOJM2Au/n2dqw2FpaBrbwbKKmijm6GF9vNlrp6ZDXS5YCf+ykXk/GXt8dN98hR
0udCGo+av4b0vD7xbhMZRdqEO/3UgrHMXueN4lmiNUk074/2kSyA/I4lUXj2784H
9mwL8fReorrd0YKnHxXgV+zBWxiHmnVCauwj/+QFm4Ti+IR0dVExhC70UiNcN/1w
02yhfHL9xu344QtV/TZQKDBizldR+m/7W0ljNXjF04NSz89j+Nzh+KsRra8b/Uex
eYsvGRak8lo8X1rwQxsgwL+lOdy19NSZivxLMPbQShYOTeQZQzLPBbqXW2rzC48k
wtBX7oo/XBROQ2aST5V+Cq8i/NJr3QcIIy8d0Of5Eo3lsR/tOb2uKwEBDHz339Zj
Tob7vik0UCsu7EUNzv5S4tQtCDazVutOUjxG7YeWvTOkSFa1QysnSYUkxiKykFrF
0Y6E7YOWNQRZ1qulN4kmOyCoQ6MsarFdt1CcZZ3CZR+PK20GjUJgybVAlHLxmIHq
37rREkP2ToxvbuvuQiVfnWkEtdHBIybUAkkiSv46Pki6eDYqECNrAoW3s8ej8HBo
uXMsVGhIIK05IYixVuqGnD6qb3ZHEWeJaIFWaQ5H1/+okhxesHxMSLgvVz5XbTIF
P3141GHJBPOI4/P29zV9u0V3LQ6UYYqZ3aEBhkwIdG0kcqVOyXd+9bf5pq9ET3jt
EBb4ltumoTL/ZP+o8VDtG4Yyhe0z1915xTnIW57AeXFHUYwvCmdQH6f8sPUPpzo1
hSGf8nu51gm1YTSNkm2b6WaYmfG7v+ilMxQK3/rGkcyzoVjlxsvIUGxSkNwg+NiJ
ozhJ4C1KdXhwQIxZ/3QAGpNE//h9u++cnfJADunJYlGXe60vTEq5a6KMjpUOwQmj
B6hZdDZQ5UbzT5o3i+9BoTc/rc8Sd0Oz0LhSvrBo7fm/s33q2YsomC496mfNAUgJ
MDUtc5o9ZWVorlmeppYWN5ViJ5sjWSYjBMkeE7vCHSWEDJDtkDtsPLJxb1CRkRs6
JaLnRoBbOl58mg9jhddoIDjXt+djrGbva0y97R/Bc+Y48ON5lDU6zJmsmP0PI98d
FE/I8qUoxCgjfjaiemXyGu42Qu9VilHhI1wa3F1BDcyh3CSwHCUdrvtkoPBQfUtw
cEuDcI2AJGDjm43Od4tMHRxcXqxl+5V5+65zdtWxkVENireEUxl7pfxYZo45NIIy
g82WFFLewnmpXvWyC1Fio61GuFG033Li/Az5xBorXzODBiIST1qaTCl5b1JUXsbN
nc8O7+vGEFwYi4oysf5nn3FIK0W1haWqcv+32w9v2HaF8YcM/Kd000BDp4DzeZHd
mMWymJHyEBBQ4IJ9hhCKWoNl/fj0XbPQ4nhJzQylYBb7BWTiGHU+8eRao/6K//Z7
`protect END_PROTECTED
