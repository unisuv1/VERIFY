`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0y4D5CpXLRnk9qhyYV8b4lG3IwUClQ2LEBx4k0JrOeG3f15gquShsjysGirsy5wW
O2/SSZMvuhyQm//fQqifcoVheVIJhkP2wCJqmt+gUcjad90svw92v3yuIjQeLjXi
GFUcoH5rwV54MnE48b4s4y2YpRYNmKV5jScFT+g3/kC0KbUQyFh6TOpLQyAFNVa5
+olQANlkGMAvetkf+AcpEcioYWyj9lLLgvGPmvmJMMI/D4y1Y3S5ZpDWFScWzNNZ
oqroJoUMGxAKOJJxZ7o8dk3qnsrw3icddBEFE8ykjj+Iz7MIJBIs0xSanXudriB2
uY9Yz7BSfNZmvD0ZSfcBb6mecC7OEAIKjYYi9Ap411t+ZYxhRE51ZrCmyngqoiEk
SLHYCQ7mpGeW33ltHkkLjWPNYIRMFdIV9qUg/MZlii7dA9/oo7aBRwsCtNHWGoSN
3AImAOaHiXmmXRUEbKEST/Kot9mhUSEoLZc13Om1pklzftCKyfoCwAFKqM3vsQ3w
+UFc93P3rca+TnzNNvF2/JWxYSZ/m1u52CAu+XTW1wkK4J3kx4f/KfdDxFarRg2S
oyd442XwxTHg45dJOcX50IU+Va4vBUM+lDi5vYLZaDCcqNE68OLjHpAZBzBBuve/
9HpQygrF/ABr6r7s4GYYr9QzVR3gyoSDWSAF6wyxnuyzmzz6h6HhZ1MChTNuSjlt
eZgKpghAbKL6gNziRdTnHvyTRDIXabZXgJZnPBZEfvq1pWxYJjc+krJq2FKX45wL
nZccboIffFPz1egaZKUDlgS9uCoL3ioLeb8WB7wr6DLSJ8xpiUH+Wtokgrwbya5I
efn6RZlaflYZR+gzrXVfwpsmWGdshnrqxArPxdOf94WmxByGPviZpgsGZqGT1pIn
6kPhbIvkK8bA0BIF/7Hr7myq9wliizcffcxBvdYP6b4Jr9M+U12IRixk11T64gqt
Tfh57WF54/oHGWhaJdobjJA7s4Ic8VhC7Pm0DDn8dqAvi8zttGgK13yzPNmXSh5W
9U8fWEaOT7xV3CDFk5HFsT4P3Sm+EBXETWicgty2k3ZiYwSe8T5c0jpKKD1a1+nm
GPrIGmJ4Fel2aPdjYUhLYfCCS54NM1nLLNJsZauuraL002FHmC+YMH7IKoLUitNX
YuWaKg9i9Mf/fVN2qUojyd1fg5SI/uaSFBgpVoLZiMxKZ4vjBaj7256SEPlVa14M
bIznm8J/dqXL2vmmPP5PVlTW66ROonQUn2eXzo/OkBqdw7kr98QUX1kfG69x5d7Q
jaEqiDuvQHmrp6ubd/Pprc/xrtofDe5GkzERC1pTD8HPLixDjkeGH2qWUAQU1eI9
vC/OrTFlbQkdHBEf7bVKletrL9mq6SpINnfpjjefoiwWvSO+Sv93CQXT8s+zbHzD
4BCUfz64xEux5WIKQurh7KEk0MMykh8/jVLz9OeXOeRkGh7ey+Qf2DrBcIysMvpZ
qVc2VRwhsHQpL7VIikYvh247Y2V+CZ0IbJAnAt7s/JSN1tc8Xmv87qmqfwZKyd/b
M0Ki69lZayc2zwWdOjIfWA5/vB4ELt+mS0ItvYzFmWBY1tFmwqxDKwjSuHi8Xb+U
7E9thYVoIkIRAiVMIPFNyJpwgq+5mVupk3/pd7YHjWJRSdekfZwxmfCbWBO+osv6
40SZQrvmrb31u48TvqI8oqjtG5W4BftLm8OHvixNAaeSOVBdbzwpwOofRoa4Mvja
e+u6kbfjKjGIQ52ELpBqdA5ka7mNVwAfFMAHl6QD3SJ/NO8IMV1E3eKdf1vOWy2V
9lAMRBZ5eWoUg+PLjxJoIeAZIIAGPEu0IUNeRl8V/jy2FX4/tYOJFk89ckyopz53
sSJFbdzokLeDRJlSNWvj687RaoQoE8SpgmnBeQh5k3WtQI4JrVbx8UZgC4maB3Vh
BCJg+BMM11khidh0AM8V2MaUDAnwTCxKRcDXMsFbJWs3BomiFQcGob3fcLVjpbTP
2FiTooyxMLfHSm4/67KMqtKov4XXTbVhUAZZaYsVDcVec/saVJP0oylhGVhRhubC
XNOjSs+hFYdETZ6li3k6vIICm92QJICrUAc2ccge0Zd3Wrg2Wwi/8cK18CQMD+Ps
U6K4UtmUZevHGykstL/n62iG948/mfPmglxIdECutx2qxOJC0Wd7ib2EfQa3b5mp
zT/cpJiVNHC9VcviNmAm3NjutTCJKIrjE8Wk1ClRfv4h2La6MZiVXFYBR3G/Z4uY
hgoLLN81RuDGDB20Kiq5EqrkjFe3GMYdEtP0zXIyvZcke5OeOWdj+C83mDhA5n7L
8OScHPuQmfZeV8tvSvq4nxJfwR+UDK0J1dyoGZbxeRJ17ljLLCb5fs/API2AY6jE
t2y0NZsTLXhw1TU0xRqxeTD+ieXA4xPOmoLk1VALKL0ru0RmAayhrAnolIzkiJLC
hxdCKpCMJXZY3kL+u0pPQASN9nCDsiy4m+W7dinqG9ZUWbKwnVL6ID4llleVBoaN
NtHgi2aFMvxRW9LJhJUOkTxKdNFcCM25at7I+Nq13zR2P6305xhWZbPGRyzDZ5+h
aWzBdmZCF8O0FVZ4QbpS0DHRpFfcFPkStvD/p8mF4/zuTxb8hqY+/ZujBKFYcDLS
5DOv6gyPRA/SKlCXUgBH8Df5lGXP0uPGQAQxbuaj+QA+Rb0Epc+2mAnl8MV66KDn
JHNV/cP97IfaQVakZBVJJ9brRnVUD832DhRQeti5kNQfydlKQYke9U/h7ye2QgW/
/NSr86GRnmu8lsvzhwm5xUcu2OdECjG08N7U6zrU7gIgFxY6EzwvOLuMoxpf8Fv/
6A/UCTZIDrtIhf0vEzZm7HXj/ePiuJ8wZkTV8wT6gQ9Rs5f3hhqlJtHAyrVeJ5qz
vU3pBjowqCTmNHwb3aHYe+d7W7y6gxLkhhW+trfZ2q9cUmuBTUlpO8/4KUnBlNtQ
pJIgqiMek72qZD4a1H2+noyJGwrvLZJ8iIlCSjDmYnMFXb/nb9P+6A4F5SF5CGjU
v/Sfo63ySfyQ9nBQ9RXbrs2EjYx9aj5IK9L3BU426QuDqeDi2REDC5iMrLGl6Ij+
4XEk75TVShFjC6Oo7RSC7WkuOvjpzoC6FEVCv4OPNGK0ZL5krTjqytARbj9rY+Wx
x9m9KyuFBx0xkj7WaRvIDHGuM68XcpHWNwdtrLUR83yNMRtHVPZCaiUEHF7btQih
DrvhZBTZsyaDx1GvUjse+DBiz/glFYYevTITfkvXFBzvjZtdr8/nM0xaAOctwrFW
Oy7YWO0Nx30cur7efnJ+HbWj9CX61dc4c63JAvCGHpzvmJamWx1FPmiuNAtS5MQ+
8CVJiiG0UK0qyIbVb89xJPUTmy6Jvh4l8IrAJncIW/W4kIT4EnqBUNkNksXCkqfr
9BgEFXj00DYY5MP/ChIqNZ6cMVR3RknBlozezPxI7ke/IzHQM1zagqx2QfLYnaer
Co+7auNQAKTcokLD6IE3xZNl/awCBC92zzmu8DKt0rpZO5armdQPoGdc+ngTgWg9
rgKO0C6WObsu7ZZ3JFsWmvw85oOkrjCTB1TQpcMrFRqM6U2X+HbjIDRq+hPIBp9l
uaUhAc0sgCI77P2hjxcpUg4PtEdHVMmo3Rn528MS38a9OFZBtj45WbI/UN2ceIHl
iRjdqG/oxSnD7hf0RjaX8z+YEuv7THBwJXhO+OzurH/uwMVimP9g723O/AojGj96
mkcj63kReBM9e/f1PCQASJ6khVVulV0EAOqxtYS62dfFOnzQ/qAiMqGNooehg9uG
cNHK6LjbgtnQT6h/0cymHTTwYJNFoLlmvFywgr99Fg+O1u2jb1lCudX2GpjkonDH
j2SyHgUFsi9mP/Ki9BhMwznPbd++JLy0nr+GWxl2DUzyUpcZH7nqkjs0A/fsursY
Ujz/Qt8V8NIQW3HsCWhq/GInWIbaad6iHvKGS4bxsRpCeAG8Ngpjs6MReVenaW2q
DTHXjtyUvWqXLBmqQJZDxe07aCzUD7c2y7EFUv9QwAIOMdO6l/JrpW8Jg26oQoLD
FUPEBZVhNAYnVlDIzJSmL/A2h6rfxFvXVS6rj1SUPDVcVCEjMzaaKIO57jy/cZcK
3PzoLtQb0ctAdlQIFAmaky9R59yDPhaeCDgIDREFuP/FJ0g5iOHNNTEnRWsHTZYD
nHvaY7LNiUDTll7wnHGKx+CizBygOybztiwGnL6ufgaSvtWGnYSF8qga8pQRJQoz
EREN8pjlbUnyxD4tIGZva40SUBoMQyVIj05c47ZRr3aO0EMTFVCTxGREU4LEyDKo
rOgtfzGtJ4S1UOVxEyefyzTJIgus1B5jHpKsvEflU8oJAs8H6wBcu130weJ3r5sf
IDaL9rgUjvO/TyT32UK6A1MUHtf7E1X/NrkJWGxi1W4/+T+ArR66R9aWzAOGvMzW
xgnr15PUBEJsW22Kond3VicrvHyhOhqkf1vhldD4qNkgvLjPnVib5tbe3gtMctK9
xoNmj///yLvBZlV2UD6eRPqMnfr4kgEB3weQawwPDlMmQ6k4z0VosStdMLQSAGB4
ZDJFNf6J9V5/KuefX1Ua0LIS2WI9l/kBWLOvAlaolFqyAfw3k9wiMd/HjPpsB6BE
MEqYrXTqMI6g6wBizMxCBg+SrZ+KR3DBGMWk12fHoyxt/Cie7Pc2Wl/ITBhWjiQE
QYKi6KwH+szdbhRkT1IR0hn4BT2HjuJisKET+mEcD2VjnNGEnHbLzAD1W6mt3znl
Hqb0vO4ElalfRooCXzpOJ4Ooxnzs8xorKaZURWXFKcSEGaoY82x4yF7K8tdjdKMe
Y/0+bTzSZqHNNh5O0ls+dbn45ICC/mLQBeL27uU4cIAZWjnfp32tPlU+PDccmlz2
yToiiGgIfvt5lzi/7s/Fkilnenz6mztcE8qzRwj1AhVYW7ceLbWOIA1ZQo44/3M9
+PmvMykM5rJ6tcEnM1mo5027yu3W5krE3qgWHqznfFaWWtZNMbysFKrbtNQVOzsq
df/l6L9iPYHq2MBsYi2IgDA1ltSxbbWce03ruH4KhIoaDkjGf4RIZLnNq5bO6NvL
N5zQT61Ag9tItnxOK1yGXpE7xFNGyBhUCPz76nLAGiTEgWJ84S4VAj1Z04/6HZH+
2YO73lFOCen7++S1xF8+UyqGTwQi85zyghEyl2JXlJYJja6b8HXlagx0sh8lyuTt
ylNLPHmYvMl8y8IPkF6e6WXYagOKKczOhzsJZRbyTrb4PHQkNZmuXkmhbx2IGWte
/pB56QhWspyUBr7ur23t7ZDYfFdtkCh2dBtQB5UhOdbE1HdP56TvqdPORb+s3Pr9
tTPn4jmB9Jz8QBzZP2Ah4fyl4QbrjeQu/VKyQ5E9GFbGWTyMRBYQebWtFmCFpUTO
3LmRO3mxyMZEK5cBEA9Nvo7fba/E5J9/pZaxw61ZHzUzpS1oGK05Rfn4a/vxNG5Z
UL8LOhtXF3Utl7IDhQBS/p3iX+yRKyI2UvN7G28tGwxGLsBuVWp0vGEieTlo035h
k6MPq1oD7BxOcLnupljJEobQn6g2VzDObKfLCbpj0/GooisChs1o/QMEZZ9nq/jJ
4Wi0ssRsIxxZCE8WfLL7TdUQEnRXU8PrygggACAIcZgudZUQq6Z1MUzM7yQdFiRF
ATxoGWkt4FQjYH346Teq/qXnebwVSVaQ5rYAqoGCofeokOcDsura0H2HOIH48+5K
BmJhOLF9dUBv/5u5yBf56Wt394caWNkSEL8CvAv9X84Tmb19lpYXzidBK15+JmXY
5pnP1VdrpMXQbBcNB8A/rbu/F7qrtjBXiE0E8d7TrKx59E6VH84FijdOOO+XuaRo
HkPWMuS++4mFh1WKpewaXL/sCmphNKKnCSg0naYyx6tewdQokN2VixVvOqK8dmQe
QsH9kSW11cSiRmmQRbsp8Jm/GDwFmGsjE3tyY/wG+jgGwaOVbaMLMR7nYQDUGIr/
nGdNQ+E7XAAi0YEszG5ojn0g8zFYWie1pY+rW6UJbGBMxSAPtQiklJACkpe60g8k
IfR4BBb1bu4sFPQHl/LKsVsl+6l/JQ9VJD+nPjgDAA2zT42w7O8Q3YZTUIPdNVF7
BPtPIUiLcwoeqmsSK/eOG4r9dZAr4v1zgPxP973yE/8NJWc6gzL7JkqwHouJ4ryy
YZ1ipPKQbwIcwvRkKkHIl5PAsoUi/hIPO34AlvY1hta/JDsN5guSdz9S+BqyR5ZX
b9hj5JTzDm7+vbdTCI1s5LoKDzuBDCXR/QkAoFs8PRU842EW2UtT1k3Gp+vEXkmV
baCsJCYr8NzsWEb5r1/bNePDYuMdCjpNsQE30jG7Twr1Qj5IGDdBmKzN2fQUSGxq
gMbHVLE12Vcc8JOrS5TWkwxG8LeUCkKKkvWWyS4JC05N78cOy6qjY2GKn8aiXEye
gyLOjGM2yivW+33gVbt8xfgRkn3OsKSsQBj/yWXdHNaIT52p1DjWtAYXyQG5By0w
ZwbHVmQkUGL5g4TX1WLflMOXRuifrsek68HGw8ZIal5LMSBgG76/DGopWdYAY3WP
v6O40KgRBZROeUW+DT0NlB9xD9nZw0rsfum6DCZnB7nybIXzFF98Iuj7HgirzEY1
BqHIBheYHx+7Wnoi+3PkVBfHV9NAd9CDCcIwwUashmBA+A1vo6ZiBZMYbjAFrXXN
xp4egMIfB6k0yUSavvZoyudGHiY6EXJKsMsgCcCaZrL3sTwhhXXFz0v0yJ/e6PTo
6LiqAtwLVi3kvTZIBB4HQpTnPBSvQXuvaxXvBxskuuFntd877KcYeWOwyQDttddh
O+wEan40g8Ub1l+hFsAFruwetlSWPFQ9tFY8dwNXxqQt+EWVzM1gnsk4Y77txAS3
H7mI2ejoXqDbZPsnHdckmvTYoCKRJqTDasa5LEnLPKSYaEgkD7W6/V+f/L66tdI4
a9VS+o8MibXpvM3O7anbSaJhUT5phlSNMW7PUKt8CRXGn+v92SlG72dDr/4nEPdf
dtNH1iWz/lzFhUf7yGFGdtXlZHimg2DkKBH8eSixR/ZfYHzIsgAb8eyDHNJ7Gs2+
L8y3fw58EjGiq7RWgwlnWpYQJ32I4c6mGILhscpbzDakfMq3UKFiSyuRusaxIHWj
2bOvkWsWUcFT/D3bzw9WVbBLWbo9N3n4MqMxNRTPOqfYrxKOZWWuZkGvLNSAwpWg
yn5pwXo0xTEBM+6BHmwYUWGw0sbs61EIqImHxgkk48PXvj/rhifCdQ3uNLrLD1Od
YLXhfoTbRoR0Imprb0yHLo8n1PSgcme+eus7peatl3FMj+jW4XFI5ltU66ALYTOS
5TINxQMZAJ5oibBR+4ULFsMUbPsGYnNSMySPvz6bUJrUWNb93Hji+0UfuAUU8hqj
QS15Dar0Vr1Ppk1Kl9/qeJLcYVrycsYYBIwydAvAcyl4J+IsmUfb9a9RIM/0EqFf
4T8IG2eJGJtfVdoSfVU0AxPGN9vnWY5VX1cC2dcb4Hc1aJErPTVDzt0lc3ppZ3EN
4vVQM1lxs7XbpV9J3EpS4aOoXnR+HfVwswTXEwVANyD3SqrKOW2A4WPbRTBITgXj
0TutOsbwVMVgXnY4a4/fd56OtVoPhiFE+NzC7PmkuGubdF8GmPYszgiHEwOsEp0Y
okHWP0kizMQJRn+6O3U+lIPzuT0faCPnMMIo0F1if3LigoH3X/nidi9Br7t+Fq7x
cRrgKrTyBF7XPR1AJUWFLQWy1YJNgtm27JCL15MmtsOiFeADQNRUNe+spmYUse9S
ITFEWz7Zn6FJRAoJ5ANeIKxGL++isnu37HzbDEq+qoFOEFkHeir/ZGPeUK8C7Ds1
VMBHGNjTBkg0BkVkDsF3J+dYBrPhpQY9RGm1mi1129LJQTVNESuTZrXwQ0hfCgRS
RbYV5voZNn/kc8bwdUkm8lsc05v5uAkH1MbAQXWclykBHzx/Yo4S+rZujVSaXu8I
X5Dnvty1iaQW3U7DXwk/byBgAIjaq2EBuFtGWk5RrcxnUCr90/xLoedR39TJZ22/
wO+DBry++p20Xkp8xSthjD2oVRtH63SSuBe7S7FHiU8VJnQhKRDwjkhj24fVGOOM
gb2iDtawFjrwaGgfHHGVYXNyC3GYYMD2FDeFKKE0PNgIRwmKCA5t2CElGHZ/YU6p
bqKuO1XXJ7x+hZuY6EbPUhf8rAPgQ2z8DSzzlgV8C47EfIRYnWctUgRqTVzl9WoW
93ZjkX0UpH6VFiDP3QX2BsnLLJzRygtVq5Ju+vX3oMjezlWUK3mAvLd270EEXptl
LnvQmVuuy26bsyHhpbbLAHLo+YoDU7uV/zE/JAjU23rQL+nyRFS5BiEXOyQiQPzw
uMPwlrdOFiX08374SIr9Jr+HOiOov0p5/xAS87ZPMVKNK8TP+hmwaYigZ/KnrP2F
iJcDUQjorZc9yuEaLGJ7PlpiFOvsak1T226H4Xa6esbgLkcpr7k3CfyTjI7h7OeT
qvbCyaFVOlFizl/peP4imxowuLnLRhf7T0+bYUl0TUNno8Tr26mSy6Q7tcw+KsHv
/hWTEun0j6ldUXUgvckC3MSEGcQkMExKQIy8ViCTCeDJAPVA6qFlkbtAI7i/pf2+
aKalpHyd8yYTvalFH9O4/ZyNhDaj+uWafXUIJt+Pu9l9S60ywaOZzRPU2hhAiKep
m/8GEnK26e51Dh0fyq98RPHT922N3lIa0zi9ft4AJSZ/8SDP+0HK//GMBc/dm5Ms
2/lWSawlx/adX5WT+bvrLBn26t1ae8GoU7sonAu7gYojaxbk7A2Bs+sLchO6LQjg
wY0l1BLNWbbKbQlYpW7qHMWRKN2KIS6B9bLb/4Wp74//om3/Bb99RofLxyxeo+9Q
yicPtSTyzm8hKOR6R69/X3uIMSLv/5QCfeuVfYJKnPqenqb5XpVH6dc9TyhRc8VZ
f2kZXgSztdEdn2uVAGhKcTa7C7y5weBR2Ts02Kb2lYg+F7I4EpmlXngudGccTUHA
LDtSqrUK30m2PitWdlrQerxgDXoezjSn00yIN2wf9SQIcyWbHVTkI58AS7KSKGw6
Ca2CpkO4WF0W24D1vUzQBPZ+rzFqZ+kprzoLJWENghDsfjC7JusObtJgJeye/bfJ
kDmk8vmWpUGjMGa/wLt0+sW9X7mrUEc5eBvvmzNdWbXgKGUQlU3+VdBd4cvP4kJt
ve5A2Kd++JxQPMqL8NEjoF/JgJfFvsFnsj6EADKqWZZwFzJZUsJ24aIAopz+JC0W
bkhpUkoi6ox5LfBDcfiFLH9oPjYrSE87ixO9866ybUYL0otxoNGvCSyNA/+uIqrD
D8jCSwhG6QQE2Z64aMM0hfddLb7DEmctXJkl9gXaXNLLI+SxD72xiXVDLTUwWnGP
CQq25g7XS5TzmZrQYdydEVf2VsGpzl6Do/FhUnDGevW4aGH/5gx3XPjWKdstQi+T
f69q6dwvsRRljEDFCGpMkuim301mX8gjb3IAQJ8EymFHy0b36UuosFIL+aVv6Oln
u16alU9QjN/qMtpPO/cRJHLZfs07SSwfJLei8ooHYSwQimNAZRuK6ep2ECN6qdaQ
fp64SQjPqfND4qJpFqTk44oCt7moLCHTRzZDR52u+7um67W1kDmzwjUODaKkgfa9
scAXWHRTbp7dq4zUleuaABnLKS7unGLRgLKOKBbINW+89JK+qQG5F3eXL2KuNat1
B4lilDtUMf70AZqjl5+IhLyGjMAQbRMd6muSwRhPmxXuW4IxaRXVxInlr92IM3tc
SjvGn3N2T1vrZ6CJmvxVPSKKSujhVe3aUf189a+sIe8l8adGa/HFp7kPgCkpdRky
Xjhpk/eRdXKi9ORO6uD19UYplsZOPW02ZZY06xMrg9ob/qN7/awqj4i15wItsSpa
McA0oC+8Fk/4m+ej/U3FO0vjyDG24Z+BrZ8cRG/09ev3OxWCSzvK4XALcnQaDqDw
TKNDl0KqKS38HBGKFXz2u/R2vsDej1nkE6Ea8WjNNPzk1Cswk9A6WGCe0eYBc2O0
/yaommPKnOPcmmt1ig/w4jBU0AAln4C+yZkZRQ3YNcs0r920ouq0/C7oHsHSHtbT
BpL9TbMymEGpA/HXnss4F3Wz9609/pDIxnlhI+O+ZMdqYkgWROP//GnaZZh81/0L
O+PVfnZ5wxoCUyI1EXu6PxIZ1ppKFNUKfOW/mT3wAV/Lj5cHAaO93+vEhG/qiAdG
3X8uKp+/A+p4GH1cRxnvGBR/uZshvjzrLE++voUEjOCeq27bq7mWxv0uaxPGxO8w
jczwwPzGCg6BdH6DnC5kq8a8hoRH+NvK127F/k0hu9Za6PTA3ZUhGYR2Z+M3AkbZ
UJxO1VfhbZFjtoSONp0ftpFMByN7Xcq/0D1KcKk7EOlGd8FJz+GuNyHwsD5wyEsP
/Ceb6y8em1KoaOVBrJED6QjoRUFXHUPpZ3ZcRJ9gCzVfi0BxF9HDWw+gxsNEU9m7
s0h0UpLu9c+j/6miOizi6WO/w0GrB0PSETsJ2CNmdUkS0E+sB57rJEg1dLx5HkcP
lGqgtTwg35yFHNFgnL2wpUlgr6zHD3P4nYavCSGulKOXsssWgNMPcQdANBfVcxKR
0LsJkLDqJWCOtu0JS32P0GNuAfEyafkgQLqNHZxQSrEs9yOjLv/0IkkaY/WaIv8A
bREZAh3H9JQ8LIN0iOrkyIgvAL+fkd5Ys/0LVDdImm/++4FfKx9gnnHFBfHh7Xk/
+ufcsftHt4rwaaULoq9v08XQOikHlcP3EsSe/R3CrBO3PapxuVXr5YegT1X84WxI
z6gg15OmkE9yvoIbLXdU7TCsKR/kvhzN4ZAAAbi4AJNc+svnWacrwNunmY8OmjLQ
9gEfG2sKoEGciSeINiZz0iEFTsZM/HHf6vgjNeGw23/mVqNzaCsOtnQp4mqzp+Si
I1jt/tuzPFDuyyz+iAJnNPU3aM7/7HQwptJp0jnbThrhw+TRQSnqsHkI55aKzYSe
GGV8zTXqvZBENys4mBih+YpmbRSMluePtYcIKBU2xDwTV+jvNSm+6G166sKrFAI7
PSXuZAXWh4V1KBiZ/e8rL4CJGAvUqNGOr2CjvuznLdsHAxjLRhqCpxi+geXt9hLU
esMT7FqMJozXan5LcaI13Ow4Qtt+zuwsMd41rRMsLwe8ytGzPTBkoIyHokwpYomD
dOORegu6JrkbCvhmuBDflU44Qd8H8lMz+0uqpma5GaztMfZ3Xj0rMA6TWUEgzkDd
b7eqU9ZQyEQ5TpLyWsQ23UXOCnQNzvGysQOlK6vPFfLcv+oOM5QFFb/yvD4FDbSW
G0B8tcPV1Y0T4+krZdAQ1DaXBPSG0qJSvdjA0Qb49l6yAIcuOmlIjK3j6KFVishG
M33oIZXVYc0vLNcfhKuH9yANut793BGusibbig0wDIc/K0s3DKszP0fDVRSLEffX
IQ7ZpPwaxX/Jv5bDauBhVjVPVm3ObH+CwBWUUIYXkUpkdnRa7mNNynd48CcFYAqf
TGE7Q4cWb5oFfr6tirLOI6RiVsRKXVL05anW1hCQkKrM1ZjNSTRRg38dprBHcvk+
6jWH7riBSba/KzQveduORlGHVAj+2opmhHfpxFrpfZnxzKb+c2Wy1CftDhbAJcZL
AtiAf35Ul9ts2p3d9yfI0IchacUAvW3xK4utqliAU5wBhiRU3KynYNB3W4U3+GiZ
1WQ1iCzlDmDguziCdjEOwe8QnnzCusuhfe7a/0P2DAptQTZZ/8xJ0tvPcqh/VH9G
f2IQV3kBF9F7ArloZDMIv82BXuWQpU1fT8ajfm3jPVousp0/ohAWI3D1S+RTLyRo
HDr+imEPai0m+da/gBbOldF1sQy+oHOLjNP+9hjoT3hzDDZIgUR2egs9cR2/91eU
UeK4zriMkUFqpg0RYpu/7DuA+xjsZ85jKvVLPqAB683qhg0c+eq5jLpoNiF4vhbV
QD9PolsvAWgF5VC2FGLjsU6nXL/Vvh7of11iVh3v2vvCBumPMaum7voOk5s2FTJT
4iBF2KiIc/mxa6exYdw13tsT4lSi1p5X5WoRBVcpkWU827TOaauFi30wnyckXuXL
J5oWysTwQB0cpl9MG0LtmyCFkmUbRlIgpW4K4r84HLXp7Jqio+P564qOIuJ7vuqq
jtip5sMwJjmzxzAsdDox13TrHSlWcZBxJqJ8I/QbBCZRWbCkvq720TFsLbtaY7NZ
+8vMNOIu9WVqdPPgkcwgJhFuCqnRHLRt416hXlAVNJVBQwFAaVSxCI8V6wlpICdI
zYBHADKb2LN1V80EOOTouDxH2RR2sexErc/9ir0iWCbQPijZ0bPBo+ZlfcL213pU
j/mSYjxm5w91E0c1nC7ofAoddrKauo/hwhmfQzLrNGWI2MkBfrCyxwA2cknDLIvR
LTl8qni1vgoBMBCFvMI23XehUiaEp4eIU0Nb6bOpRScVmS51OjtCzW5YUyUSbOWN
2gUUR5k3pzHQG/V8hVPwbI4zMhaO2/soAEdW4ZKUQdiVKdqrOPNY4fX17BuirtLL
DnA+SSo/MGIv4vhAho8Kc1c35JxBLsSHOXo5qAZehD4=
`protect END_PROTECTED
