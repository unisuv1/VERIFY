`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2ksDCzzZxJFOwDU962PTTseFhJuXy87KKXZU8jpYFaLLVfChxUO8bEevjE4X2WHZ
ReHdD8KYhCgICPUvn13ML//Y1QczjA6a2E737oHU7HJIW/tvmsqG0GL5F7Vi+ex9
IAxuKA5bYQi10UzmFvbbeJ4JtlwCR4FK+J5xJX7zUy4ut7/dwK/3hKmMPYbDo0iN
VHfFUJsqxWB8tKxu45zD5n+GK9NZ/soxhvf20/iaO6RF+XhmI8b+Tl9KTzoCBuq+
44RzrWCgMYny9W1QGTOWfkODjDq/EWuFyQBKjgK3kClUW5fiI821MIO+x35qxiWW
dkhZeubcP04exO7OHPeea4IdetaiU+6f+7C0oFA3+DRHqC8xT2OG4Q9qzaXyEZFd
B6kcqVZ68NcP695vqXOfgpD3RAmH05SqWH15LVKt5OBfGRA78QkAQtG1Ix5TDN5q
L0Cf2OwXQfalcb/Iii8SobW1KmXmIOFFDdKJOzTUqZEQTG0gX3qnY8JYjcMP5sSh
oC3aWKnFc/xkbuTdWYLHiMSWSv8oiHaxh0D90IkmwU45Us+Ks69RBS03rlcIiwDo
4TuzbRp30KdzxUkfpFb5C1A709d+BvrFge+eaLYq3NXXK6K+H9CtYEB6c8boiCHx
FhyTzfjXmgmZcUq2EGUiGRchwFBt+819APXFtO4TdMJDsZBMueHC90CBlLAStiy/
OU+lcobURMnVaGH/HlrrZMNUc4WOMeYjCgOjQO0ekMkqYq1VHuwvXtmiAZp8+7T0
xnaOWna3KeSzWQPHttx41zlkdIVaJsT9Woz0q0+H17kanwKVVj5VWI21nV5K/tFk
ClqWuDH2bPe89JcfFsCd3EPzTfkvcrAFEdJ1iG5EOdwAuXDL8UqRglFBr3VHT1PB
Y6vgQkawraP5b8jQzlStsizdXiGIF4hAbwvsWbRyRnzjzxcPIYEtSLcHautyIvH3
uw3uHKBabgTA27CqkxSGEwUZW+H/ASItSGoyLvQAefH2+cMpVNm0SSNr2QHMYUxt
KM3xVtpZpW1VU8eG164wR2ckBRR7WpuIEjmlcvKsWOiRyE3T0YhRaOtirPKcq/JQ
e9jK8nAAdbTnaPMV3GSati49R3La+XNiYrb6umUWeVQXYEUBZQau5+nLFIhvHN2e
svWFuK+oCldUrzjOfFxhriIQl+lWf0eLUaUGf4F/+tUU3BXP59Wfl4Fwl7vJ8hrF
rcFw5QxVAQD8dG34usLUdAA/1NXLsutxXlnb0z1o14uRLGBxamu88zwLBIs8/Wc5
Yr4UQsfZG9WdBx6jFIVhLG/nDDMWJ/aWsdM3+c+GHOi1zLP7OuusMP+9hj02y+AH
IR975T1ihNv0Jn3Oxk/jpGfcM0+12nswCXZmPKZBO2SWbwrf4Nypt0V+0s+ikr8p
IkUfDSR53ThCPcMcwpzkqwfulsIN1FVxxHZwegeWLmipNoVQXVu5SfjwGtu5LTso
TX74L17JxqirYleY6SUq7RiEn48igv8XyDvzRSsB4VHeHXhAUWxcOI9Ia9EO1osF
wfVYotG14mxSqFaaT+ecEzuZniVrAKB74xzx/8TT2qI7UseYFJAJ4HqYHcKbpGj0
iIiYuEEdN4t/HgNdZixBDmwfH/jWrgfUVowVFpJvE+FZkHJ2b830cAvU1n9nlRnB
MNGFuzWAwp8sz0mL73cwLoQ1sYu2pok1FwuRsVCtpz3gvwqLlntkpNleH1iWgQhv
6LX9l1rIM4DmrxytkqLa9M8TdC5DupZJiwmtFo8FT8uIynmn0ioKTRrWHpdL+ulq
LKl2KAzxW6Nqq4WStlAgsxo3bJOZgTwOjdCUWluQdb+kj8nGJZFSsjMGaDdVhTW6
wmuvJwZncpIQrZ2Cl8UtoGNPysP11SeN5xG9hEMQEp0J1Xd54HYQ389sxYLsln3A
VlW9iLUyGy70C4+zruAtcmhJAe4gs2P3Y91PlvUUUl6wSILcZmHq8BDYkHfbJ4AT
/4rRH7eQ8wusC3yHxvJcBqKBvHcfLyZ/XRvvLXyCRlPf+2eSoiEXocCSz+uXYA8b
pHOt6oeYiF5h1wvxF62WFGBM7BNeeQUPrjvFz+dnLM0Toc/Xv0JYqpxDGwhvElWs
dXKVRU5oOHfdgtlmctnK7OoQ8njp9BAbJgMj8Dlzlxp5VYMdRCqYRf0NzA09fMJW
LYCNjUOTlbe5PjmtOknSZbLsudyoq3l3dEK+uNRg5BY5BvrsyM1THdibp0WvxmuU
7ZFifVDMjIivjCIfSz9a3boJ36HxG6j+A2ukZ8HQAxZMxCU48SMNeFE3pTuTfdOy
mBHLsm2AViaQTQVwroBxs4Lvpz+622f07SPBkU1kPu8g3jFRC45MuM9Op+YAXYlN
tcGJNH5O5XxeS0Go5LBiyn2r5+ulpwnfyByODN0z7TGkYmG5yiTGdGfolZI27FVj
8PvAz0Jm6hPDS5yrsJ1bfUO/P4bMwWDYpoJQ251R5yd+AeSpN5jA7Q77Om8GHlj1
NYY+H58WNc6q6gVR6HQ7wN93Q3NZ79L9JL0B5BtQ2ccXCwzM4ODhpnaZnZcbUQWb
cp0p8Kwlht5cinYVzTOKrPTZVQwD+ut1APZ+me4x0cbQ8nTKb/4ciwfPR8Yvbh4k
0fb4TypHVHIkv/5ImqFXQOPh//PsuNs0bO0D/QAOFmCb8GKS2Pkc1/SH84pFPk3b
vf17Wxz8h/xclk/SUWcpixIj/py81RpJvvmoAGaOADuvpXPph4dJF4/9AYVJtD8n
P3WkGskwBbKTfnL7c2AP+g4smp5+h6ff0x9B1z5lfcDkHouQztsqp2pabg62Z4nn
XSPwIAQwJE2823b5qRxb41hpnTtqpxw8tCKScX671kuvkR4ouVye5EqZbohfFys9
59nBVlH1xP3tO5KKz/lQ6z53AV6Oa2Wk19+pvTBE8NX9317qe+9QBQK1B3WA0gwl
8lqRsA9vOqBK+gTnXNaOZGMdDAdmvk/PJxQzur4PMAiRZ8n1zRHjdzV4/SS4nlvB
1e5wUL7HNHEC2cQ6OyGl97Kw83YlCxHRwHrLmBE/pDG44m/GDJwAItLIy0TqeRmM
vvKEWVg+ZyNTJ4nSnaEijVvJ9ufZ8Oouz+xaM69P/zH+Cxrz8eINOVjdy+YTxU0D
S55wjdtfabL0lk/OFy/9SU9eqS/hVFeTHzGhEIL5F8AnqpOxahCDgb+QEfbKdFkI
jQ3DrVn8b+HyYlvKfyil9autOby3lM8THxLax2jG3k35dlIJ1APGAX+CITePCvyS
qlbbIO4E7WaM/ts0p1oRV+iXCutfZXhQycrOSqKtSyg9fsWau4AVAHBbaPEWzFAo
zxLxxMhak4I/V8S/eLCOYMNJGKWNYOrq3oYRohTqTdsRtjYILLI9/CnGggTpLx80
2w8p4l9sPDPHFAuluV5kxV8p81enWjsnM021rL5eqg+WPamMidUi1aKfo85ht2HN
Eck35MuD1ubGrJlMZsPNqMJsAqeX2e3B0zKCxWEtlm83dT5gzaYV4FeX9a8TtRZI
xYJkFak6CzMzT++9WghAB5KHd7xUO4rX5mQKYClr2cLkYvgFaAy5xFAXDEsG4MgB
IECZcYcAwGk8u6O39e8ck1S/DIGzlZErjrH02/m+X6FH9ZrNvzL9KIpPKepooBVI
xfZdcyGYmBT6Ggq9nyxLdCcZ8ZyBFHc3iLty0UY7F+XDQiZ09SCw5dugmJvGlwFB
qC1vOMeywi98YJnkYzRw0g==
`protect END_PROTECTED
