`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D8FZo4cQBHX9TmGzV5i2QImqbxYcdluSK4R1ahYF8XravVc9AKLjJ22qkl17hO1K
3awp9iWfGEOY7ac/gd1Ze4HFWWVJQPen4HBT0xyQHmH/XOWKptoQ17zVI9OvjEXU
gJTkqhDLn6nxU5VA9PNHrHKmkKKRn+mo2ip/Py90cxO8rRYbzHNcYcQ1fYW7K6cE
kk9VP/qGkflXIMJ51t1D+JqoS8jPgkJHkNb5XxtbHGg0IQyE0SYacyggFzi0VO/6
IRWsua0QAlovnMI5m/V73uBG0YtkIoBd1ALVwvGkMytgJ0mYMdNNg4/AaqvCTeg/
suhNxSVi/UNL+TB8sZjK7dd+K85NpFYwb8vVJ+j/LPtJGvTHIOE1dQQ60dKnhYZb
59HyjmHO7exeMy/hbNKsmY5ed6QYiatjw+8dZ4NvZW3LvY/97JHaGJvGKuajuFZs
Xk5r1zscCNYuXt6EhxBxjlwsK3JrtuJQkq1dsSA+50WBtYfcFQyLREcvzqGLbmkO
n5/oOBcsBfm+3COzilM1v4y9rl5iDd4O95e93bSwpMPIDulYknz/rYDdpgokSWQB
EYqpgckCoDonybCuCf8ZH7Jj7Ra3V0/HEg4hNGSQxIkTNXklJkE9eJUbTEmOxOaC
I5AGJg+0LYGD/SvsC/q1wKjIzGfgIcHzlj5wihl0lFsvqBAS2MFoUgaHSpL8ftb1
BWWfwJ3kQ8Lu5ozwraPYG80D5QNStT92ISvZyn+4KGafjOt+0gEMxd0K3Yb+M3dw
rd3TakLLtMnh/FqO24mXoJSgAJyWi8Q+vNZSs7eoUg0A3quNHtArChynrfIJbhsJ
bOKsPWmhg3qUkzOWgP2MMIvmCd6Wh+R+tGiIeyZ2VmRBb5z7p591W8jkxM5mU6aW
lP59PAXYR4F4RHKVwo031k8HEoyYInJOtaC36NvwmmA4TsIdNTT9+NpfcKPDvih1
iLm9Ur3oIU3InikosU2xAWPO3H3887PbXA8H5G/8yCW5NZx5mCWG5s6bOFCuNfeU
tJeA+YUp0eEtPGvhP3s542gtlge+ErvZ3f61fVolJZT6lp4OcAwdiTSwXrqLldDO
bCLBBMATBG//D+MwezFZu3d8k2kUVPHF/VNlSy5rGDy7kurml/m602EAJlyY7JaT
AemQOnOK3+I5p/eTq/j20gEv0SBmmjAl9H2G1AfSMTsMk9SLRj5/chhuSXAJDavc
TstXUJGBTRcT7aOpECKdQw86ORwDj8ZD5gWTeLtMxDi4nSsYwkSJVaE2oqbYtYCo
VA/Xprk8s9aekt4/TGkk4lzqocjEQLTbQUtQc7KNub0xXYvyVscCKmZrsyc5Wy4n
lB6HG+NtUBwOZdV5uBEh9A9Uo1YxHaggBVvvZcTICCXVjJXyxgnC7lIWPicvYvXR
9qzNP7T8Gj/u4Jl57GFAtGZRYImDP1hzM+0FxYedXwW27GNK5qntU3iMAxa86AHn
9JDNjdA67TxCVG9nTkDrwv0gTbGl9UNdMCPEVHsdLA3Ab1HHhoD8cGW8EYOHbyNr
Xent/VXCsXglAMXKNmudi/A9FbZmiiEDCn8PY7ZAPfZv9YS4lxXyvrqHmWYIjz1I
IRX2dQhJipv6tbD+CgE5ewlXxIEcwuLEpHSMH4U2KfOVqZ9BRWd3E2tPeZ45YPbF
t7nda2YuPMyfZCoM2/xZv/EIHYGFawcYSAbCE/GEqC89q75sFp/zP7jinIfYy6Vl
gawZgmWDJojQh5XuXSjf3JTFViMwuH/nHe/8kllsnb7NaxeYeMAju77A9egpMyxQ
hjFsxbU0r2chui3zbXeZEVy+83lUWmhTY8sAUsVxfT1WVuc6aMD9+Y1UCTiheMNI
Tj4otfHGdVGiJTRJaEK5VlLc52Uw+Q2/BhHPDL7Amap6Fxkg+EQqzYoRSMWVwy34
kkyYyMJSn+FNaVqA6A18P087Ai9PBTum/x34DWmzumg7BJJuBC09HdRPd7bf6xdk
PcMD5F//Aov+CLbCktuIjW5fmenG17p/tUrhb4278W1HTmSkqezdorWoPWUuXfNT
TWmqyNgYSvCaYEtqrfnVhY2LiMLRrAej59THNSYSA94h2yNJ6aVzyFMRyArZv1jY
tzTroHUwUbyZ9DhnBXZOuzDKJz5Zgis+j+4ABuVTblQlR2aAfLPnziCFY4Vi5qEv
gnIG0/WKf/SQLWDaQe+3zZLkE2x99DrDfldS5yaqp/1SIPAIZq+/6OSlRzF0VJUW
uu5C2UmmwnkjSqIxMeob1/hurah32NUxoPyKP36GBcYtvboAsCwUejglRNAHCyrX
rvh/Qu4C5RK9Wwhogr9eo7h4NH9QmXXxS2kEeVhntJpcycDJ1yAocf2mAUAiPe//
h+IF3nWzIjwwL6g02/rwd77pCtyqNTbbwmXYtOPHg2D3rLL67eFSK9bTNqQWfaz7
HCBEzM/iGq/acEuLWHs7wx9dkVH4iq33K/O95tZ2Ra43tgY7tW+JTfugNn41ZoJ1
8YRaRVJMjbKP3JZxSeDMiF+9EojtZLQkVk43PtNmkSV8eBh9JPs3GktRwKAa7pa9
OKKdR3cf5A32NLzcZZJbPjvvgRl02rpBKPvQ69bh+8I2AwswVOWhbmbAZQBzRwrl
zK36AlLcLHJmivhETwAAgpV2lip8bPgwZRaGNwDZVT3HUise2M+LTcDgfyRVvl5q
wh696S1GWzpEf+2DOvjjdN9XP5ynnCPuAp36pnPTn9l3QQzXTDxP+cbzEdnJWrqY
zmnV4VUv2o1ROtRqgIl/okPsOVJAKGlJgIhIJ476B5aGcFa43DuldYSqd4Ltbd+l
yTDHGWLpiHUl7QyUkJFr38TDzkesYnEQEMDAXDgaL/cpWm9yWNWC6Sq2pivqiMf3
/YN2vzlXoGPRndXaNtXir9WO2vxPkqgOZYLyazjFL0mERSO38aKyh4GalKVZA08v
EkUU3EOqls6PJlQhreXmXI6VCxG+KlPAfvGdY2XJfX+qJTzyqGve8TIU3trrfLf5
ts+AH72E7Ix7P+bJNGOFUrn5M1ETLHX/ece8WHiNRIU22271EpaejnVpNeKt71Wv
ocwwGnCcm7qJCL7HP+O7M9ZzQbrrdyx0WG9sXVAJyCl+D3Ry8nkWyfMJOAeii9Di
9wtSIDFHcLO1508cETPamVILpLB2M1QloSsVMZcNERw75S+HBfb0IumzklZvtnOW
GgmwdfeFVFV8STOFltPqlZnOM7c6NGXIGlrlINP+A5853OTTJpdeXjciTG1fRvdI
vnxOONGWPFtpNT6iXPEdZLPr98Ndgd6PWRwY/jxR90LO1/6XMnsf1gjPRULbPKwt
IC4tsXv9VljeUKUa0Hxb0IcBYwknVzYNXdc38KbYQRqP6H5NMAcFpswp9k3x4NBh
gH0fDvs6KbIGlozhZbQ8rKC0BnDJiSlG7WPj01JTxkQjn7V6JAH+e4yrNXkwIjph
iknskgqDyCyCZgUx1LobmEYeToIZH/+72XN2znERE7xaiF6W+xuQWNHjZW/y1KmL
TmHMvX7FgVsB4gtgw/10ZzqFqYmZMP5QF2M8zx+xcnAYwFBNoSr5d0J6PJytsTTB
XMkkpKm3LlxU3TxpzcLa7srgyHQxe4tB422EbF5PtpejhEDCTR8/7rdGOioTMeil
dsHHWr2iMleOXwcJsIkvFZG0UGRDTzBs3EOPvpkHNh6li970QTHsiXiGXPq1Wk+G
qLpCNlWLA2zWuxO+unxJIssHU8UgGy6ncAtsMuuF28hxRqwcEj0ZIc/UjZ3Sl2Ai
cwu0r9m66A61VdTHVy32aq6nTeCXmTDAPyPtFn1/iQPcCxg9cGUd+2BKlawsSxgG
BdekldmCX9xoUxkUO42RHZQt2g49K1/xJBzy4p9+q4Bh1XZKJTDi4zYmlibkwL2Y
WIK5quK0rpMpNxuQ/imWyxILDkrFPZ3JAIE3dOxO2Haus72YugUSLVoJd8TnWjxU
HUiCvOI0tB5VfJv/YjKS6fYna0X+9rncuHOSGiRXAxmN64yDisMSG0IQw2JkyA7P
5SbVBSHxiEfSoIsMuRVq8XY2r4T1zWwGJR0yjrtZBftAimx4fZxaxT3et2Efd1H8
kz6eqGXBqp4nwPcfM6fg7YIM3bQAOEU/y7JF7UyTm0FhUma+xqprZ+EA5TI9JNaQ
ONUJabcJTFMOYpu1HRkIcyZJxKRXDXPPjOKnT17M3xcVlsungYb4z3xBtUNyoAjw
G/73ak+UPdC/TZD3i6BZwG8KB3t36Tl04rTWMi1khQmDhx2xAM5UOikK/xb0MF4h
zbfbe6Zq354gtkrLDfy8A7HYovbSaA+TzOAqwFbzKYByT6ssY7aSTEvXYpiop828
FjhFLAPbEYFNhxcTAzrOQbRK7Cb9iKHDBBhX9DcERqbzNB5NnskQRCv98zdsVlcK
Us7eQho0OZR6MwzB4+uHywdgwZOsSDyvzxLbs4qDhb9UkQUHkmXG0f/UihSfwnOV
yGT4NEV7fw7DZxTivXNdar2QfG1irE/jAaJEHUYckmy+K6vGOvFathE/GTiDmTQ2
1S3hTrSyz4qiqpY3hI9OEzNz85DoRbEaVg/4hbJfNSipVALeEBIUPZYO0V5707i+
7xkdypCOl8/B8ftpIyuZrx+fU/XQn6mkWxxKXXumP+P3JgHj+b1iJ/3E3or+gGDS
hWrA/YutG38k7VToJQEcU/ttc6vsIfCUZisfRb6YfeZOcayHsZJqGNXnoBDLLsWp
jolNqUyOJ7SeCXqUjsgZF3TL+HX77XS9+DHYz2VQjOyX/xcX0v8Wm4Sos+D8LVZO
QvQbVvx7HWuaPNyNuKpSSn2hDmAG6dGFayHTxbjXNE2vpZiivuuQlIw83WLZ/R8E
I3CvB+XWa3R39IcB8V7B7rXB8/5vCJaazZtvSIA5dwh2/6ApiUB4Gwj84vaEzmfV
eWx4wgVPFQwJcaHmxKOu3xyaF80LRA0fA1Gsr+QbK9ODo7xuNd4IS1kM4kbEy2D6
aBsCliDbU5Ey2BRiyKr7Y/a52Rza2mISi2Pr8n+P05nAiJ3y4Id98OG6Z7y0Voa9
6OwApqww9Offh4fQWNg+yBsfZOm2smtVlyNYRCBdY9OpEKEXLpBiMgXYHoI+bWEg
1vQvBs1YkqSufTQqZuA2Q9Cw2Gn9HIxwjOHuWqUYFlcsDvWaaY1caIlL6CoujsH0
28m5DisLqvIAhC4jfAiRyFvME+PECwHLCDpYHU+ktJyeMp48fwQhGd42OXWH0yvR
j20LSfbq1HGmXE7dvDZzP6gHCUxk1GyTVzh1YZy1GjXSVWzkqJ2wUHe1dbgt9JoE
xjAhVuA3TBPboJqqEVr+C+jItt8QFh0yeqpQdx3CQRGn4GIZ04EDDc/6XvD4tR1O
dSmS3qnazYLNb4DY7S964KnTk6tTxn1mW5iy3frtYq2toEAKI/my1fIG7XMwjLm5
G86t5yvglhE+lAFkd3APDAs0cTgKvQkEyExM+QxAnKdUm1wpUXHANY+zu+uJ4VT9
jyjtb/OKvaTQEsM8isoY9eviO7nX7Prnqs9CaQHY83f/ogIKNU8GPGweamAA9h2N
Ob3wVViyYRN4Wx0qhWgs4avCxfD7b8a0ilWSWdRaJcD1Bhdx632DFtKvjUP9qy8J
6p7d0uO5ghBGH6iqP6c5wozhI6pmtB/RGKY1iyA2kBTrG1JVKbtbLB2yjqA6QwRY
O/8/fgrx/jnYbk0OExjEo7lh79ximGIpPIsaTWtMsWKGpzr3JJmiJo2zSZC8H+Ex
vH7jkQl4lqq1DBBd7eC2bEFf1Ew6YyTFcHkueWXy2L5Lfmj9bZ7dM+SIUL4ec1Kx
c+EPs6R1uQl5BGxnA07e+9R25zSXZZi3YCmJ5k9c4W6To5MRr/uoDXHyPQlP8+ee
vj/DasIYcnWDn5WDGbTtln9evb6MWA5ums8yb7GWMu9SClmd0LGsmz/ZlKZLD/3/
y/07IcH9P6MuW4oUKIC2W/Ubr3kXD9TPf56t0wAM3G2McGhW4bffCeAUg1uv3BJ6
0YhKaoVLB9fqbM8IhYUNgvgoC0I+PZwJSzvaE5QcUnCxfudALrHVwMsNXubfV0GG
yysr6ECd2BG4+f0LdVXTt1n11RLuCMd3EaIw96mZ+1+4D03LhfKlBrITkG+AHN/s
E6w9WYMADH4zFkmcC/QNMABrfQKideD+qB0ht9tEKX5bHSkx1dA2BH31v0mSmg/z
fFlGcMoaXiiMRxxeTPMwfiw/2xIANP9PZGkSYLQQiZ0OFfTVm9/huDQgfDg3Mm5e
TmE+7GARRPJLd/0a+PnFRCFqzvyuagzZj5/xsdi6olQXwdK4QFq/LJoKhikk1wJh
7xHNiP2vKtTsBU9yYts4REKo7oYRESu49MqEYW7WJY0qeNjgDN3V0aJGpY9flF1o
StivPCvF3DNNHDIJMsPxK/aVG0binVDHCMMCOM8gAtd13jOXsFccSzDdNFGqaueL
tlCguhFuXvmn9Y8AJugrB4KJSG4vKFn9eKf8EYzW6In0xlYxMm++NCpQ6HTXecng
E28HNx68Axe+h6rhqBdO6RztUI6wmZ03g/PISX1a6K7OwfEtX1+1eWf13lpLJBeh
ML2QEOUrnkkZNSRwKWFybc0/iFNc7n/Yf2v8NXfFRer8HTSleuEfqrVIL2LQCEyr
gcy0iWYLjZN5+4EH8Ck9QhTCpuZ79e0YaoeQQM0FblOPpgY/wpobopv6/tbeBurE
zg2LxZ0OZnfh3ywCJeebc4mfIIdlYVyo5Q0TrXy0j5hdpbuHRbJd2wo8DUesmLyK
SJq9JAaTj7W3LHeQ0i9r8YRbBZgrle8OoeTH3/AM4IYXLE7jdp3wmuUuPZx0dlF/
qXxAOj5x/yTMuvpJ2jpp3MHY+Eu7oTv4XaMXCiP67Q7wkXyknOdwSufi1ge8FApl
10zR7oVBvU0UubgjShPRdUbx61+cZ1muxI/gH38U+y/4OVXRsTQz6DjsSeB/QPRC
gj9l9Op6MtIpoJtz5/9QyqVd3AMWWBoZfwF9aYNeqJJfoYAorsHMljSg9QPUFWTK
IifVbz0wZ3wC2/l89bN/74esAfMcXngoi+TxnVEXkzwbOQIvjf9X4oKuSheV1kcu
YBja5nyxoaVqvGZz/Toi1zaBzimGRu78eHRdIRVndloW+2/oUyA9linOaQS3uQI/
aD/OSH8ZCxmG3iZ/MEXHSQA5uLgs6FJfYu6Jdi2jybU+zg++HeGKVbseNmpipNLw
DSsVUhMEe4N4BXBkC+fzAGpRqRNQYGJTHFXDkh9gLEb8ObAy82PeilNDbRkvQC7m
MPEiqklGvTCsgBTV5hMqnLJ3ZOW86RbhB79y7V/2ZzJeKpo0OH0daD061nzup/Yf
Qn9AerBMMvv4+YiFhykM3UFXsx0VflR7NX98OYLefQie4QyVJITTse14xEAVoAnP
Rtyy8CSTBkdvRXzS45GSdIXzGPgAvyGFrTrF9BPskTfJjcUwi6S4O1pb0WYMHgYY
fSXpLXYHrhL9o+gA2lWiCLjnZnnbZGc3mDI2S8TOTRQOHwxCLVZ2Q4gXq/yLsVMj
Iia0Um5cv/CFhoP4zUhyVKEL1GhGwt7Zx9kApatyi/VBSpA/JT7gad5V/gxww/gl
iv9/jVkYjJEn9vhPEFSXZ/H56uvNoa/gI4N7VVFselr3D9Z827R/cAULIYlB0Xpl
I5DMwhiu5jbyK/ALS8UxFd27vUtgzF/aFtCld/k+nox0e7jBVslVUfPyyI8WAEqO
Xog8SDdVMjttcTxt5eHOxoUhR1MHeVldL7O+VvpKcOheeFDETeWAgBohZca3RPNx
d5qYQAt3wTL4O6V6THQTjM2XuviB/NtQh3N2l0X6VhoVtjTc/bUgiIsC+8F/E7lY
uiq7kuapngXElA0znDUJCi6s+V2y2MJMYTeUgXDxhdJ5FEmOQMXajz3bBlechZyG
uG3FIXiOgaDKCgg0Wc/FcUVT3XoKOfsLdTnDqgWsQRCuP0SU9bFTlNWLPDwezmY4
tLfXAHntgfULnCHFDw2t6MlR6KSBgJNA9CDRiTvJMecTc0qa9mO4BRZ9dPmfneDH
TcCwQk74ZUNJyenHHxllPx8YscOrXJiti9gJKD8Wu5IHF20F+VjnYrLc6uNAPvRo
u0vm91h9JQH17ke1h/2Q1O5Oz0PMwT0PZthHLA3JWUiq/aXZIAkAJqDoSsnvZ3HY
pnmgmr3Yl/aUuXJ4w25gKbbbYQ3PYHN154q3XO3lX8LnS+AeiWCJkq/In/pcjVj6
1+9h5q2pZeUnssATWnuCx0uRiegqIIdpifCKWRYqCf0d94HZm9o3aAZtZH2e1gcO
v1FOfO9T4k9uDjqFTANhM9aMcl3tMLIDrTbhUonnUzZoyt/lckmaA/mYMh8JEQEy
8yi81w2dlE6kIoJx3RMZgi8Xq+IG6Pv9RmmMrmzb5K3ome418OTGShtvTEYfKizp
gOBaw2ysWvG6FRd5KPrkx/40kOpE3ytD0MEDxs4BhuxWRuxW/yR4vPRsCaJnp4Ky
zieFZCbqnqjEQjSn0Tv/nPxyD/2sYr3kFgqvnnsAc3ktobsz4S8B9Erp/2t1Ew4P
89/hz+CuNl0Ksd4laqtPcNrAo8j/Oz1LfsduA6OgzthTJVsRpjs1mP++qQ/OFYK0
58cUGdXcU4cVX3wVcCsGEUngqjI5SfE2op0Rk3uyyCfX56ZdM+GUKzHjetuMjJwX
UrNVGhljytsEhDHbG08PCsQnTqMUDcKOA+kQmWe1c4e1dwhVTjsMLeaGd2ehzWHL
dVb/ReiewNSsgZbDsoYDLVmvyEI1Ma9VkEP2i1TtVEd4vCCgEYkHhSp3UchxxBIh
KAP8m1a68fBMoxQcBG9t/aoFYgPfdn1scZEnqDnSaZL9ClN3f7D7QmhdgQx2vCTD
irZCuuB403cZMwYzzU/6PgsxJVOc9VCqJQAtTwGPf8ScQ1sY4OB9Q8pQiFI5T/MH
+iFwQktXbs+/z4PSc0Yf1WA2caAPY+zbuI4XnHfX0N7540nEeTUp9R0mfIXvF2Kn
u57J/v7WcbssUai43IEyacEUkCqUCiq4QYzE2QnN3/x4J+GLjmhgT74AC5qaegaO
RHr2cZh5wF+ID901KYT2cy8cd+OHHoY1ZEusMoAkOFMgIrh/PmZA8ugwrrbmJ/lr
pLWJxFQcud4kG0iWqo6LfZNDzhO1FnHNIwAr+aS3aiVGRq/lQW8nAEQEeNC51Ox2
Lu6XNASotARTTiaO7T2eKRyREGzjW1gjnDota+xxJ4487vgz2nDqETrnE5x53LSe
dSt/Epe4Lo0i8IuqhiHDGU/smX2pw1Ng5bPXZTfr5R3GrtXAKUtI/2EBRan0/ECl
SBUrsVT5I2LDdxRvwcVV1koA+/Ryw8XSSes4z/w+DX+SU5l+vOTA5WwxTvp+9Dtm
+G9b/PFPsjn77nHZrIjYwhJk2l/2r6VJSJXF5uFOGuBzeaV+5j9G3eTgSJq8CeP9
0DYVP7/RMXuBCFcvtleBGaMyz93QLWSREGP/axNUWsO9Ua4Nd9NA5V+5JFP/yJsr
NqjYX4nZE9axFfpkln7fUYEr9e9Q64srGhedt76I19d7AQ9Cp8BfDRu4zYMrRyth
DAQyQyGgOdik9F6wmAoR2wWdqzmUVIapMERDOQoomoRneHHQzNRumTV8e7IHbGRm
m/IV+Xbtl8wmcOSSSHBO6ee2bypya+/N2f00FbZDpa2LLo4UrN+O0Ggju7ZUZric
91gmvFrptFK7nVt2mhyW2Dik2UxhYW0XqkqjPApGuKYCQw8HzNYUDQtCMT5tpo1l
6XekbS6hITh10msGq5yIvI0IMG8gqgUjrjekiMagQ0rfkwhSWCalyEjkZz3sin9s
yJPRMWitGD1aCGs4feT0pMmRh3YJrbVVgyAV/78WJwwGj+JX4AYQI70nfBaPp7a1
Ej4/ITSoOPcsWwxAJLljgYjSDcQSDXCMizwjDmZkNTF/hX3LiUqi8o9n1EEO9/0x
X02q1YD7XaMt40D4gmVoiSGlTQPufSmoSlLpHUS3D3iPDFcQiMfRC7B2SwMaiTD9
DH7m40vCtyFYNbquJM3/Xt73z88OdLkZHokGoEvPWqns3O0KGr+apWpstjbTj1sv
DIieWBU/GfPmeNfMKxc/kuUPfyqKI3ubQs3Il8eO/NkOGdaQ/rlNG6tQcxiIzv0s
7rK3R3ukDTRhy0xPCf9Xq96MoN310Ov+uw4DCDWcMuSgRNIfpxCDxTQP76OLVI0L
JFO3FkLBgIa/OaSsTtpMqnvYrnhYsxKccJYudzif42ahoJkmZDLmcK7RuFn8L8G8
xfqCojgqh+td2qcrIZ64IUgpLQ+tUfqBMMYSnqD3N3Sj8J9k0W64QTT9+jSyNHvo
L0spXnKHoE1P8jZliZJ+r3avMOKiu9vLpecw/BdfAm6SN8vDLYYefctX3KPlFMG8
Hn0K7hMAgFMl6bryUVaf4npZ3/tOCWwb7KlRP8pf6+74hlO2qowRDDodF+FHlGNJ
CzIPdSmeAivD144Uh2p/HzFM1K39X4HZ7/Yr1H4fPHWvs9cxIdbSmW36wPw4bwG/
ownsF4hzEeqp0mIawBLPykMGf14GMo3KzJ/zr6mKKK6aF0z+WSguc+HkPNzoFVdy
5sRxNXcWrIvrM0iY1Dr3dEOtdeLWJvoFc2m7mHu9tn1hPHG0VB3z285NzRbo0Pze
E2qzHk3kA7lF/8C/NnCWiL6NkUwQDOyV48M21F06fZi1Pq7pCC1asH1yim9NmdAw
q5neOZeMtAaTA8BRulzzxSW7qRxj7WQl/vYzMKRAMNWOBWxJfoy/I/w0rmA0Q+Z1
Pk0zKEws20QMPR1wv8vuYx+UthyS+JRNSVKz63iC+0TzE5pwTphhmdexFWgraYcJ
dFiUnZOdzw/uCAWgJsIRH1b2I9I2LcUkmR5Uh9VVSdOuJASsevk8vAtfZjZWYsDT
R1HXiQqTGVCl39U8Fx7WXbT0DNJL0TcgaqlCPEhgpTX2J/JjG9BksgkOs3vR177p
Dw2YiessEdUdpF6Pqo0ExCj7WYfPce3zRyPp/Y3O68cEuRwgNBlhJS0ByFyGIlrY
rVoVqpADUECWsuH7L+c64n5FzJrN8X2mn6DZbnpVoi9kRvS6FvegGZ7e3sbbrSe2
UaOlroVWaOSw7NwZifqxJ9cNDDpprlDQDFK+WptTzd9vjou6gJlqbFj9eqhV4gj/
dLTsm7mkWNDV13TsbKdb8440AskX1WEzy6KtK8cwUt1YD1hmOHll0Vy386GaUecV
W08oj1POlkil5g9pRxtpS2Qm5rEnOWreKNscVp7r7JWXxxE29Wt1vk9Y1pkxPIiC
9tAq19gZQc2ssaUMkKNUTfPACtrs35KcPZ073/kVWZn6vXVlmmPNAgyDqIJ5DmRR
nszuDtYgo+MgWPZkKYadV9KaelkjswU2avLNv9ecel4wKPZmMmA2sPncwvbZY+kB
e+GNS11AADt+E2dVsfT9O3KG7pG/6jPvN2c/M56Nvhtv7i9q6n6fv8h1CPRy+QPi
L4sC56/lzj89xdSeRVtt8o4al8WIQdnCSoyefeC40MrxwzZIKRhDhxkZCThKemPZ
cOiZPicUAd8VJawcueyjF2UWaM1hsvcgI/wzhB3+R3PhF3aYA3nt44/a88dj3ugS
EqZUTRBOonZYR4l7Nx/DmPI5k+4u4jnKa3Wb9XoyqZZkwyXvjp2Ufg+dhP9MAHUO
4edYN4FZuZbhzJxz4I+zMUbNJpgoeos5cQ/U8zMYdMzGxFmi0jr+nrvo3bwHAdcx
2h+DcKMZ36JPiOesUkLwV9CGcDqaH086zCoyTScZt+5Bpw65Yos9m5ILELWXvwZ1
inmMjoTnpmkjqflFgcBrkpqLbUlVS7NGcFSHgFhTUZF9JtYzbswpB1ubjN2T1pwe
Y2FKb3li/10/3/GCUMmWOXOrNnfWmqUV8NHRHaJZaHMmS/Z0/7QepNShWxCopK10
Cv7LqEQcFfNQJsR3BEFGuAep0GBpmzkmniIeUhtbK5LCZ0vDrlgZjGXl9xSon9CD
sgOBvpuEyTRKc6Qh0MO7sAsuxaOZ7tHfYQ55h34bG8nuCOkDD40MSn4tQBKVMJDs
jpmKN1xLAX8p3XKTjyJ3JseGb7UJO/oWv+HfhTaCxGeZIBb9eL9Ce8qPWFRCU7Qf
OpJaavus/WyFafU2e6GNTb04x4Tjxu7MtslZcM/d8tQWvR8RPVL+IpnT/LpdD1GF
ua9YElLuAfBgqP1grvLjMwBIqzEOtf6h1+g1nnA4Tl/nG/nPlXCQrmIIUnhXiE9F
bFUjn/IMHNQjdOEFyqBb06KGE6t6eJW1ac/6+rO2e8MczvaMj6KHN5nZ/5Mm+mJS
988dqNjSCJpPf780RDGiKfW2ghj8heXK3lDj75bVQOlbGCK63iWFNBJWjA54kcBT
DbumQRtYYv7+6IfQ6Pr2PjltcJJGo0RNry7YAs9g8nCndLfLdXzH8Tcdn0ggFkxN
8O9mJizOAzHb285/MrsHSEJaO5enPOGFhBTrymfx2Qh5Y1B4NNQFm10Nx27aTD7z
+97BZHFjny5HyzzujSHiVycj5yW4QaUZ4/7mF1x6CYuO6YD0aqV0WeLe1Fy3AZPt
/qRHY9hb83+JDVgQH1v23N77ZlZpiwiE+iYqEFwAOzqWBzelsEnQISU90MoVp4YI
x0OsXlydMbVgXc2bBS+Ubai6WCmHxlKM5HbxrCzvZyafvGMgmf6GiSz88IxbUuKw
g6nWkgC21jY5b7WeMijqe1ZbirGwD0CxXgWyHJCJfJB2vauowCOGLU7nXBxiLv0F
meSiMZlXfqyNttk63KGO6da+t/6X4nYKGp2Ag2Baery2YKWUXNoh8eAt+HQ0sAZ0
Zg7n2hrMCdYq4titQlXF9WiFBX/EJIcZBiIHi8hfd56JiZxtVYVh0s+Tt+Shxzal
D2u5oAkmTJpa0hxhnZb13TdtsWXvOM0U6/z9QLAnx/Bz+jpv5L2wj5l1O+ecfKtT
wSstiAzXEkOWdn7gxdN+Ceiu0PxEV0wXQHCk5rvJF0ws2hs8zvkE1AWkK0v4CyX1
YPMtw+ZAJKlx7HZ//EWWMyUX3V0sP2xbji8C2hD82GWrQYGKdGc+AHaYhGa1BIX6
K5OKXEY/znVd2eDERK8wUFePuyzcAt/yBV4AY1+vWmyveTJd3HZE9a8a6Joew2Ta
KGCNdQQZVJX9c6N/qJBBEDpwv7guFHAyLpwP/czlow705TFGAE7498DDOUaTu/63
1KU6W0nnpYslBhM9LRVM/sABAduffk23NiZGxegEMOzSu1iiz4dhjIezM707Q50o
4WAqXVN1fecOpdJrUvE5yzziKfnz14fKyLn/N9AmtLd5oInZQ1/2Ca/AkSpXUoT/
0RzX2cEr2sPveBez/W1MmtPl2C45R8EoUifXhxOCyvJ/Jb2tUOfSLYJ2vchTRO2N
mp9+aDOhJahC7D4TLkkdzyvabfbxJIJoq53j4OHphwJ/BFOWKmQxneSZH9jYZj82
UZ7njG+E2TjeCaLns3drsx9VOxa7dIpROtZiZL0XFvo3NFH77H5e/22l4l9z7+UB
N/tIxkYCOIGA13zJ31wlfrQqW3llh9Eco6Lf9V5fbk+9ZrhjNJS8jAd7I0Xoi4tZ
35L71QcAKExyVDRUmjdVN9GjK+wHVAtpiH0y7tfY7GesYXh3MXzBYYkKEqSy/9lM
mnkgM5VV3WtJ0IPYWw8QylADzlD0wuTKmZZczNtKsZK13i2qSODYafWTHzMEElge
9C7Wf820GR7qhQZaw9jjlVovnvVe/clWnA8JzdDD9b6h57aLuuRTwm1ADhv0SFGX
NkkeLs9ws2kOGYKoW4JPZlcWlLHtTpiLc9dCabXvkYXoXavLWa6qlZsqU7UWHeqD
62dPStwMiEPln1eql0i4RsbbBibZX1p0+oS28VT6qdINzxpeYIQmlwPgPXafyymh
BpzP5F/leVJ2UPozv4CVCkhI/1U65uZjh6LJ0LrhY/AxVWkS6ze32ksaN/yev98e
8xvajsmuw+SiqoFy2PfVU8kF4yL2TEVxOn3FiC4MpeSj+AH3BNeISb8vqRZYKGKA
57jlCZeRzDhqylWZ7vCKGXoWTtxRI1TYrJeKbdmBwQN1QVsnq1+fp87dBvjMJ/fa
Ae+hOFn5XGuzMV/UAzPohgqs3RHvV2CnR+xM5JuEIzRHR+qSMEhDD5tDpii5CJAu
lmaL8TzTA4afyMZKFU8FIt2UTodgMxg0wC5vMNMu0osihN3yWK6JeFgfiB1KNCP4
pgKBT54ZCZoeQ503ETugp4KMWodTrHoZN5twdugv3vjJKzxItuYB7Mx05GC6uWHv
pcBuJ6ZJki+VoA/iezy3LTXfMLMY1sTFbFZk5K2/qhJI8x+WvolF4p5Catqn+er1
bxh4e8CnNJt6TUbCfdnfECzxPGBO/RsiU0aQ/Co/uevdJ9l2wJh8ffJxdSO44KND
NKhir282xch7hqnS2oighxzG8+719HLmQVKgJqJ/OGQxqbuUxebXyQOjPy+TZfgv
GJPqeLbLhgVPO3k5lbCJi7FEdEioAbj/3fAjE9RVJ6URZvu+jr9xaswnHCkWExUh
F13DZVxGeJdHxK8YbGqrsJR9SYJdw9gnEX3kVCjRRN6pJhEkJNvND2cCvWWXMemS
ERekyO+dcRoPcv35NyhE/6wrIHHw7ikcwDEg/otrUfAghfoMf43fJi403SI3GhDc
INt+Z1jxtVhiAAtmy84yFpQOygh5KiLO5zRv0NAW1BdWT54G/M/it8fc56nOmUEx
EguHXUez+5JV7rJN+CedBjmXY8tuzH7lEZRk0B2XugWhFRIUhiEPYAatm4Jp/2Sy
rFPgdQVD1RNcrxSG4hZFVs4He40PfZh4cou4K1zhkKJ4V8MLBUsETk+BZxrS2BBW
bJPS4dimwbLlKjA9rxKi1FsvBBZ5/pYiWaKZrl3btY1Sae1iGGtel76H3DnGQlWx
wPIb+6fRjW3ibqk4JsUykKbsxSOHiACyA/76NIZsDnsoPXYw476h0Z2VtIlLLPDf
BtzPbkfiF5nad/jdwHoSlmIHLhia6MsjcSmlw71/cG/j4e1FYLmu28kEvfKB52H8
Iw2ZNF+W5y5sQFOZzuzW9UJhONfAAzRCZ2p/cfQyKyFVh4URGJ0UZbwSLbiKxp4w
QKHY8jaihXgL+glFkyaMe9PTxVJP91QUysUK4o39qmKBfJZQW2a/homp7Ke7b66A
yrRgulTYzTrHeB6bcFY9QWxQGa+1cSExhUbohahSkDizvaURPOqMdl30vMBHpte6
s4yXjLoWMv6Jc5DBeZreizkIf2Qw7Y4QdOjZHY1RKoE3tjdiKTGPORg9texSKIPU
D7hGeVLNRMzAjeMLRBCqxejbx/0htof+HBdMgmfTGzE7Y3fS/oKr+dn0a1hN4Nle
wkScPCnM3og5HC70yHLPUeOQyTrHIR2GVNY46737WotiVLIoO78lKTjzcMa8V5oe
qdYGAsG3sr53vHG4bF82GzlO8AtL3/wtOXIon6aSmPHn2pVzC1LWeXzaR0C1saqL
j5SxHNIZk6xp2oZvraMzJavXfz9A0n6TbxBRwbwA7NoLeMWZByxc4XewUOEikSIv
v8TcJ9NDuRsilUnGB17NGH3ntYc7full+50nMz+/rGCo1WIs+AOh5XPGHE9klORs
408z/J91MABKtxbk63BwI0rIBHgtTNq1ehsxn1KeH2+optmnV9N3iwoxW4yNumGM
XfSWKzxmoZYGl0bln+OP+xSo1zW+XOGKV9GrsBZCkYeUpxpkAO3kAxASVXkpVfkH
PAcJzVBCnVgjgRIOWPxZRd9s5LlE7TOCxmbiWVoMl2IKfEcZANOYDmy0UnhZpc0F
mEVlxI3On0NvfM0FOawHkXzCJn7EEch6lLhRcPIa+NN35wVur8VifHQGFD15cG6X
90J0Wf1NBPQIpcd5u1aanpEb0vF+nLqhpa/3jtTeZTi5dfHnB5SlFEUUTaHWY+qM
jlXvEkU0hM75fyqFGXF3q4r8eZWnlM7MjLK171kVK0N1yQlaP0qupK2fakugP67j
fucRp/E5Tt8n87exEOS57QsYGQMGTkCWV2kkgu8S/EnntAxnze1qDmALKje6GNJo
zVc/6p8U1qS0aS+2sAHcZIUreETOnCwIamVKLX+btv+tHHl2J59MApyLJigLXt+X
xhad3Lg+ZbtyoLfnJGR7dMDobXc5On3ASf3wA+ws2p24t8O5hpCzsNgfKDB++52u
8olR/nX1eC5cMJDmKZ5Xkr3i4Yai2twdIx0AXLHKJNk4bXOUgmeZf9Su/kxtsI9h
Osp+vmtH56h6Gq3FYuyK2VuL+Np6Ms9Qq8z1tz3TCAQom4CDqn/IZBY/e4zPjJzw
Ar8whUZkroPU8Mf71OMQRMlrb0vFlrRnFkWA+NkbDIM7HzoQJnyXtFrbjKswqsI/
8a0gCO+n0FdO6AC6piqQvNvoHOjcTd4x4aK0XGoS8Xyx7PWBLmZ2itmeGwRkHYwA
xzGvBPWQiDf0LYY4laaBK6mtuGMHdodtAOhg7CDi6utIJUqN87TdKdrMjvQ986mn
kvEerbpnq3Hsbro9eY+OE4RtODmYjmUMWJGeZDtEEZZv5y7itMs4KQ9nNTthDZl9
opKhh1Ofyj0clV5qTZjXjvusIp4g0vlN5X+LAysV8gZfSp5jSYyHnM5CnMEexmKu
vmooCVCwwilmjRK85Y7PjZsz0G7316+1hOHoeQaGIYyHnajjKZuw1+Hb9KdCcOhG
BD5FiO2X9RrCBgGvwJI1pH2QkWQP+dk9ilvDGsWXK3aEx6aNfn5ttJZO3b44n9Wo
7GNdtjeiRXGS7Bcf4Zz+21pZEIbLtSlgHdfxvP31FxPI38Tea0zJ+iph1BK37fX3
8mjS1nRlp3VGP+V6lf7h0HQjYwI4KPzxxVfmxA/u/iED5uwMwL8pj1pdVtxoYUEO
0mWxiJjAuZk5C1/Kvv+a4HGqy/TJP86wwT0FcVbgku2GR4v2OPusuz2aYfX5Ax+g
pEJ+XNLfBXnPLjLwtSClPerFepgZjqOTo5aGEgIayFflm3tTKlalIwPt5CROpYdn
NVjaCafFMnSsbgtzIUrBRxG5sQCOmqYEQAl8aqZTwQJUnXtvEafmDCe2CFiqXfXF
bAGxPa9pVNc3052v8CgMMDfOFWAMM90qxQOcn2NOXJ++OW/Ug0HWrqP8/yUF0AwF
0IU7QQ0GB/6TFMPcyz71ZsNIhIS6zYCpCVa4Q2pFpTi2fpQOjTxB267gt1zf804x
HWJ6Lx7hqf0uB1UPyqZnSll0WIlXy6v6dW4CXTeurHZBdWIVk7/e7j9mif7ferZi
eHX39YxoSgm/twa7zs2NOduLJ4yKXRE/Lovi8DxyLVRpgA6FbaeEo4R/qiVa0m+z
Gj6EVwoi+O1uu7K38HP+9aWj70r9+r9KerxRwhVcnA9DpHwcJCTrxRTKvv5JL9G7
Cjl20EnsyaH5tirfjcTdDvq8t6CYq6qPvDaqpFlktnTF4i4SrbWKH6LoEfVbiAyR
oERkV6wG4toCImpm1xB6fOvZ2fX5kWvA1SwhS8fSiUFzxo77qDJsQyh0YBl6aQkN
Uq1IYEBGMQ+QeX43uVgg8tnzMw2YTyU6rsedjmnpNSpQvRmAxAchZz0pbcvW5r1d
q0I7fSL29qlWz0tbFua3Va6f4bFkYfWMBWhkXnfSQHmiSjStS1SQpVuh2M8wfnwc
9NgCyAtekBR47n2wXiUyxnmJN9uSf0PCdqHuydMSrZaTK0c2PULRKiv3GCd/TcvA
jReMxLX3K2QL0ZV5KP8tqR121kva/nhy8AywkXnunZEA4LpPOnAvxtTGz3MDNtWi
A0Bb098LH5Z1kfJQvGP+0NvLs5V0X2DQoiKMeRhdtq3OzRSkQS5r7IbMImgkMKkc
VQvqhoxFFkAQgmZ/EbWzNmcsI4KaZMNuuslhtZ4xd9O9lASqlQpbnSAHRP665e8K
QaUv4UAmJCMx0OrT886TT5W9pxD9yEiL9tIBJESvb2DtD0jdiwvdeAJBpkXdbht7
OozDxrBV/06wPGFIs0x/Ns1L09wGGFhwrxWFt5anmTFyfxHBMPFe+U2r7uOc2sTt
WOWjtLOeREInmWFRY8HeROKWRTZam2RB0ZSBajp2KI41cV5gDoFHpiVjiS32HFmy
/+Qfn+Qe+58UYdYAw8kZD/H7mm4jP1cgltcyrJ/dC1QWNF4bka28BASDli4GyQpu
M3e42QWQMC4+S86cf+5OsqfJTzbMnVEzHHYzeG6TSf/yk7IZIVgoFLQEg0DwoaiP
unA0MXEm0K2N3prabm9kNz4fk0CoC+03O6AC0Esl0QxeX8QxrXtHhKq2p0/kFJqZ
PcNWhuBqhhZMai5cEK/55EnUEF6H+cNVpwKYviqMNzHKh8g+UOhiYPDyV4Q4g7A9
fZ0vk/9GB5Yn1v3LnZPpuuhoO2Eree8vuPy2mK0MZ5KIkIIwY1DXiv91kmtj/Mmj
CXwBU9eg3c/bZgSh18LIY0UJrOLeyJZ+n/A/qQR5z1x3CaO9GOpC1X/EQBpdIuh6
xg6NEyJzKiZChaMdLUDY7S9Kkf2k95K9um9FzyfxLvJnPAXXRy8LjP4PhIXiPFSH
WCSoULdMz6xeo/W1G9mGMJu8XNb0qdzWaHFhLsNMvGA/VYLhzAes2I+3TnqFMonR
ocDQNsho7w8ovY3ZiTq1BtwycPYlESKXeYPOguOenl5zTtT6lyuMUX3qeDQnoWj/
Zcj5l+o+gF7bW9rP8+dKRDaD9DBa6IS7+fxouYYh1wgGgzFaxGqXEOTwk8ka5rij
KE+FregPCMKYm38WJhW1unjpzx8x6zebje6JF/a0EdhuzN3XUS/ayTtZzm3KYuNh
sgEj0/c9v3nZRpTEArCl7GHYV9bl9EAssJLZaP/Ie3RFXY4dm/3A0FVLHi9yV6nX
qJWL7TZSQv7Z2/ElJ6qbKzRtfPMkdpG588mSEW427C0sgx6q+ky6VL0ZmmE5hpyK
Jzl3LGB64XITyVhAbnWBCB3r5zIifOxtkqtkoZ1OcUYrn/NnSSdXQfMpqhP9Ymsj
ZWB5BMdYmHBEkY1AB+SJ/mgoEFtw8IBtR5YX6PGf3b/dNWopPkTczdmkWZJTfDn4
iew4yVuJOjLp2riVkHVJSUGFo/XE2cJnea7RemitSsQdmJ0f/PHj7g4LwGyDR+jL
h1zSPzQmxVnCn79Lb0J/wNc+YSU3UvlsW1rqNT8kaj/kEqUBA0Q5Eqp7Nl69bIYY
FYLUd8uPOTd/d/aaoEeO+Ju5966waNVqIHuNgAfhCrBFjfcS8tMx6AJqurdbHVlG
FNjU4bIshAM4cqJPyw5VfPmnNC3n7FrvmsEf1LSN6cULo9UMC2VEFPw5ZAy4YkIW
QKVPFsdqtfy4sDDvilyqjAQGikMcSGZYWMhmLQ/jAlNHEkcb6DrIT3CAGtOxD6Rx
1iOgdtr3wQTZ7gECFW9zBpNwnsiRaLFf2bTRiSt78W8x+5nmq7rUXYvevB1DXJoC
G+9EmvyLU1I5x2HJaszQt79M62vmvlSeeVmtBMPfno16Ch9cQ9qN8mFU7XOWLsoS
T4J6jpWeFDNf86arJT8QXH5qCJidK9hmLoMjdJUsfbVIjGTLd78RahR0ej8BsYcZ
NBu6xlfeK0on7+IGLRdsK0wZ13Gp+LVs8/+fr2PNMH8hdKGDdOd1dkV7LNseYgUm
Y8BqRW8LfSYVQg9gA8Oqg1fY2vo9u+oXowZAxPDbLSsruqdtTeq7sp8pDe30qzkL
+whmUZcF5lpt+ELwDN9owDXXUl4ETocbPV/8UpFLJTFZ7Fh84CxfK33lhjJXEegf
bU0MvVTU0aqApPdxr2rhMOkZwgjc6uct5XoLW2cTvpC6I2zW1CDX4PPWgMruRlTC
6oAybZPu2lTPdGvWmg5kL1VWK/CGt6jrBfD0hfL2KNLm7YYF+FVVNETpvJSocysV
Yl+l7dklD19ghOEJz70R0/TGJpoQl5QW/qjqS12ejkki6co7IktT7N1N4hVTEIrX
NjucGFNkEESEXyzSEoaeF+9sS9Pa2wnG5FTUadBBkUd29YijqG3tXsU93qrBzMK8
i9HEVCeEvE7Yzev3bLMzWvMQP6z835jJdFuqvNktco5eJnN6d3/JFqWigVpWPDDt
ytTWgPgP3XU0/Qxsl+3jXfdOnvI73KqMOj6byclgEpVjrRsZBPsG0wdF+P8gjPe4
Tq+lPnSLx6hCNsZvNrWsHS6pN3GLYL6bE6ZoFFvUr1M6WqDheZUtAGsfMOX9BFOJ
CCL3BLL25Uy2iq+tycBWGEI9PZYPxzx1k5NyoWeB35Dhz2rtRuItgOjmjnn2uJ97
Ni9QWB6IR74UayY1gAIic8KTWQ2jU212JmubvLagTCOzlV5dQc7MJ+uxIVwVl2os
/xJGT+3jMtYTBQwsRB9Nrx3LEe5iTxm+YsJomi1wwnoMFhCQB6TKrPUnSmMW0fpx
4meup1Be+7nRj1zjRnOdcLIB4ZdNGeNTtfKBvn8hUNj1SdrkjD3pZJFkP5b8sHBr
JKfibGbysfUYNGc/IawyKdSC4zVcpfLrymoJaGGR1S5VHe4xrZwQIMgjmIPkWfnf
AJNKBRemkxOD8A8WeBUqFxs60ZjokWOeqkF5cEYe1zQxZFa6LWUHi1NlVY2MMUC+
5MRpTIY7ZYRfYQtWi2ydxVc9h1osy43izxlw1TgcIsCe/d/skWZFuwmmKmqtiA4N
u3ixKinEXVmrhM1zDux+ZjyiCPPOJgl9ikAeAogHSrPcZ37yBVROGfncBtBGzg2c
5paxuL3rCemyXsqvEADa8OyvDfqJ365Lx9b/hajbWiPSaIRsqe3/w/NFHNXcWYcW
4FG28WVzJJqTOkkLhb+jcaTXSSJhQmhjrNnNViKCzEri64gciktpHK52z6sNtIGO
H2AYZwWp9OUcIP4lE3p8Hi25QWmY5iZONT+99Pzstdz6COcCHZ4nld+chRZTsC3L
pEgiBvmH1nv9xElfCDubpaaDq4Vh9GYRmIr4VFwrUabu5SMmpg+gM4c5mNbHTQMo
FHlQmbh1ORd7i4mXqybbW6rUFUb4AL1AWyjRNG+olhnBYiYp51upkOnTI7qoDGOJ
NAYe6sxeA41stOv0QWutqLy2N6wIgmLF2veHKL5+0pb9Dp1JHE1JH1HUp9HkH4xw
ZHZ7GmY5BKIIO4NBC5k7vVTB4Kc3uKc340b3RWJjM2ajlbjgTHVDdhUSklgJJoV4
CwZGPazgB78rIqmkJ3Npj1KiIphdnrlZsm75m3R7BGSygYEwMFzpAtFwUWD6qzBo
qxgIV48m8u0Th9UdyLdcm2I0fh3+KiK2FIMANLwDLH5YYYIJp2wnYCtVbrU2P+CC
Gf91F9TJ/D1o0VOvcHOpiVXB0glcGNR8IXca6ncPeOOBSW61FnkiafU9RdE3c1dC
4vUCu0drrTdDI4bUH2m0Wf37qFqda28nXs8qw6FxpNrg7VuzXqZSNZ6NlsHiMYzW
HHUF5wUTXt/2quU6kF/95DQnROhNhXoitCqTQchiCIzN1AV0D5itHMZ7AfhiM06e
TYSW7ETjPk8B/Vrlf19bPMgEqOCNIbvPKW64foOWqpsH399vMaPv6sGBLJxqaECL
PUTMRlxSWFwhbsJExlcruAbsFE6/f3uFiTHpEOxxvS6kr2DabftGC5s+34SSe1uW
PuqrLkDK+TUpD5+bfn2QSZ7pQBJgWSTmXNJ+1Xy2nV/c3f6LJ06RHgb3TYoIHAt3
lTe+CtN49frCDWHmnHiQDNZyudjaUJuLTrdzTzTj3Y8U46uvAJbZvV9no8gHNOl4
7VzDwBaR+fdxKwta3BcbJYuxGJruSI/YswvXPeftn6OBfDgFN/mzttmt0kZdOChz
ih7zZvmTVWNZgxBdbHTq6ZXPHnw9lklqEaTZvaAFFkDO0GTw6mQhvoX1yt2KhTqP
wISyiVXmuxw7ZCxwo2vL8ETEJGPfJJ4XhnWnNoCmze57AZ701gSr6gwj/ZwkPmlT
+O8Ayx3EKVlnhlFEq7B+5GuQvmeCkbBbZf6pg0jWtp9bk6wHgKIE30TT+NcO3t68
c/yG1SxKhRWX9s9TIbXV0xOgZiRu49U31i4E/UbLF6WBV1xuLGIeXpe1atoCOV9Y
Xu5OcQqB3FJPpjidtKJMCktCVm239QSHIk+KneaMGhsBkXBBmAdCW7T+BZU0oKW0
TjDlulB74g6N8kOCwLGSr9EF+8HWSso2wqsvAyd1gaTi3aU9T2kSwGQGUXCVYYKt
IK6EWvqEf61eImqrpS8ALG+suDzptaS1d7CMPTvYADzUt5dc64IzHfRX1MqClA5X
XLxDtbMTg6dX9I0NiCHry6kIG/AQIsxgXE6Q0/fR16WmbWinsQkeC6Vw+Pw+L6zi
P+i/dwmmQPvweli6XChN6T8doKp9eXHZjy0OC8cLfc1U6Lq4jSLzrcbeZiQk5qEz
zipjFTdLtBzal5UN4AkrEpPY1Z5+9pmcB6cOEN4x8R8LD10OB6K97RtNHH1SRrSM
XvD6JBDAXheqjVLjyo+rQBf3fv5xZeuPpZ7By3w9ruIUDyPj8PM7dU9aqdA8h2dk
d8VeaEZlf6SVUUIJIqDg4GK2d3mCurC3sXFhR/yTM9J/r6QPOddEqzMQMpnpVB+0
r0fpGvkBBe3kePqrsbCRZgn8J7lo8SvUBeajqrIKCJTUXMppLrhxemjcwG3JuN0z
ZQsWXeTeiU6lbgteAi85ErojVsoNpivtkV/1Y64++NSoQBEXORIoLeIMxWYKHlac
gi4eIvT8tfIwC7XDTFH6LkgUSlFJ8gBUT8sYr70zkZI6dZKih5Rmtvw3qC0xyncd
1Row4cheKeEAy1lXKSQxSV5WyxGzzQ8rjlL3jRfOK5w7Ry2B5n9ykSlhj+Fl2NLF
MXxNzIUAN6yF0i7WDOG8ugGsBrWXqbedqGX4VT2xfTxAapyUIIxCEDgYtBw2qs9o
ZVZxYpCplylPHYT77xA1eAujHGm+Fab2SULQWcoMbWuI/U5WoEVwqA4IujxRLagf
6Tgy5ohEDMM/tZqyEaLixPRO6f3Q432VyFC2rkeXF9fXGX1kqRvcfvFnBlYR7kv0
LcDd/367IgJnn8RGLRI043jD9Qf1zqU/3i3oEnd3aepek/KI2cxAmuGGRLvdIYTf
frdcm5KUlxqog2QoGGc1VXWErta/osnt/n1AVxBqvXopCdmbwqisUGUWb3C42lfP
Q/cWMpqsp+8rNiYMIzTJCMVlaMEKH0q0JkV2GYZudKJwi6vEN39AdhRefC2GImqZ
UTdS1v81Tqn1GvAFL/vRfIBdXIAinDx2rGarOcBiPIJ2GU4UfsLNZqh1HFfeyil2
L+H6rX1C7CQtdglke9E3X1/dADee9ZgF9rQR8vv52AUl/SUUM4GG87PDVbYoU8AO
+yxBuR5EbiQaMGhvdL2VAhA/178oxsZdC7zvho3ao3fRVkors96xkKATZrpm+Le6
Xof7XAjHonS8GZYDNLPK0c9nJJaI/HlIU69rvfsRZ4fuOB5TJUzs3SDa+PPUUHgK
qTcW3o9Xzat5TG3P6vyGbZDWXIKVZBQpTBanO86EYij/N7fseP4zcNGM9mIBOOhH
nDoNR3ByvTW2W9P7badhxBWo/6CsnNTJZmLtIrXD9xJa4ct/hx/zjOmXJVajG661
0S64zUqJkgzbm5liENS8wAVl7fCIIhHMtya0Cnx5rR3MAt31vPWMMmDgv9Y438Od
mS0VjNt/G45irsIr+6YSClaon3FgUpMbvvLdUBV+TBu8W9JuN19Md+E1v1b4f8Qz
7N8hURaaRHZB6PdHqGljoDV8Mta0uj/kpNBYJtz3Pur/6cJFyBZop8SzSk7rT79/
pq5QMHifXlgcOy0tcSz8P1HxI7LSwCDn6wtGPyEWS2xJCrcppv4TTuPWVZclw3Ih
9yo00R+eZsPInYxt9RPSpgSUFZ9JhMGsEPmGSUpO88rJ0QFRAUh58d8hRV5xxHEv
F2+48PSnIjj1F9xsjJOCyHRyAJ/AE1fOS8mTFJ1+mtXO7BMlmDCnJV/laIp8jdTc
k6qSXs3sV/2igjg3JTFwdXwpPNAs7jniCE8YUjBIDIG8RXStaKHddjvtQoY23OCN
ZtEK6FSznOQ4+GxYsorZRTOMgCeM9TUGdOkjwOFeCWl0JZOfp93VpylweCCRW9BV
yN0tlmef/OF9yP3aVhQ+qo7BlZI58bxdpU0Ek1QJB+i6MKr55+zG+StUeQ2gPnjj
gqXsPc/cbmofTuAV89wD3HLe8wqRFG2niX8qkX9YkChY2AjzG1P0IJDZTjkW1+9g
GzKpSEzep1Wpxo5CCi5OfW82MZ0C9qeCdGgzzIFQGLt2jCxhtP+d4rEZcG5N2rIn
gbY06zgngGDHgrcmyStDpfsqHO43jHgzXfGKbeZnALI+mbepXSQ3p8/kblVmkbRZ
FfGHI3BAVNy9gqEEjX7hqkKCkr+5P5hxVhcXCjZ4nKYdazbzjDwQ6amCyzeJUfjQ
/qcJAS9HujNcApDDfc0TXtinWpTHqoNqkanP7hIeg6dTTP7iX/8c+n+yOe6FJ5v+
q37WW1mkrPvb5njUyDlHYp7FSV+/BUfxboTud+muru6J9qCw+mlKjOnUe+tQyfG2
umRoQM2iH4cDmVRtU9HIZ/feKZqh0lJSOmnPZ/rAzs+l5P5H1kcakLXYOh4L5p+J
jHCHum8HCeBC4bvyU19AFy8jOf0D+ysZHU02tckI5apvfZxVp0CapDZ9le4iuuSj
1t/sWLr0qTgJikJa6jv77s5GVP1oe+Y7U3UG79m1B3VSLewzqyUp4F4RY6vQ6R1z
LLRntK3zzc8fXc9RnkhIS1RCrly6/FN3x2ps65BbDB6DP3IK5eOzBUpGohccCRKn
RTwlN2iAGniPW2RzBk+jVQCbmnMFIqVRICeIuU++fn1qBkLm/Qel0xd+AchsBjnf
kZ/PU//ifLi0WejaugXebvNds+8m20I4iCJYMk2iAcgKp5WYk/TphZ5wfJ7FNkIH
2Ncpjg34/Wjm8c5iGsKfBsSXO3/6eyK5jP3oqmc+WEAQcRm3nPOJgXwWKrsReI5v
WgSKksqe0vFkwc/4K3I/QiyVd2ubAI7afMfT319gTCZnGybrb6e94vjtadtIrW6e
YEZmDQx855vc6l5qHUum0i2oaARg32eol8MGXZPxhfdbP+KaaOohmW1+neyD1ok9
kAZYrsc1ydxccpSUY/92MB342R2t+SU87F/ykgmfIJNbCxtDOxTkayonhF/2QEgR
tNQ34ZSr/dnqBCR8R2d8DF17Ix3TsGP1NiG1inVUD4fafrDUBg3rUOO5/5hz4NAR
8CWU0bTbpga4mYCNNc95ZYnqU2lKmE6FFQ3nTOQ44NoDRSAPPzyJEXDnCcI0wgwp
IrymEs8zCrRMtse/nItjukl6J3PXsBAo9fOwJMFosChLSBDKo7rgjNf9LdSJFJiH
iP/gfYYzczRITpM6BpxQYJFD+aJZNkiUFiBuoAToxSYuEUtP5QPnECh3+Sj8dM9j
9oQ9OOkciW6c8jt1tUrWvTohw82ovLZQge/aF+WQc82A+FO3dsQpCCB+YfCHqXr5
+7Wf2jSeNncFlnl1O4wA+lRtgEqVwzlI40+6W9JhndZe4g6nnluYe2P71tpM9+kT
o5mV63kgbk4kGpavQJYmSodinEUlRY7n0KPf67Z8XjEQINIdR7ZevpOFwfaoDJ3Z
FOXiAEvFxS4aBLpAQYbb1q872neReSxaBW00bXUaNYD0F5hiaNjncAf9/5HzQLtI
zdtglGO8471FtIPio7BcKhx3rN3sYfhg0ds4n2l2Db7MzXhEA8WYuSeCxnQ8nPuK
mjmBFBsdKENdytZM7PZZ9hFUypMdJskFKniMWeemN1eE06mKmNCLc2cfOwwY0RIS
HNgqpgjILJz/tg8BesGmumeEpTGLI28Ft+YjHoRDxAlx4sX+ZRwBOWqOlhX/8cgC
LTCjuZcXFPVUlcy03rpkz/fzs1oIKtTKCSsVnSbCLO36/K3zvSTILSAJwf6iiT6r
c3yR/XYugfzzbV66roR8UijV9tX48oII2Br/0ncgUiHzgqih/JPY0nbOXbfTCPQ2
vTODPIHCtZiC0LJbjs4C6LdrnFofl5nxFQMeWX9/lmknhRhNMKsMKyZXWR9C0Hgv
HRkKHSI0t/41q7IuvM9NOvvxPwt6Covb1Am7E+wKxwhaqTw9gHY4f2IjHQqMJ55A
0KAd8Hjzkmzf+X6/9zArR7R0xEBLZ1bdH4LJz6tPkyJ+x8UOt5s6oBLe8Bcq4d9P
vw3AGmOxOm2g+c51lykDOF9iKSozSvx1lFYOThWHa1rG/oldZbe+SM5KY6Mgmvat
msttzGSjgI9LeWDBYJ5fujBWIl4yHedmMk59J/Zzz28T1jJi20J1CJ5VykT1y33t
LogrsaRgUtTd2fwuBVV4KhnIUdsehH/3lnirdFKjZdVwnAtkoboQeem8LqNSqVDr
utwP3WxCTWHGJNQUK6F7KiTEHtsuZ/Kd2UKPfwGW2rFbkKdiBREmsx3v/5WiSRVW
bG8/IuTeRUzykLEPvQYdBLuoMv9c9wUupegA11siMAQKcIX6ih6x7BuOaORmeIFl
/WtmBkmSuRHl+ane/o5ANIPSaA2i83JkxbdEFEO1EFcg3aN4SoQzJx8ixrL556w3
ymoHg0ZR0yvG1vw2qOWDIq7DbYW2WvN+3gDrIIHHGXz8GguXj69aBfCLREEitNz3
XG2oM2NSVn6LlQ/vqlYOpVFc0JGT80vg7D1M+iWPGBFvP+EFbtu+oC2zRKXetNkf
Wtd0Z6qn4hudDhGKrpK77Fcm9RORTHdsF3KJudKCBAK8wVfkXXGxipM8ra2Bj9gv
QM9PMRjF43k2q2Wvs0SPZN61bKYz30x4+u7c6cNfhOM8omXSm+LwPA8eIug2/8zK
S3kx4qmWs50WqNbLazkUy9o1peQsqKMitKlGthcbd0Jk6dw8wnZvAFKC7Exe5nIr
iIOQEfdDwxp4FKk3riwQxUXdxiqrPdwSw2ZQwGtgV2nTNE2gGpfQ0XWvYEN+/NoH
LM0sx1FqHAf4flb41nuIIAceNTwK/mR8h4lzJMMEOShsAHu9+sS7/o6coHANdb8D
uV3GRPIR/Mk9/EZ+hSgiPGr6ej1a6nVnvmDWm8Nv8D4qPATBowdn5p96SMEzHUGT
5r1vMJ8aDjnfgxMD/7AwXWeaXqNnlIeTobGAOYttH9AOtUjQ2D+pQB0aexaPYrjV
DbtgVK/Aoi7hN4cbvmllShuyQscm5EBbu4Q4W/b1OTyi1zz/kvTEZ2rQFyHB6OJi
4/zuPvUJbCYuNwcSqEKgJGpJYJCIdrbpJW2S2tZPO2OMxKnCjm+2qv8pETIKIH9c
ZjW+/zwmIA1BLtMRftTI6vaT4DHmlucg+ARqpLCd6f3r07kQCLdqNb92JK2NFn+i
qXTdyP86lyhsDx/YjbEGtNTisrrF2TS5kUg/qEUBae3c8VHp/kNkvEfrm/okZbwD
ALB6ROXZCw3gruUR4jifosD/Y/S/VVOpY0EFWfjWpnjABf2AoTfk7YvbCLwRfl8s
/eWXO6UT+pFa3GgnClPRN+HOfUIxO/hVvwjgF1qpd1GL+dqqkqLdYj00IjD5MR18
wxdL/IsQUVC6HBz6ihlAIrt6qxy/BDBZn5ENUnarw+hKbYgikWQUPRa7ZKOehWHn
edIKBP3BkGB1UR4TCcJ5zY119j98VCadgopH3Hd465mi/kUtvl9qC43rT7Pb0QqA
qS9SlTYfKRDaVwU2VFuLIa+/0my9Y2/oteBzvEEWEwoHfFXYwgYLKF/Lsc3ii+lc
0q2d/o6iEpoE/Ae2bSfTwUE/zHOsAswj0/rzK19os0IW56GvQ1e5MJpG9uvj/SSH
fDas5nUV1DYcIW6TyX9Vke+chLuCjBnqxhGTSCbdZbNesFHBVVdpghb+pnn5MVu2
LxIHX5u6OPsKBhWZ42roGUQ63vlQadzD714n6eqSgJjN0tkHgT8ksB94P6LIa7A1
+53OAb9hv9rknLkpIdJYnQxl5mH0Gfl9F1NcLYbHEeEapfaOVTxQuAYn83AEsO8y
hWDvRhlNUPBKQRwZcSEUeWUJNApZ7MA+eV0lsPlTjbLkohhns+DhS4D3MxMtKYhP
6NrlBjg65NCjs9+LoKtmr8yMWKCEleqBjFMk0rvow1keFC9JQQJAc3nydcyItcon
xZ8h9/k4LUw48CkJass71rSIECS7moJPQbHH9lEAO7Tr7H/SWFq0rPg6IPY4Yp/I
1e0kRULGVCfNR3y9GM/OauPIHo2yW9Gk9GLqSDr92zOVOPp0An9Sql5AY7cBVr2p
PPEZYhuB5O+Pe0jjUi+Dtkspo8ruLhw3SPfSVHQ9lni+rfEQJMB0y2guf7XGkokt
E7JQ8awp9ZuAKrhsf86lbVIdy/1f4QCNVExS5ucnxYm/3C7nnSjNkioX1yxS//RW
foaGbz91PzEJ5LRgcyWKhv5cyyJ4GaOu/kLYHjLGoHr8emNRFPNAPMNvttqvNVK2
6yNfdJ6GS11Nq9/Y0v9QKXyjkLqwcijByAYsPDphFvhqsXO1tRdU/WJawEvHjvSz
73V2bCC/+AC8GrfTKJFVOxuqTe9G5hm+Pn24J26cdqKWA1+lovd8VimkZOXDeezS
bbqrxszc+GV+uijz1oX7b/ihY9SuqNAjekN/wijv+OXq5NVy2onu/NtKwZl/7EF0
udbqs+yLuLZOIfKIN6EKivS2e3QkOpvqJrmom4wbAR4Ovhm0B0g3W6Emer3Ih6Hs
Apt8SWh3yzEk/JgHY2qFk/VgT/u5OQ/9ESpB//6wDbSZktvvIRge5fH31MDKRPqQ
fBub7yYrDmMfnxghoyrvQths6ZjuK0pxbA+tQYSrQit5BxAnqSM2/qwOCl5aNzpH
w43yzwPmwEsB0neS5BKc/fYLxG8R4pT2Xun7ceZkgLWX6CtFX3wGkSTT15lNq7Wi
VZOMKo8x99X3i/MWMULa3EUXN/EYN7T4IQkiO35Ko7KUCuh+Q1di78FMf1FLh0u1
4LnwOmsqx0ZEGw4GKWeLXvPey97eSkYWXMnXTDfFHY4D0iwmzo2FCDf+2ZMTWDCd
g30DTWsmIgCor1bTSnAMyiTWqtHxxOMJy4r6Oiv+ztPhIF1Z2jr48x2lWMFZAIrl
GN9+O00N2WVPngPZNTg5YHYmIzOOzj0BI6yAAShyd+/ky7iUis78hY5aa180o58N
dqVYMjXl0bPj62nsccG1JmREobVL8H2oOP5OeA4ptK/FaMn859B/g1c7NzREFhl9
Y1gQlYy32PeIzepTnIbPVr7wNhkIp5YTs9IZ3f6WGXLYGHn/NyfbRKZf1SvGX7tl
gcEX7zpWGi8IZyJSMKgrJz6lBxR2lGc/0npuVCGQuLl5XaOSHAKic4oKTAI2Hn7z
qCmusvhzqTJBY+/eFrhLcqRCRNE8LWUM1CoAfLnMoOmUReGmcotNugW3dssb2afP
sEDpr8CEz5ZzocLgUEBEgY5uTlZ2TDnLByYDeymItuSm1FNnaJ5cjatpjduJ64r9
0HWN/bMTMp+xdFp7QZiWbQ2QbZxD4g1rRP8daCgVfmx1zThFZExcNwqzWP+EDetq
/lhxctY11AUR32n29YIrIBSGiPFXspVnC1gJcUwNtztacw6CpITjnzsgcLlbJeMM
A4l6HAADKKgIb8r2I8vrCUwCCCsKhcyF9xSRrNczLxep8m5t5Sr3WtocOjc1QcZj
/s9K/Ed4RiekKXl877aW7jz6SK32ISbbqo1EqLUt6927o5xVtPiIeLpdwLFlbNZ+
T+RrowBvAb+/Ok/BRThdrQQX0rgjSu/IUBD7bK2mBaINzx+8m6HcdbVQw5I+kPMy
Q56prPgKAkWIL7nOBGT9efnWh6fcPuyzDxgFcXeNAPREEzp0B9kVo41g7TssIuP1
IvH7XLBLZqu2yLBAdp56Cnt4KcQn/uwvist+8mENA1YaGsWSGbc0znRU957pxJo4
4cX+8oNLZEkylqkac3gFSMQ/UAx0hbJDWWv9We+4D28gzcR0oOBaXb8+bd28Wo2k
zISfe6r06VAGt4iqL1L1NcpQh2M4cGaRT29qw0OyUhX9NelAkG3LJfa3YR6Ykmos
URFd6Ar+Nyd3pby0teaXtj0ML3L16KhJqvB4xfX79/mIM2kbkN4iMiJM9MqW8AmM
YmdkstpM/OkK7G/0YZNt7d2pon8Gne7UJ+zrJ56tyXhq0thxdxcMFWKfzmzbfHf4
H2OqHFfpv0xzjpZn65/TJP+8MnhisM9IcnY+DmIZepxy6ryZnHIRi69mubQ095nx
CKn1foteqnzOGg234pYDqyZgSYKTBRDfwy9fkV7T4WXw8ys4RdmF64j6UGsqBT/Z
m8r+oWwEPVUrbxYJ+vqs8o2cbJe4Rsrhhe3L7fH69j7yolFV77CxcShI94mCK/Lw
hkB1XOQK6L8sVi6zu9016eN+B4miYDHkP5+t0FjT+tQ6KpYT+gxLGlcAiSGpaaHt
xvYjNgeLga5jhN7UH3FiwnleWuM4dfH1MI5b8SgZjdZ1geIeEbtRgzF4wCBbDMqP
nbZdHIaPRjgfvHLk8nHKTGdoX0XRJ3xAR0Ip908VjOVqlPkpKFosDM2o9J93liMH
Jh5dkgIfO/pFJmbsc1bfbR/InMCk/8D1pW4ixNw90oXjP7+AbaJiDVTT+Poy6+b7
HtFvK14rb2EHgM7Za3nH+/HpkI6eeP0LWmeL2ATRSGMHvwBfkWPrQ0JFdJmnvtyk
vzKckkVOzYSN72dj/vkWTEDeV3xFxpxVsjZdEG3f14Odb6OZosYgcpUTVZdvawSN
Ejzd282MJxv6egpfBTwqJ1WC10Bb3lLPGj+4/kbElHQf8X6fFmhvtQ7sOTnGRSUE
vvftQ5XHUs945iBjWNj4UhdIRPEVGVslOkS/ArrqAG9EI8TArupMtG0Eb7s2H7rw
j45enB/ZPbCSmqlxSTBj3vhhlZwe+lNLIMk6UJ+Uxrc5qEvf6yGJ8oqAppLmZGVw
5xwlnVt3Wuvzoi5UetwtE4OMAIgyIbys77h/85zIBCnFgFijUvL9jVj81Olfuon+
oFn/hMpbMED7DmzZSX7doEWLeUGeGYDiKTd8AyBEhs/X8xQ6GMUNmM8gRu3o7fiQ
KGFH77kSCCGRnWOGM8GLT4xt6xIhEBm8JtGMFi9xRrkYkcd/9Rv0/1eUOsXpyjwN
JKZiFLAGmLfClwcYT935uKyHRDD1IEjqcgdp0W461kskzSEa0agUSxcYpgr1fjLs
ZXrP/400IgSx2bLf86cFxxrrJUw7/Gvx0Wm3UjOaJJxg4RozbcAIYhqB4NdcRCyK
P6TusD2Y4afWnH3HgQa3x34p/jNfqq7mOa5WCMn2KRYJe7N/kl5ZkVs0Bb5auMvm
s4DkplK6it5Id6thdfbIy3oAhFg/KNViXY9HSPqOIgjzTYxn8ols+c8O/jJW/dTU
JaOcipbJvZ1r4Z4BvnuS2grZOaM+cMjpr+K9ioTV/piQfO8G24kcyA6RvmR5AwFv
TkkdfBZV5MkPxplzkCvHcgVGN36Hgld41dTBwMSS7bNDW9IRMY6NtVqDuJJKe6dB
INqkQD3DSDWT+4h7hK88j+Y/JeHADkhCz5RJzjN5sIgZ+c8YVDeLh9jLs7X6vxm1
UbsbEaivP2kTLVSVOZYLmEpRzz6sDT6Lis8XzYopedyCdJNthIk5tgcmXB2FBMVO
DaSL9IQyM34Y0X6qlo25+zAVPdT5TDwKCtuNpER5pjQ3GNPOPcJp4VITVo3CwdIa
UOZoVdxB7nBYFiMvhRbFAgTopElBU/aVtS4VnvmnvZhN22M2jmdif6JhNACwyAMh
ukRSo0eTo2PeuvLAFmDGG0MGLH8k9cUvTgKMDwNQM0hxKb4m+3DySKZ95iOD1rWn
k9MYVmSafR7b8pXORtyXtFr5ipWRTCtN1E/67u9VVLBVfbjGq7C12aX6rrPmBRUk
Rx9q6sg2TdrYElcyk3i2JzSrcfyK/1NneUBEtcL8UiGDb8fr+Cr12s1ELrI9Bgpw
a44xfHnoyxE+g43wkU1IdVPT3olgoMc4tQZNOklSBgZiCqzEkqTKqrFTZM4b+bCE
9YUW5bOc6grraLu44iEmQGfxGoE9am7BoqO86/3AA/oZ3hsXQLYCtNd+OOVhVRt1
eowI9vdkNX7+yFKdBSnwzYwYLySxWLOiKqTrYwHbEKEeX1xYL5vqvFwVPsLwxlUp
zTZclEmOko777KJH5YfBQ7jkC12WoSgsM9V0Y2FA9ijAIIXnJPrguY9McHqPgBDO
fhvQ/eo25ZmbnzsBIY7+zuyR+npxf+SzNQ3aI+Df3yrTrAjmbHPruhFVNkMx9A93
XRp/b46/lbQuT9A6wIAUnqw/a2J68c2mizpVKpUv1re/4ZYAq+kwrsd3ySPwa777
b5n4MvBXPulf80ElxnTsycfz/642g/8dvxZvdTWUKew0hxjH6XT6kuadImm2XW7v
UhTQLdRSqZ0hsefKfJ+TaSqBEGlPkAxaOHYMuXSwaSae0BcgfRrVrB5afmeodvMJ
MrcR4vG+g8zNMAVCxLZe5P74xjQmXsgdmgzb3F1G79IubWpqT3lTWMZeq8jJFolT
TsgehF1tMQXnRMc68B39V33kZQtzXEtr57FyLctdafq9Oym55uD5T083JnMV1hCe
bPx2SxeJDg+zXKSveq1PVhV05QlbjPQg9ierY2HQRYrKnbhSEz4irQG42xvoWNqF
AW8aWlGZVaWVUKvmP0Yb5bILpZ2RZOypKy+bOBkBbqiR5pZijkkm+UZvQucGLAky
4Lyc1lc18TuSRB1fdXnMi52gz5WRMoIQwWvy29sYAF5eNHrVzY/DGU6ARkqFIhLP
zelQKcXNesOlmCfhaMelRv1W1cC7Fq0EQbNDcZ108gnWKaHH5VWJ4gEYe6vY2sM+
mTzCADtVm0s4V1Tai9qDeWicA5WQCllKS9rdxOb2pfvkGw+DQY8/yY4QZgsqmSpi
mwJ+065RK3JaSjf8ZOS0X3u/vmWq8FoYC2AbKMLf00b2XkNalFwkMpbAgmz6KdIN
9RA9nYRIVMW5g7J4JAHKnIQ++Ih9xbycNwpJbzdUD96G0nNAqymj7qEMVg5IKYJp
d1LmWmrkyHWwghrD1RVDryOmdjr1vvyCXjKJ1Duog5eKtHSjReuErCRyD/zxU4PK
ByCUmNG+Ix6eAdH+l5ct9fhNJRZHu49yGevqSQw+FpWanYREtZULlIiwU/bPuu+p
Q6/kbZiIeNtOqzMugS7c2b47rQBKTU6ukZGU2lKlMocR/v/8s3xhT3N1RxYH9DIh
bEBs8AWNRqit57ckVYiTP43vWPZ1yjGlBxRJkoKYTPOXEbn5Bx4tnAPDrX4ZfpkO
GVh8VftgGx+d45zoecVKcjt5XrniJrrN+LGIddOZFxy/bBbrVAWwSQUfHJQpepB+
Y3oOrd6ywmzbKXDYa277YsnWFecOH8WaP10Ucw0YWXhdEZGS7E/s/Oe4RtXNSPTw
9jZxOX6a2iqNwyUGmwrmqju8oJzvwxsQUofW+uRHBAyI2So+HkMvVTGpenRdswEx
h2YxLcFKygGihT7IGLRPzn9VbXKFhxcvcu1OUrXa2vIILcIxYhkPggL/wB5GRKFL
FoQVMhG7qpb73TC3PlViJnMzj3z4O/11XIeqHuTdpFJePlcQ78BF6adFpmE3cG8P
GnYqsRdPwYEsnR/qOHbndAhYIpp6Vdc/Rv2Hj3lZNHqvXlyXhz/tIj9m3T+hfSZ+
cAZnCGq2WsvxTbbFfnKoVDFFLPXX6vHcL0LpSRMjlnkSICmHmvo395OkX79S79p3
k66HQ94C/Aac/mJs1PSugL6eHZpsejHWl/4Tdnbm3aYyMubbEjiu1bBZCQr1bMdU
iXuW079XGACupRY5VVWmwo+qqJ8SJ9gy2+0VaWA/KwpvbnaoGxHWBDfPaUPiiWQL
JQOTO4Q8ym+1LG0HmZ3T7Gn93EqNwPrQcNthrTzNyxFu+ApBWraig52ZVIgdUIgc
1GIZSt/8HidMjts0eIl9ntmIcqd7SyUTBmPGAMqniYQRA+WycgZqvqhJ246FvrTP
yJyr6Hn+9JWU+nK0K7sXhP+lepcL8sqCTmB08e+iP6qGY0a1TIxbag2LzQ1Fr0xy
xgUQwE4El+wiLqmcudi/lDgzkBU9rSOtGDJSAAPoAv99IbRR5+DrcdCQGxjnHwSV
r5l4TrICwWOblolLviOIo2wahgvVow8CBb79fHIVpuWQ+SFhbz3nnbQOujyKUcBq
Sw/Hyp0Kh8jNvIl32LK/wR3nXAO2Swg2kV7dOnxAEOKkqNPJZpK1l31QgV4TUhbF
QetgZuhclkLls39rZ1o+/0RLvzOv9FfLU7ZHIiFCeUU+7rrDhKl4QIIrI8lItduk
OP+D77wRpsvK2Z+ScDKrPX3rn5C3AHBukd4zjb1ysFjXWjMJzOM+tYyttjyZlylZ
3IZnCStX1yuBipLV4k7f7CaY6hBjxe2Y8urRBgtda+26YUE+Ux1bHPYlDPuXCzI/
rrk8WXw+93505gBGZy191/2L9FTyjhdVtfYM+bK+gNZ4GIhuHiZeiomZe33l9QBK
vQPkuMujwL/RnV52yoZWjQ4vh7ND70P6vDQh+gRsydJyvYliVSTEfsyB2IMvlb1l
NNOr1RggU69E48zYEK4IoAuq8nd5cg7iCuq4XVbo6WlFdFscn+C/N5phcRci5bWw
7skfo3MpoyxINmK9H/okv8qhqjTjL3ifcpco5MT2j4UcqeTdzWziXT6VPi2kWZwY
hFUpfxpC/+DFt+YjnDPIu7YhYWHHWWaDxOkWiNNbKkHW0BjdtmObrFP32Zfc1rNQ
CKfzkGiBk56BPkEVnq8qavYqPgCLT6Tjz5kM/wu+yL9ajdRMwSm+GTYcJpRyngj9
k4f6LyiXVSZgDM+ssejl4MVhVHxXm0XC7LkZDnWAJ076ApusKgRGFKU8IaMTnfbS
m+XvAAbaVc71Rk1lndLJUODiMVWTW/CWWvY6nu2EawbXDWv3J78O61ECLCEL7jv/
aupd02CObrlErxc0CP2KD+qucr1Y2D8zyIs6Xwgr0783eOd3eX8ACPWiKRau/1CZ
P0c+VpIXTSh1VWBCmlnn0qyMFdv6YnCIKbgooNbL+Hkdw7nIETGRQWLhHkpBiF32
CIEcRPmF5WZ6LPA8wm0DtHUPdHAoen0UMzct1UQcEW8/hEW50EfTCcpsAUUHCHYk
5WhSqSO1OMeFOJ3ED8GuDKKot15zj+IexJAo3hCsGjD9YBi3uhzm4N3uGURLNSkn
/Jraxkz5iAGl5ytIxwRrwoHQYPTWHaYWjJOFoRbkh1txx0rS4aTYsDRjfuu/iKfk
39P0EZlYk2GHPDZNUFP2IruSVASYSagesm/8ADQKAJsDzmXoZIurlpGeRTVY+njr
t+16qW+7PY3depFcB4VUnV8S2D/2fnBUB9OYUarLfLu9GaIJoq9CnY2E7VnXpL5B
iT0QM7qVigtGOB0AO65v0fe4vvmDwGZJWsw2sGmqlSterdoswpWB+xqjIi/5pTmd
qs4EkT1+bIx6O7bAbadynY432kKtJawSjg4DDspBMIer+csSHAbMbrLrK30djl2Y
OnDC03wljbTK3iBaXTWfort7z5wpFl6lX7LQ4el59UnV/HwpNfzRc67/bHFCsGCw
0jX1vlhDYOw3AELYOWJuNOsEGlI18gYe9ygJRm9T7YR2WVmgxoJC8Bn5wbgBq56X
Civrtv7MQifpSkBXTmDLWgdS3lYLZi9dWxQpY9n+AfKB6j1Oys+lW+TM9I6bsyq2
R3T65ihfZ6rbVETPrVD+H7wrhPrmF9P5lMKhLxRun88gTsVWlD0AkTe4vYCr9ylI
qEkIbkCXJCUQfdAullYMHP8qhQ1W/ZyoNruWPJmd7qa2lpQj0BaF2yZ0yng5IVIc
ahFUk+hfCFVRF9/KQAwtaTtJ3sPqozB+AQyd+SlV3CZGczNG50Yk0OdnnSsBXAzK
ghiCMkuC9reXP5u9le+g0xJFEYTYzym5QujoejB8wMbiKznFtIDdxSgYw/mfTUim
P0aZkoOpILqgWplddooQy2FQGTIGqYpQLjfeG7Gd7mdAm31baZPLjoJ3ZfANR3ft
ybGUyLK5bUvleOx7lxqR30VNKYXLbf4P7zE1TbpOTXByMk5DIM9qyX8qMojtgDyG
ehKs0qlXmju87gcqZSCdDGeJyalbY4oHFGFnjHdSjREcb82QuC3Id4oKjAa5mBFe
J+Nls5SYiYZPXRr5wcRNN178DWITzKWOkpK7nHIwo5vKlcauvkBIrMOC0gPRG7kY
9Z1vm6Ou3r9X+KwQYKs+4OwbCh538hyg44Ub5PPEb4gGnh6R5XX7q/b+ayBPkED2
B9aISW5TuutNlaXN7uKZpWp+uDpDABB8NgitHOQBRsJufvm0j7HwH8l+ZirX9fQq
fj0DXl5aPhvmgAzMXKSGE6lKQs6WkeLJDz0/yg03wSb0+kF+EKg4WvLKlcI8s/ng
NA8WSrmvWJKVH39yTBc2wRsEtC74J4aqawDQJ255Q2xDcrmjzFC8gQ7tE6AlI7Oq
3lh/GHcdUcT0TWFyUn9mnpEaCCALrFYogK6bQ5I1iktBlB7YX6Ka5uYhBYZkdNRv
FDv8lRQ0OpHqQfEwrctIiT84EHVMjqnNybq0NW652N61qpO+ombGwllDICSmMT8a
8N95QdPoq96cvxyecJLxfGI7lA51pPS8rus/5jIltd9UOTlWmkYCtWnR46zAoo06
LYVgajxJIJ/KG/Bex+qcjl8bhQHv9ck2uVAHzZUAtZOX/yiN5UEYL03llAtY0QW3
mf9Bj7g1Y6+2oG3nOiFEZPbmCQ5EwiEANBMT5Pym12/lp0ncxBKJOJynHcIt7syu
pt4Uxs10gmC1TGCww7L//ENRtZR4K5T1B22rXzM5bYfVeJD1zJHNVZFpApTHCB1L
mOzML0OlnWDiJEhbRohlolUqr7UJt5fJkKvzBGIVU29EDfm5FE3tcT2U5DxBzYDO
ZrxvKkJhJmrEZ1MW7OIcFdATCTOe4ZHsMM88cxLSTnxKgDqoAeaqaIF/Rc5p8b1o
PylZ9cRLoq277bI5xgrCg78ufCowjuxdoomt+I0XDzCnZYKWQNvuMP8ug9zxpSsO
F1q2V3OED4RfRrqMXeVwFXC1D6at+eiOW+Xh0Go9ySWXX4n4BApIHW+GngtPHJR4
lgZL71GfbVYHLC1XFjlpQwpaF8jQEY8hnWGLNM3yaJ5PCV4E6hgRFZr8gYfyPm3T
nGDM3biiM2eie2+xYi2r6CIX9PVxwpybzGKNKkaWEA9Z+M764gp/m14xb7ure79O
LfAzSLpLn4lVv4OxewMK4rZjcluCtpo0yl8N7Yp4IlW/fxj4wvd2ADKA5rLjrSbu
RhGBt25tb9T0k2VHUYa2rQyLQ/gOCC1YTnaI0w4Ywc5wxXYzqjNt2sVCyT+ws69g
MpIyWtf7UVKZ0f47EqwoqsYZvFKU6VVU6GH6WWHLzOJunqkDqdx6djQuUab4uovi
8zeBdjScr3D2mY9ZxHRBnPSft4tlF9PDUcRXWYvJ5NQ+MieWbY2Bk9owhuytGgcR
BBVjlyKqUl2B1l2YxWa47KhR8w7d1Fs4FJfcqc1A9l5VTBZytHMHdDJFIVhN+Bs2
JR0bq1/qIDWO6R8kEE7tnPHUuR8J1Uqt6AEqD/WlWfORdbf9cXjlzuTkwJ5Ptsy6
uoKCxlD2QFSnDpHKePV9MHuT8A7Hv+3Fo0LTqEdnoKCyWbHrWDraItl2OXEGJzuL
uaS038VIDdhQk42dF0pMdS4lMmjGliojXU4qqZWIEX4oYjig6sPp9J6D9P0EmGw0
J6i/enKm8Q70EILHvmuYNDwWijRNDMMjylqsocmKcX8nkAvvqMaV/K4zSgGBN2Tp
Z5efhx+9lZRBsGjR7TXirXphPbAzzGjzIZEiR8qJPAutVn4EnRt3Nu1oP/0SnRVS
QGeZ7vc8m1J3jdp0dKK2GL2YTZiNbz15sr9jqOJXZ57QAFD6b4YqyV65l85iGxav
4Zn/BTRlRtWvSAGRs7mfBnIn4hhTxBqIhDqye+mGKKzW4AeUwVOl8fS1TZ3cA9OO
7mBOY+SA/x67KsYLco2H9RGd8yS67SMsz2qzFhp7iRI08D9OMimjsd9//s53EoWv
l/lE1Ls+9fXk5GPC7TftJCnj/etVCsO9+3uJ993VD21YnM0fwb1ykhudtWMlT23B
qtUFwt8m4zlo1YZD7j2Plm9WPyPHqeXbeZ2XojiAcbpbHTDAoMWAXBRARLSAVIFz
xeu154ZNVK/liT3GaHVTudSdmWV88wE0DG2HZzppHufx1RlETmuTMLkD36i33fFL
K9OLJctTr7Oc5lVSbymyG+3yW1Ktmp/ziUi7gdBD9mwRTDXZA0Tf5b3RE5uvtbBq
0hl3zYja3NKuujx82Qmw9Mt5nDTXdJXla/77f5RJRKhhoY4ldy51R6T7dI5wGlUR
TPEZzsMyQy5TAJA1t+CGUZkn+gzEMAkbwDLoQ8Dw6LoA6FozDe7zbDSZTJ+C09ru
uCjKTabRnt/9JggnAB4Z+lHd+16dl+U3q2odiPQ9VPov+dyT7GkfgUpIMaZaNoLA
BaS+VTeD3VNRdZRcCWM7AsqFpQgxRtqqviOfp0LP8wjF7bsl+oVDAt54juOnsD3L
H0LAxUmjStx8et+ryvFOQFS8LsOPV9MsXkEhVLr6lPfiwzTodmmBO56TBA6CimI+
ONytwd+aRvKVKcOvi0vRt3tb7u11SWKpqCkG48PtlR51Z6uTnjXE6thqNjXOu4yg
RNwDssbDd9ox5lviJ37uLpg77QMArrBlkg/+aWrxpYi0O4iGZnVHHHfdJRyr2l/7
ohSU84kfe6KM1lvVAhNMh76g6B2pgg6VSl+868YtZ7ERHVAFQ26ymesTy+UoD7b2
BXOZNyP+xxSNpjQ/i4j94ZGC+ZBZP4Ti3l36MuhXukWY2cX9sApq0a49eewkrrRI
ohdU240JdENj//Tef0MIu3r1qzklipVWcWKVsh2y35QeYfKaDlFBeN55AgYpUzY1
N4J57LciGVQ9impAmyZOeh1dj9oqyRAzBgmTEuf2tSw7vzIlZVXuifgTgI7avv0j
mAX2ubJZl5SnwNvFLhshM3CSVldS6GOw2Ov8wHRNBBmg0NO5F97cEQlxXUA83Oyk
yJ5GKSsUp6tMUoPIyVbMkma56oMAfDuahbTgtGo7YJjFJ9uEVzXT4cvyuHmPej/u
RnZy0vVnjAVCGyTWSq6ZahMowhIYi7mh20tiNxf3BbzA6EMjHClZL7sewEj9KS/m
RHyDTMiJ6dms4mgTOYrVoLXsr7++t9iS5Wic1PGJRSsWTQHl8p2DWBNP6EOrM4QG
jOJm5Hs9jLrvViuQYX1Mr8yAbgz94InsLi2RLg01A954S7GBxPR68ELow17ayM6b
dI9vOh3AcN2dEezmVHVZ79cHs4wqlaHJlNrAH0OtqZEu6a0LyCdPDgcHSWu9ZbWb
aJxna7C5cdhBa4fEMC7B177dljfEoHZdBWd9tsm4IqMJ87uLWnM+7q2wX3MVyb3O
xu89NmszYJe6yXjihjT6IgILV6XzzbKSHI3cLhFfVPzJETjcTCSL+ogIYms4Mu4e
94MwX+KqEKhrr78+2L7ZktzqeLAAFV8Wr26wIGzzbXE01tu2gpnRl4CLPSJQCH6a
p93yeQfhEic9hNPOdjR1z30QXzmN8v6j8ZttGxPI3V1zV7e7n852/cRAU0sjqgg/
U1tSQZ9id0NRXPdsmuK2/RhqkSsY1Lx4ICzw1XCDl3YC8zUaRx10RYqstFiCNKIB
/+J42YKCJXIZRypTuWal2oKeaB8AFgRQ+7PC3DJwo0MB0FgVudoAY1TrjHEO16VJ
uYrdyqCpKqsx20x8+7a1QeeEtjdaFDwWbMvW0IkA1Bpt2QYqwkM4qfbs34z3MpBz
iMI2fv44jlO0M2V/JkY10G3WZ9gBgM4lubkm1YhgKvHKiErGbkxPfNiZzcuiGV+B
nHNoANR95kPAGkUl16mqilpxp8n/I/Vm0Suxa+Onjh0ig8mOW+H7wNzusc/dqZU8
VphpKk6OTm8w2npywGutLT5ww0EGmBrWBXPyLMsHPaX2rEeMiDKmUHkkhI3RzQVT
1EEZN9Isjg+DbhP6xmeDGsfmMOqdYS2N7qV9nLF7fk+7tboP2rXEcNdDwP/K8iwQ
CLwlhmiNDtblweUdvqXGfdTr/Bi7xTb+GsfwE0zbrBVMNAhCneXxogb7MQD+wfJP
3ILtM182Um5g4fHqf1b2E0xSgJDg8K8kBzvkel41pIZumeU1gSBb1mFfoKtrnzov
mz8ALKiAsIuxEZpLCkrQ3Xjnlc2uylgIVaBZiJZ0qiRwjXO2fhAVAIv0tpKbl5Yo
4XlUntTtZjTYa23d8xulm/o6zcjCjEdvp/HGYgLt5cFpDu2dQkzxn/eAGwqf8I24
FOOZaQT0ZmaJSwSql4dpHiAk5Z/+OaMpirH9XqVME+GfH7ZqmgsNW4F0ruPlCpbQ
qLyjfaaAZcRPgMjgipEx33VbdAcpcOyKRowo+32c1NRWOfd7PzidLf6a9+l78fEp
pYB59sKLCRSopL0TgEx6jfkZ057gSdD0y95p5lkvDMcvykKYtUNcfLOtfaJFTPvP
gTxgDRNywLN6HwHY8OavmUkZ6GEpbtlTkxMrtkaXmpKSQ2U/X4TOzo1txOqFMXcX
9XnvoMDbSiKPuHef1XGGOzBBozg5e7y3rM5rcc8CmHvrfkfBRLtvPp8+hHgZpthB
zp66liJ1bBKFk4t23sZK7d1Q0gq/hXOdwKgCvEn+wvQ79Tpe5JwHQu0ux2T8jSPQ
G/6yeLM5YndLNuN1Im3nUPJ1sAXRkgrv2QskR1o6Z7BR5/R7Iogtk3G3BiZkc11x
/zudWU0Wlvl343R/ybzZQcM3VxvKdwGPNFgpLHtwpuvcLg/E4ozNpxI0iKJiRM/g
58OZo++YTLea3oeTINrumTvaN7yMW1MCzWX/lG5XWgiL6byGDRZgMzTsAm1IH0tn
Ele2fqobTI0pwzpp2r1E21pZFYPOkv4SG9ZZYrLyguEBWMBazL9DCgtFMvU4c4LZ
E0ZrlmTC61HeXtYnKA1rJfCZIdU8yEv1qZHOdGLFSSMHDvLUuZvNr58oWmYe0Mic
mxjMcKzZtxpSZK9hX8yM+I1s+hfRdnuubqK29IyTB3pSrHlikqRQ0aoPItySHzXg
N+gp+naF+Td2L+/7ggXXOr/NgEhHFmTGlwMvyUSUKEUVOdNfNOZVoMSzJisaGAIq
yGusZdfZG58xBL6zYWi/CH2mEYHh481wS3XLb1keERQjbT7EQlB+UkbIyp6DXUx+
dca+g4GeaG8Kf31Vznk3oUv2sCAhy1dpZwpyPYS104l5tyOOexRnlr6lCmgoKkZP
rBUDUJSWUwTT+0dUcbMJc0MiX70I2qLJXd0xjN82niYqw2YCnG4iWyl0qq5o5tQS
dpx+4cRvtm2r0gtafauFfNNJRXcFCUObg8NnLEXY1yfDbKonpkNQaMx4ANMUIRCb
yrS3AdHt8bvwKNkXriIM6R+rUekDzxflo1kXstBqHfQgj95EAXf8CWSVTrHvVrXt
CjO+kK+o19CCRio89KLsN+t6VboqPW4gv0Dk8Q9J0saGWN9WmIvsJhqV7BbT2iEy
bKr761ZzBjga0wtaD39g22oXu8BuWERSVWAXRdv4bgHIWo6+SPpzE/BX12kSowoN
kTXkUMhe4B345sohXMaF8o5QX0zNlgQAWQp2TFTv1x5UCCtItbc9iL2X1Kfz+qea
xTIVDa4gTI5RRjGQY2tHq93rgAznwr8Z5OvDPug/ZMOsgqrSZY+FDAUl5EAJMr66
noeTSWVF4erQSYhpk2CzzIt78m3BJTDuRnX/VeZUljOPKWpcZ1lvgpJHSz0gCb78
3971goMkimEYr09uHpKxLHG0X/nf9vf6KMtfatq7upmYaJZhig209KlwV7VW6DhI
9ODx/B+OIg3sZ48ne9tngtcLvh4GXYT6KCjOFrl3Pbpo65JcELFozBR/lSiMNA4l
IXUKMNs37sJmceOFU0s6VsPSjKCTWvzjLwbtpcyzKbx+uYIiWdcaUpWY1Tiv8Zyy
zlfC+leXY2KEgSDTSoj3fbfuKKSWxX31cFXwQporgr5YMVTsLWMdbUurVqe2bx3K
iqRq1NcOUY+wa5X+yVf5jYGFEeWLw2u9m/ywFr3b0szHjomR6CEvInsU6mxJA/km
2XZSN56MyZLIbWGEUyZsyN/t0f5BaiglfIIwj15tnHEGv7x9v/6kjGOXBkUHTfu+
kokqt2PN7oAX1T66+ByJYsN2EXLEQbot+z22HwZu9EzE8ibcGZ0ZCqrZbROZMRwa
G4J4epxrSX/EfcjjjJhPhSmkdMGA9YsGVigEM72o7wly26+Q2Gf5zxBw27AV7Gfq
AygCxPwzeeAPG1CB/bZblEL8MdhDs4t+tsXMoE85AQ0Sf0yHR7397Vk2I532n003
wO0P6+EBzepDukgbkrhu+xCioDa+axQn5K45aL54EPjnUWFPWa1t1/0V22k2aRrw
BvPBKdK/0h31SIJBYkWibmKmuBDzByAceRzatyJerljxMkPRfVO9/j9U1ao8Pbdw
TMI7VDmnVg+drpT4MabSTM+RKPtofTwgvCWASBvJo2ePH57USR3PJ9hzViRC9sha
uS3aY3cafx/TjONsIRwWmRyXss5kIn4ajXRkt3AAUYiYlh9Y5cf7OjlCre+cKNDM
GCduNfZD2AMN88ljeTITBz8fTdqxFtBPhYnfEDmAOXRv6nmQZgX81c/QKGM6tW5G
AiovYE5RKD2Erva3XVRiiPu1Vs/CNjdEDDuLQQlBt+Wec3wwefO8OAwbyrzW2Ti1
tq0JVUIOHmg2ZqtZcl7+3wRILnAsbc1rDkHRKrDPrC1dXyhWMhX1mHp6FGPohPWg
hOniMBV5Ry5la+HYS6DTPA47nf2xPPyXvD90hRWhz9qlWSK1RNpcHtHuuI8qcx9g
QP1ai23/PqfYxmJL/4SNvyaFAy4QhO838gDRu/4W7zYLcqt0QVWjy9j15miPD09O
a9f/oxoEtcbU9by8kdZjBk3PxxywEgmLnb0+YLlpKkOTVoSXixQryEULslpqsEI7
F2c/nGVjzA5GmvdK+offSs6vsliqL++UA3ajHWIV3Vkhk2b72h7RFOZewFsLqWrh
xlo7Tj+dIJsp1EDGyfp8o4lsOfJhtRMTFldNoiKh8b+mMuOxx7+kZhhx433aSvaT
orz7HAJrhu9I1NaXOPLinlG1JNjFSmU76cPBXC/naHiOayK4mT++BKm6K52Y72hM
8USXkXK0si9maPnpSxTlLhQ81CVXDR2yhHpB5TntQ1ixTZ/pspjOfFLWKVsw1/mD
xbH6PT/ww1LwZ01uQW6PjY4cbFoqjxI+SpzW218o2BHpfQWrcoDRrCVMdlBWB+Kq
AVtXfel5Uo0Ma8ZhDoVXF5a1LbdzYVp30AsvIKcfdXt9clk1TMovwTf3cpnL9Okd
j85Jc73yCXfydljqPx9U9WZioDkfhD2hDP9oO+JzaS5aMEaMJGbvaNXBwCMfcCbM
yRYA1xERU80eqPlEi1rKV6y5OAkpuTkvASvLtcYIxgFZFjW2387Aku2ajTpowICJ
wkWz90k6V9XKrkBY1a9f5bVR1kdaenGrqjE62Vjp/fq8VMEXEShaBtMZJenO7w9c
5ilkUq0WhYdqR+1jOFYO/IW/cNUw4LKqyRyvf7tjI8vLaDvxl/GURVgj4SeFX3nH
3DExkd9bDUHuJ97Z6c9EHek8CEMn7ApDwedeDnKb931ktuRHLa/wXJPNBi8/69eM
2VQT5laPVQ/xgxl6JOKaRqhmguJQTZMsl9EQVZzEMJpE3n2JnA+t6MNYGE+7hEQ0
aeCbovFfrYEzZzjmFnLUNRMUGyMx580w/lBW0iz5rLgQVC1hqhd654xvBZ1LRh9b
zF6VqARL0/RDXXMXluA7lDcYysNDd7AgHGuPXKUyY67o0SY3/XkG36zhOAvdeM/i
Pf7xeP8VMHz0AbjAzRCEC0UJd2gcaa0wh5x8K37y30nij0Jr1m3YkWBz53MKUvB/
y6tFWcuB3mJIe/dByCzgNJPkNJTOVFiva0AG/sCJLY2wEZju/yk1DcYOiZgZLLfK
ispDZkWgBC7y2S0VCKQuh0foi4HO6FZ+E526OV5QIu3Pbssod82Z6Qn3mkYvmveM
scNnVLHOHd/xJy43NO18BTWwCMJldOkjOE/yo2sG1JS+S480BE4Qad6p3N3LL2nV
hAbLZXXz836cK4NC79Yr1Sses/XDkHAyPYn9+umSNt2aNx1LjP8lmFbh3fpEaWBy
pQOBEh5YqIt/yy1Kc0/kDLQma//8gmqlgIv3o5HeJjlX+7V84+ZRU8sY9IH4qSnW
2vK/WYysrkvT9MX5m3xEBZ1NrBkzfQP/XnE3lNbWITmrl8EAijJ9+2+eTrEll4X2
PMf9Tv6T5jj9i+TItm53+J0upK9N3JSVuXQl/ciiR68Ms3gTwhNpy1gsIjmn9Ljg
gQZYZrGlszC+RAoANdloydjDImBWkPjIiD9LwqJAMh8+5JAhlHuPoVBmcZdJtXtD
QmpINexQk/lvCbqtrjjDUbIrqcT2oKNL6R6QNGv9NmTHrN28Yl3GDIxE/mYlvzat
UmZ8+bE294p8P/+2raZdkc/AMy2qWzGwITErkaTRW//MWqJK0L6znFmvxfEgiSQM
oa1cU5j7rEcW7FW35R7ApiQ1BHQk/wDvu595+KQtzECoe/6poLP2aHLfKwsVh8YY
zWP8MA/qZhEBadQ9L8V+wnOCl48h+TwxPJ3QouIMi1+VM7du+CWtNXlxXgCLJxls
9Dg7H/FWj5isbjeME0BmSAyjOtWup4elM4xVyb1Q7g2fABBzTa8gstEccabVgB5N
KfreND7GuZSDY68vuDfdo580AkDqZchOaNCqwetfdjK6bBnirwOKH1NEX55UHZpu
W3RIT1YothN1fheMHTltMWXHnxbgfPGWKa7Am1pmk3kwgW0haF8etYaw210O2eJo
EQ3+M5SwEMAeF855HVQY8gRJ1odloGmR8q6OB9xGQAB+DE2dJM4bEUWiin0BKA+M
xt8ZiWqPE6FfONGyIPof1GNHtlvloS9atzFQR/Z3nFnDiGP0DTSRvpSHtQLzOF8u
mZwfZBsFYmwinDFsqKy2kuVHgLmdx4Y54LJphNeMtM43S1x4VVVxXYYYwVshoW4r
V+cPtakB1htwa/vNmU2hCSEugtUbpPKK1l+KXaVNKrmdTFva8DjOn9UQT+4eYbTl
jQzZihW9qFiYnoeOoaMn1+QJDbO9RBzVDZ2h5CkIZhcYS6Qs8RCJjzzY+3mnzqNF
kzCv+1s6Z5UKIRmnF5OUmKA88qnIejqKuZm6+ANbMsWyeB4k5iVWtvDwaS9N4x3N
gw9UDSBsNuNps44MNAsk/VcI2rjjqcWU7/reMTqMayY6l6mHCoET30ow2O9jGCA5
eyht28pKK8NpTiajPGLjkQtgAtdcpoKhusGCSmvTU7pzViYndqddfsA38JcG5RDv
bdwwiltNqH/rZrRwIOBkvzfv3igHqnxcNXNSqCvt6TxXI//Jh0Y4x/+RWHayW7SL
cFggabKsRfuuxm/OQa9dj4uMoXrAY8UNuzXxUKLjgZGLD3RRqDy4j+UhHaH8eE5Z
plQTs4uOX2HVI/xPgbiUl717Ctio74dmsFiC/cWU1QEVl6Jo2nhDzQD6axOvt2ZF
bAnjx9ew6oCPSMIfssLadPAwi2SDagj4Fj+NN9XNy75CuvX+jKHM0Ji46wB5+Gjh
yJrDHkH44xIty08isoifd6ecvqw5ajwyaY4C9TroQ1w9Dg2dfhdwgUR5JQ0ZHOPc
SmfEAgSqdu+Yn9J0nbZxYXplP0shdjJsH4YdcLVdQI6v7t9e8hj1hOkKqlz9joBR
20JZQlZ+4P/wRJHbcNCw+zsPw/UDAARk8okFzHK3ls4wvSaXc1XHLVk1dJJhTcds
6WyoSZTJR7YcUPc+Qqq6ISfhq2MYgBZJPEu6HTHRy+fcPnM56PAkaZYDI9bI1Bui
8Ws35NbuT/ModlraU2O0IDVyOPh95O7EN64cqcOA6T1g2bnI7CraQ9WrhI+gzkBh
ahPYq6mEAd1Gce0CgUgo6lZA0U889nHhZ/ojK95HFOcac3hoj/R5O/IZQPy1qGQH
kC7KBCbCdfwbfHZ9sDSX5oGD4Fps6ENRtEozaLk7iqJ/RksGqW6a2a0bFDEFHZR6
xQdskrXXanh6VT1YqbPVQMVdsnnxuSGJfBl3hfUniGkM1P/mWd4aTwlFNizhcktt
g4+DakkuY+/jCwaztWX45yLAjdRauukpiuHcfU9BI7CHdnU73glUYbFKrk84+QXR
B/CptD69oBFdV/yn7iatnskj7nI/ha0KPhyn0Boay5qjtw1ceg2HZhuhT7Ou97E9
3DWL54R5TGdF6sXxTvTe2QOUniBsRNEyIWyvZODPbaO0/gtvaZi6bJZqeGAyYrpY
UmA0sUw9oJg46TzecU1DHIMEddB07zWITJWnfN7yGoEw6s16qkA+cz2D8d3cBwF7
xZ7IlVOd1rWduWbk6Gv7c7TChEfYlOlK89we7pVu8XrJt58w2syXj5TlY3re+JKe
VdXbupJqcon67CPPoaICxdpQfIHOk5sugKhIj7OO644yDuAa9LI0Zb0ykEngPhZl
Gb/PPKSI12WGCdNNz9rJgSf7i4GRyUHcsDYjJBuxxbQSOP/LFGhodObipgi5eZLy
jC/IFJOLjaSg4Ih55cUomBVfaNSbsUHJaYTnDkTHZAkow3MkoIyzI1Hv+xUy1qn7
mDS1CHxM31ar2UXuHu7OR0i8bMbUR0cPa4NgnlFLGpiOyKYEGfEymDh/hO4HiUCW
5JeS3o4U+I7PI60b9mYOkZvNP5igr9yqCNe/Lr+uyTAt00eCsNRdJIPo1WJg2bah
JuFKjfnJ7LP6EJKDIbRtX5afsrWUCRptf6Ivk3qKp9aTg6avL3qdFAoVarH33tZv
1+EHDxhv4gi5eCkW3cODDUxDHZsN8xG151s66bPrfdI0aeNVdqFvuX7Wtl0hilkR
WabpgSBvq1RWpIKReH1wb0rk85eMG/kYYnlbrpcduT9SI26GTXNUBiTz0m5kUt1O
YcQApwDB7fL5aFkCJ8Dwn0jaQH6Yo04jpTpQm+eN40vpqaoikqjO0JhfpanFwSyA
7yw6Z1devlu6ArS+UQEMNHC9SOfELIlw0BsxX8HZmf+U/r2aOK63fiMZRra8p06t
V7+Nbu/EkxULnThtfhj7Xdy4TxNyCXW/1Wf87qYxxp0GHRCHoXrRAvhDLFqqVxKb
PcHQmlhYnwB7HhVpEJtb0PXtU/VGQWBzjaQbjh/opzure82oXjfEn1DKs4RitWiC
/zGsw6fiyXJ1V4aivjxS2WSL87sM822JutTmrhu6I/v5c70CBqd5Z/3Aamn9aBIV
iGTULF3/FqYofTPGdPDFSpbqM0uOPYyweo+hCCWjU6f9xKnrQJjoqAHG2DuTazbO
77cM+ShpwQmPeaWLexaEAia3TZnP3oVwh/wPL7rya2PFy7aX41K3KlvrKxLyw91l
9igY0gRM0VH5rSfWpFwLO2Bn/FNpyaLvqaKjLt9Yq/i137CDeGAgAdcTpsT33l1r
K4Q5trCeVsyOi75DlkGhQgkoeQmBckSUA5CXaerNTq1HrFcpG/9TYSmohCij3U/U
ncKJS79de9whTUrvzo3HrPlKLXB/b9v4vjEZC+k6irVgBTLDtMMPmZXXO0WQimSd
A6i6CH93qyC84qeIJeLfhj+HlVY9yyIIoJEmRVRJ1AmW34dbGY3w6WcFgqF//EU/
RVsLGRBweH5wXdAJkJtb6WAF8jCRbf50tBH6CJRQygthNtZEopT4WULFZ4DXcQxA
RtX1sBT1ihGxTOJ77jQlup/gGdgK7eHHu331+k0ivZtmE6Zky8m6+kZ85J33jCtr
Oy1wu4R7VGHXGqgjdIYkAsVuv+H76d2CZCbU6cAqMd/RjgGP2KD9SJcgBk4UTxZ2
252qhEHi+wxUWtR5tIHT8k3gKLtx/idaTkGHt7BZx1Ndpc/JxD6VJj9VQO8/LOJS
KcNbTUnPtBEPHVUko3EF98l1S82zbr+b/lDCR8b9t2Q00UYsCGQM8p+4QXUcuNpd
XrvA9hnt5goRDnuzrkOWGgoLQSDoDj7HJ37aKWgl16LvdFfcnTC41jEmSgAiLULz
R7mjUh3tzPH/dt3rwy3jUHLwKCoYT4zK3HFhfgexKwTdnZxeCaUM9pzMnrXT8hCg
TVQ0O9egZ9zLtL6r0RUC6XFEJ2FQjb+KxYIhT/e1PTVslqG24opJhbsiS0KV1RPG
hjRtgCXlPJjz2vf1nDS3Nd2fBPehtGuNnWTc1AXQlHvLq4eCdUY2bmFoub2vXfdn
QSr0r84rQBHezyF5clUVoIlrXGgSKU/fsQJrF0Ge09aSeSGKQzw7xSDzHtNqM7jE
iFPkCo90NpVSU9P34KG467AvaaBw+P4GiXhk/ADh5lcKOCPylBNgSw4deldyjwIR
1HIKXSHUr4t+4zgWataCdHqpnlTrS6LX6eHQDcGJRX0xFWB8w/6n0Pg8RnfP9mZA
Cxb1aLEs/ZDxbTCW19qkVAHfsO3pZeX/SRHEw0nhM92N4V18W8VyggwMH1t5l/Wc
5gZdx3kewlfWsErYYwQ7TKEFTG/Im+3GLkwpJ3DWuEb63aC+L1+cSY7vw48WJv2P
HuFaArYd56Pm/FJmEJJR4Yp5oNXCg1eKvOUsrkvC+IL5vvWYqhJMtT+FJaBhtT/H
M6p6N2U2ocT9szLBeHCuX1kuOLBFjGwQexvYYg8WgIZEZ4OPkb0Ajvr9bhDLOjJV
c7BU/WZ6aUdEVnxNxjvBFMhjAMtKWMm8vuaefgEcUsraNj9WR6oVWx8HgZ/0YnFt
e7g8SC/7YkETyjAiF9UWvBchlaewkgqbGChOZhFN+sBUqq8lyfFqY1Og3mlJU9Nj
ggSSKl2N1APMIWu3PMPIgxUhUCy+acuHMA5LozmqqgH5f34AtfvPzCGeUI8EmFkW
GlC3GeAsskr9Br15aDdkbkhjHvgRNU4FnPaMhzvpv8hNutGGi0WXQPcfynS7KcBF
ECErOBsh6N6I3+5CkxjnwfmHP5zPhyNjJeSoAQzhi1akbkM3IjGBwhdN6p065QU4
DdA9WHIFh6jOyGWRKdnBjW5pcD95HLPCvAUYzyHzgaC9jaf9UcnfcDh46nXtVIFM
3woFSdJUB5JrVXIBM0EDEgO5NPYgRDy2NM/qgo7Du/4po2MRLbZvr8mQCknT5lPQ
NroQC8K3RmRYFU2cxzR8bp0N0e6nSedaKs+m64lPcLqk+JjM8ULPqxgrr6HuOf2k
JGqm+mIBDwnTtYJlIqSxkzmhvIfLnIazEfSp8woevzLG7PrbXD28ptunzUpw7hRM
6S/8LuXgDjYRpe+ceH5vVkJFRb2svRen7AiahqckpLMI43hEs0qTNi9A7J66jaIk
CwQeUcYgGm4OZqflRTq/OkAqfbJcJYf2ostlvn6rmF2aYmzS2QmPbOlUat0l9Fzm
Q6nq/GmUzxLR2855twakLTBkCxs6ckpq/kplig6/A2aHPK3jQt6+31aFxlDUfrp4
4elQR8CiNzLUJL/zk54vhiBqZGlcqxQzqc9brdg36dLczO2MIJjjMnozZUVpUxiG
E4ZNKbbl4yJkxAD8YVOjFqPYP0DO/SKfcsnj/wDgX9HCt0Swjorr9I1ncpus0HNZ
XNsoKFZORSFd6wzjR1uhUZw00+NzFDP9DrRIA1TtU61ftMdc99pWhR0vv1/b51hu
LmZAAtUWszsGHQmGdl3Zv/V/zj0yZTIVCcUxoXQQObRWC6BOR6vixo6HldaHXHiQ
Cq7gGgjie2Ri3ckBvB2gl/vQto6ZoDe8AQaN9KCUEfTH/5nVoY7am/+aif2gllk/
8hWB/disseJQrqvCgtImYy1rcyDn8BRVle49gh6FrMG32kaOUDmkNoj88ebMQkF4
QnkdBJkAPgPSktSvyBsrNDY6R72eP1KsCLFH4asvDZuhGOPatbVGS8ZUOBYUfGBC
x8unr+2WpSzedd7vKqwgTZajrgmZmjeKcTDn9pi4XTnd0m5niAhTYJSriSjbFjJu
ezcwzTnFAyA+ZURe5N0NgCWWmEjOQczWEqXw/OqpFPEDgJubr22qtJt0eoF5fGN8
UAVs262qHcalR+RMylE3IXrglRsIIzUP9pi/0L83r9nth0mRVJQHIQ4VJbTlJYSU
8NSmw4X8C6AIXm+eYFTmuV7WyDkZomkGNrRMD7uwsNG72Jw0dv9m7rQ3AkWo+Z34
ZaECCHnu2IGOZZECQCriZsgl/0aYr5cYRrmDREjVwrWTKfijAyszgG0PKIYmJfn7
vFGUYRkGt1nW41Gba4Jr5Hq5DKmBme0/PAtZCl2+o0MuXWBhQQJB7SOwx6uHGZUJ
HIStLR6ueD1Kk9Tuz0iRHq6JZ72tCKcxaKi8utBtKPeIbJp7B1+bu+e8Ox6NAJgV
Tnm0TopOf6Vihta0ko7eZladuDIH70J71XVrdvH403VBKMPe7NQV67jnVknojK+4
2HdICmntjRM5Ehu2dRiqekP3994xAFPiOWZ5VXF4Ez9iaLmIRaNuub6ewuAp9+oz
2ZdZq9Qi7hu1ryLWgJBtbY8d74DRxDn55apDjcUemDhvkj1MzsaDV1ye9sJyWsbL
PRe2J7gJeegL6WXwyHYJ3C5SD7zeoyDpwd+SnMvTwo6GHAPIBFAsD+H6j+CkeXau
a8ybEO597+nsLcayWqbQIXx29WeSmW+6m1pkP8fmcE2BU/jBNxHrp6d7ZZl2LEXl
5SKDQSaISSg3brS/0+EgNpQjTcv7IM9OEHfKPtbMM1KHEEMOxQzzJpn4DKKh8ntY
TgEMXjqAfzed7ZxRCZo2jVm9upfg7pIeLbbawsLr2vyn0dIbeVC7cLAGpyick4ym
/tdYS1xnUtqUvK+yHLsm8XHeJCNWHKVUxtdtFXlqd42HVHdktJws5C9xHXhmW/cJ
1MU+cFTDIO1EHuV8Et6+VkXDCXfXt2noAtSm8cI97IcQMagZE7TP70Pq0W26ieCp
09QKNZ03XE1yGnm237F5OqJ4C0rddoRXFbxuTQsmvTvq0OP1xPJgMGtYw3ktZeFm
ufRKBbwFDTSEyitmJlatZjfKlsVFotttGxflQ1qNOevDMGcr9ftKlkaLChKSvsaI
uhPHlhTLXXJJ9AIEDdA5IFRygNqDLpTvfTkanVXRThJS7NDBSH+i3UFQibJE/yw1
fKN+MItHHVTEOoVqpZ0DPW/OmH//rUTT/9PgF/xvXUcpN7AGAl05WpIiGu/Rwzi1
Txjb09l+4Ebixo6mHLoc8ZOcnPQAOpKmcbyoMqoskrhll4U+NCOOCPKSxPmRGFX4
ExtpWoTnZ1ZqI2mGuwqzaWZKv7FDiNyrrjAap7X5q6IegIxYUeyOyl4I/2P8aEax
VvB6xjpONKb0SQCcjZg35BBmREy7W3SoaEG8O7eJiuppncI1QvdYLlNBc9UcdnYw
yH/6JgAtqZeinuiKeOz/GY1XHzRkGF0JhV5tfCY6yCLEhiu0k79k0s2OqJJR8zMq
HXQWlxf2iUDFcr2nC/u+w62WYGMX06YGcgkCOVbiCKq8fnqnYbu99MUiELPwzLog
7OQlvA5eraLqry3F7Bj6FdVpoLaYsBp50drYS94KCUaRKGkOhKWJkQT+wyKthh9r
INrWJKl28WJBGBv1Rd4og3CfbRUoFxW2SbZ7eUsEqbxptEYBfrgvIuX90HqTixF6
ZpENoaCRJHzbnGEGSeYi6mh9iPWZllzetekWYsNVCsm6jTkXwtUcURvGeWQc+z7J
YJW761N3nem0+pXwsd/mabyBNqkoRvVVpsuI3cM8yyS+rYq+BuDoVL2UC+ciX8u0
MgimEsscT7ZhB4maUr1FxI3zw2+cb0qeWHOXCRt5jDvgRH1X1lUs7wGfaVhEP4+z
Xc4J2fkxITDpg6sWr5ZaSVV4oZ/BQfFlbjq1OYy8o3kg/0db/66K8X0URqai9ZqW
OHNReMvGQGoIf/jf+Xcwp4wBmrB67R0zTldnr1Elwa7ijdmOrB2ukrZ0O3CAyqGn
CZfrbRRmwkTaXWK02OEbliPFFfFPBg4HgUQpPUNfcO668k8sWIv1I4xqx2EogDO8
c/TAta+r0kV7KKOwaVCHJVUq2iV2C1DrQuvM0JqVBVMoIQt6ek7iY3U7Llr7Z+Xt
ERwkZb0zhmAM2nnz/8Z8XxUXLfkwGPp0XqPuUGc6HxA+Pk3ZfyaVFTcvjuvKqf4w
LOOo+4DBE6kDxbTQQj7z3h56nYiRERGVmG4udwVVZmX9cbOGbHjI0pdeSWDwclFa
4KJ4ve15ExhnlJY8L/Wmb+Ad2G4oPFV9pKWEeN59JVpoC2FwiuVzfLASB2dC79FO
ywjJr1jKdsRAPyL/lw7R87uX7T0LEUgwrDztdVHCQceeylIbrLVyPYhATcQfHtQa
2QIqjX5tj5GbcsIJonekrmZqpbzwIjj98EilpqTrq8kckDGIzrCl4K85djTRL2P+
QvB3NWxe+xV/qZwCDiPK20V8omDyn6ZzYwNWtgvoCYjM2hd4Q9zmI3uhkkwuJe3o
C8EUMBNmv1PiA7qsDuWD+P2R1f04Ry6TdS1Lx6brD0KBPjoLpeBQhvpg2I0zJPOw
t3NInDWpdI3B+DPvOzGgEtbLprhNlWjo1LS+2IolzgozQKSS2qgsNK0OE3+CMBsW
S1XE3+BbhC8+ShLEPBh7aULzK1EUECVVXJUb1m1Dvtuwskye/hSG+vKRg10kzTzn
hVoWonWjjrgrSrR0OpSkL77ssfuBDCdqUfRQ4p1eWqTAawus58rMbiMrrQ5aegEQ
sl8+lrLP7poUvRWfF0zlTo9Z/IX1EFFxuTgX+L9YungTTdYprMFkSlyCuLv6scBY
X/3B/q63ghDFXjKgEmdfHR5DFmyKPKRN8fBr9t9Hk6seVNA+m1bmQP+NgwUMPSXF
gPMGpdLSUlIten7toRA9qa0E8SRw6PVJeAHjCUWn8uGn5Br14/hxLrJGdIeK1lwl
xbbvrYth1V3OKE/GG/tttNnnHEJ6SlVpt4DVdR0yqUGJQiVzPqFMWsq/yBvh5gfM
8HDQW4DdfoxM1fkRbV2jVvxqG2TCKTXfZC7+H0dFQ0sLYwQAiyV19pUX+vV3yDkE
LU1dVzkRr4AbPaRlDlGb7WrpveZ+fWjBrz0W8RPraPDxy4Gtxg6K41sq+IWkZP/I
WSq1mBXh6QKpx+RzQNNTvSQ6CFtujLOTkT+pTwYI14IwpTsXKn7RTjy4ST7zETXV
0P473ZJwI6sRm0FdLgXwOC2tZceyhtO/L1Lz01gCMRwnp97cRAa9E2eUZqN8u9D0
QTFVvs/9GvRp3n5uVVvPDsP9iiVyNGm74Ak3kPJ+6sRcLR45JKUpqQDG+K2mba6f
pq89l4/wtxX9XU+6Vpi6yQxna/n2mrUxPINXT1Q0TCQW12Jm89b/dweO94zlo1tK
+H6h718giES+HiDL/icQnFEf98ALX4AqgYi3qYx++hTux07lxD4pmPURdKEn4IE6
b+njX2V+YJBa0SsuijE7ZjiT5sXKZ8iNRG1cmAzeeVRyV5vq5cfX36YQ3DCCir6M
2wvDHzPcQu2x04LBKg4wa6F+RuPCNF5jx5yB55ErEDZ3iDfrA2i7mlJ27YdA9klk
+dmbieG9hYJok3K4cwCv7kXhzifITqSaOBqrWv87c3L/hdiXMtf5TdzJ6UyeJpOy
YrL06GrR2me5I3AOXzYEQ34VvfEA4R7nfdai+Bf7ctz7O0djElJPbtRvpubEZUOL
rlImyBHuQPwZBmcJA24oXCRcZNjFHAOhLJXiBeT1cEacFnZ5ORfiLuMlvvM+eVet
TLGrMbjM8FXxwyoEoQhaz96ZSN62ltzKBIclKPFps7/wq69QcZyrpHvxMGdwrnqn
/5ijgCEEeNA7/3RYBg3IWdmU8D5UCB7dDKYjTzcvZSGRdvyzZLR1lX6xjRGEX3a5
G94jlmXPw4CgfdTMcYzQVhbbwtDb15dNqfc3pSdDAX22/iPdHaSkhfHlOWlJJfG1
H8hmydp8tKty24Abg30ikowIcxAaqVtGqHKAD8p/AkA133yOWXnMfrEcvwKLDK09
2HWWMl20Onoau/QbjITM+lzAPD6yd4RjTjan70iZM2iP2UTcUUb3GXRGzvVNyWFD
RVfu6X2z0PNORkVzKd+59vO56am19BAHewtbD5ABSpnAlIkQtdUMUSGOIQTDtZ92
IDP1K8J1Gr93r1KPtpErEjdVFVYRGlXuYNqPMDjjUaRpdp4FVcU2eispGxIfvT+S
rsmVBKApRi5WxO+o5+OgEFoemjQRpyj3i6I4c1FMAO5cikrLjdxA/0q+u0qjP81E
yERaPVV6OcTe5UUMYlVlDRhsXwxF3Ebp3uJY2SSMY17XSYQtjK+3qNd5Bi5quZdh
a09T4pHTO3gi730F8QY2Uwk6Kqv4JIJuUrAuufcGVlcg3yJYI4kZ/As+Oxz0NNPR
kWWIKzOvmT+s+nnSxwIulm2swBZKpv/8YuGuWFm70PrTsmD158oT7we/Ff5DU4i9
74GHn7BNt3tel/plGaA+w8AVaq2ZEUYADW186aAkkr95vJAAKBc7h4RQlTfZTtKH
lQ2bwOWZ9S8O2eRkWEx7ayXpv934DOf1ShHARZwvKSS0tnQGLXDDEIc4n6EG0xa+
XkZAmPr0flsmUbee+G41+qKSVRYHpwvSo/bgA4g0JHuCDNpIV8ZRDvytcIVd2sZX
dOhJ64Zp9OeCs/BS8eyQjriOiBr87y4B1FShDP0Wn5VXyc7UO+NKBKfgwiReiFYb
VOUrwJWGNCg0IvGJng+okisC8CMFSWNvD7cV+5mtZohm1665JYqJtY/D6LqZwqZZ
m8dlnDp0T8HW1XHs0BrWXREl08k5nk/wDnXueRMvrrltVjkhhqc4Ubd8Qn5TKAA9
6fp3G/dHA9JW/XC6cJZ0vTsevexg1m4sFVynFzA+Fkl1d6P4R0VmP3t+iZt2ZYst
DXW6WdQA2G3eIDqLtMQSv1WKB4Y0cIoCAQw8uVoCycwagUEUm2c+Jn+QDjPanN/B
7xu8klfsUKUAeHrqcscNgBla4S0mldGvfAXIhY3Lt0CI2OasB9pdxG8a0uUdWfH+
RwNB28mnDERq6cZGaT3JUNvdM3UxK7vlYPj4SRe7Bd26TJWZVpZ4TQQLwGhzo/yW
7VeCcHs2XZJ5bb53/MuaJL4sFsju3LM+c+6HRbsup0X6mNMonkr/MRX9Q0bvoxcn
PQnqmnoitXXuwSgJU5lsNCCP0DFTD8G0jpT/BrqVAgCrFkpuVCspqWUWEjPNrkNV
ti/lI8teJz2bow+LLn0ztQxHuFI2akpKN3IpgAOLcdtpXVB4eYEtLSyoK45kHeEi
Kbu55YNGJumdTzVhYiV8rxNGCsRWnvoPjn5lFsOh+96qw4AQpZajXvdrBeUwXKwZ
DWGuJIsGlJD0v9GOUjVXaO0xdFtWMxzvuq3Pfb2WBDpR6MWCq948pm5e0uMd8LTs
UkXQ/Z5yWBmMGgVmxlcTkIQaGlETODO4p24lpczFsFj/Tn1lO03YMvAX5Umfm4Se
zjtpxmwRVzKjwMv6geos9AVGt7tpOGLW8rcSF1nUIY546u3XlM+zIANKzeS+pMFP
AREA4u+hGRyuWTglhXghPbTo4Qkv4UDMo10wHxljJq9hjYEAvltVuKgmTf1C88vQ
X4oMX7WRdcH3pEFl5SyBwvp/vTiv+itptEgmtt11YlRAJBTJjTAwSR8KMYPaSoAu
EsPDPkYc1C/IKKpbUQ8vdEL2WUxCqKzgA7CkZzSto0DdHWixG1twFWgGF7iweXZP
t4eQp9YxnxPJOcagiMV8dVY+ZSyUMA/VZK5NRaL3fAIENNTVtspe2ONg6BwEzKZs
5oqhHP8ehKnOBqOAL3bb1B9l3B4oFtuSOcYVWUYOtADN+y9G1R/zh3WB5oOBgIjq
+cLYSNE/Mw6xJhvPZK10IcnFOW0Bwp3/LU/skqXDhsObBNR1kMfms+1HUKCqCyOT
ABEDP+X30JJl0DiC69Gw1j8LUXO/KSHmrtrehwrz9G9PK581hFjJQl7ZNcYd9YuK
tX8Rxb5z6QYDZt+DBg1xVJn75BeS2GJMBfRIhnEfhd+BwwFAAqbWhwzG/oGTeMlO
ZKneX2ATcMNwjSIbPzXx0zJr9dtumXsv6LMDlQgagL1LwG4jsuIL6H4P9Zc0H7v3
Im/T0Rl5bj7DpHAOkljizqGY7k2NJfCbYQqv0/o2JMtfCmz1YSEjFK2WZXWc4+SQ
QsTJ4Lo17JgL/jNdIgk2R2kRzIcYnNdHZIfnlgK+8m4nL9xAvyV+VCVNuDsVYTOA
x07jEsX2NOFEMcBr2BkEVejEuPO1b1dPGKM9E/8djXac8sGm4GHiIH7YbufAhaPs
snpo35jsVZM+aZCCcwoWjwk6O0c2isfRY43wQqkdmVVTyRVcM4LDVh4TgzI004Jh
MZS0oQ40mqnl/51wlzmIKQQ2l5uJeA2xL/z3x3OJw4K3gVw2DusBr35pVlji+U+J
lu3tzU98ZymHF/owoi/tIPKQ5vbrGCrgG+spNMWQFor0WBgLgjYV7BrcONCt+Xvk
BrbqiDMbesDwM0p+oEl3PuOA+PrtogH+aO5U1fsZjeU0tMo2vHsGST3bwXzgr7D0
sqZ6kj+XkFrQ38RO14UfSJxUKVG0cqcINpNo8e+ZCGgIoaCWkwIrVWhQFxgbeyGJ
yNlljI8o2mrar6Pwa/8JPNyLxmEfFdsRXCN+YLbUmzYcFGE76ezGRtSN7uj8Lh72
IMXpdVaLXfWVBDtDsAzZV+tkJi0f+4Jb1NQNURP4G/Ra/wAx+Ai5PxQL1OV2Jhw9
ClItFP7/TMK2Yel+NhMgTAriRR/Qbo+b9GcrCv7S+qFDYaUSrOKlfeKGkpbCwrc+
OamTT1R/zpGh0ayE60eHEfBb6KJhGSpvRJfby15Q2cIUo9iaF1CrZXz+bQVKCOuV
IoI5wzDq6qG8PFONN6JCu5Sxdt7WW7FGZZ1RlG2qFxoICD/V6qGg+BdbjFwAmXNU
pNkVGz7M8D+HHvp/wuJQsbkwqbnsT1/mwDfDI+JSCHTNqs9Rf6XxPmjYpUSEQDWO
L88Ho55x2DdJ7poFlSSWa7vQA2ehGD5SKRiyEHt1AYB1cLumRrie2TpEJSnFuRbu
2yy9vVxTAvD+vIgCdc9uAuxUj0f52S3fPxwI1rhY5EkYSJoFs7Jyhm+FU8hP83/v
mQaMyrvfmjHrwOG1HG/AQGZP5suiJ/1ONLKD34vBVavyf3ZbOd6FpLmJDE8JULJx
3YpslYotqM3LrfjjKEnZJNGVx5EcU7LooUdNWMUVpTwaijXrlfBwC/F0EqWTYtoj
OX82btNnAN8g9stpPLXCfSwpK5tfPGRHibqWdnbRAs42WlNktZgo+o4FyaQr8k8W
LRioaFglkbacYKokH6Xx/2sJd6XP2Cwp031VCzIIm/cTeZ8AbBKqqREflRf9clvt
tr+otX5zP0607nwb9QihY8/5aYdRFhtg/H1qJqwr2ZjuYbGXhAtwhUXvxgH3K5e6
mezCRdH0LPa3FFpoupRIvpxRzZpA6Lu9WkvDA1ma4F4nkoagFkL1zdpWOyMxt8CD
hBNefHtXNUACg/LPKpMyUir5z45fk87qs4uRbs6O617BMByLI9NN8yUnPuq52qyd
uXtawnNWmXZZF1c1gnTHLF4/C3I0xPeVvM27/h9VVj7aHZ5W4nA/9sypnoIi5S/s
c4mLhm011kseQ5DcnBND4P8A7HukGuq8CU/f7mXg0uKVF4839jLW9pg+5QvCCuIu
U/yCx+tx2qyrr079Hwz6h9OwqIP2iCU9iEVGbisGubU2Y2kQff5srwXwNOw4/8cL
uFdlBJXJlr4b44ObRbyghMvHa0O0PMVofhPiLouZBQNVUJMaheRUR/ecbiNN5SjP
lC9a7zu7fQv9ynYB6sQpMERTZxGK01/UV9aU3j3vXz/fAhtCJp0KMelcj2EKRuDP
Y6JDl/eXf/4tenJ8CClMMePLaD0rKEPx3dUaxTsHrwWwmfRMLMZRlcR7Z1HKEdna
dd8bi8T4Ino47vLDfwJej5GRYFpQqljZcgz7pOsJxyu2POveZJTbPeWewaCAs90B
CpfPzaGMlzEchuIamh8mtPDO79gEtdD5wFJSUWuZaNzt9X+UnROYKK4EdWJXE6Su
z7VI36aKhWHQOKggza8solvKdnjbvZlu5wdTNCsE86XfEqfYNpSWnUZYZYC5HsyC
Atz0ZcozqMR2Plwp/yEdPhBm3fOlrff388/9a1dRBuvuxXx+k9DSqoYOQEiKy1x2
BxxTjmiGQnEoe+IDhD8gH5NDBL4zOK33Ew4bkfpC7NArffwyMpvaRY8wQ9Tx4/Yy
nEplK6axbfiHkf7dvPZmpV/OZnI2k+OXFqODqSjHcl7VljTG66vC0vdV2MCdDqXE
9h8wpZbo0Ota3ysnYe7Ai90GEIg7A3sW7+7abEMmonGNYFqPRCvbGi9NrIUTNOgT
G9zeQIs4PQcLQgCPvxSwd7XZlCAsSLO61ss8+uxiETv4auuoXJf7ztSAFS7HtgPv
BYj/az6ZwM00Se6MFWXPinCUjCUjSeSqNntjCq351aESF/DwnwgnWZT4J/I2ScU3
mxZEuDjNLhEcRa2fBs8SST50SZ8LpwahchRNgYXljnUqgI6rOR2+L7yFCBWrkOBW
61jJkcIqxirUfQBMfL//1zBJ7sV+iA2uGXJyk7qsyY/Np0LHnhSii+8P+1+VrEBr
8S27CtQzQBOPTXLFRGAGqlJX9XCm71s4w3GiRJoL1EHs88u7Gq2BSpP6yHFBn5Zu
VCK+jhe7sLkgQEqjfPL3dlUc22q/80crYMxc8zgb9Vumtq4dPzPDIihGVXOmvz9T
a3N+/8eiaPIULBshi5Wyg0+xesoaQrI79vz8Y5oLJVis7YLQC+l3XyaP9vwBNyv9
QPVnA1Y2PlhugmXs5/cs/pnFWv2ET2XQk6wr/NQ0/GlEi8jfWkF9sDDqXo112wYV
cH86eDQRucydxdF2NKZ2RSq7KRtNqnXYO3vdSUDznNmA72bjOF4N6PuA61WsfoWh
M6nqlhdReKK5zcAM82Pe2fOVZd6PysgCu3gSuFBhe2mjlaWNs/Qr6+djeudBtf5V
WN9i5mCeTkEFOt+lmE0X4xFfbiVTFBiSxlWW2KhFBxuAZA8B0pc7hgUPOGdRIvoR
HbwP1iton5cU/uCjkbG2SZNFR6s68U5aTYIDIujeAACKwWO11Mm6Hhw4QV+78yVH
Fr/+7587TA8ZmXGLGDnPDHZ8aRR8wh24DKOQLEHozs4xXwA0d1V9y5zXMDdZr+VY
GWIeiG9GjnvvLvdJ4BXZRAKT90Fp8/ir/SGXDuflYlZyInxL46Wmutdx+dbJ8MJl
o/Kp3+sSBEkhY5zSS1CU8NYHoINwrSKmdrbk2y3NST2V9Aba7GItBfAKOEIM+YIQ
ESobgXxZZAbJ5Eifcki3w4jVjSoceZoMraoZ7HGpwZZyKOP3Y6Unl87/IE75lBkW
qRrHE6DCjHDByVD/XZLnu5jDS1MAGf+WPb6CUkfs3xdGB8gQQIHioWkHLBAHDpen
pYNy0b0BtfCDBvpPQdX5a/0zEXcxYNoUmtlJTZnzTeqjxmvOPJ78vzhBgrZ9kh8e
LBvBPmAvQlxGWrVCyQZ6Lz3xsfZ5LyG3VVExQ/y1q6cp+KLTQhz91tK23Imzh/l8
c8PF9rP20lqpqRkrkhFzLCmxtgkJIQcl353UmAygTo69qxVIqrjGSnW6RV6gd1nA
z/1lC/uww2sWOTADj6KFGKrS8XFHnCXKRN4iZeHPfW5AtqM/z7MEr5A3MN6rTuVv
Kf+At1dmmDQo7AeTPa5To5kt5fycnUmsDO2TCeAWsmzBkQ6iI0qJ4nsuC7RwvMOB
Ea+91zbuv77ReFcUnfjPcZ5AuiCSYaqYReCHlVczRpnH66cLQ4kGsSMNt8BJCGAX
8lYCaod0XwKo+sgmHl+VuwPm/KV19zwMFlQ43LbDL6o1UpwR3gjarariCoTjVMoH
lecQl/BjJeY65G05ZKhSmtTTdLalhKlCFCRMpkB0ENQUGZKe7qMprptf42So11U0
1ZTHn2dYxTscvCbtYS70/Oma6Oodr3XjJ/fahUlzmOf/VctiLBiJ7XbMih6baZmM
K/qyYArkIXS8vDJcnZFwxv+uFmKvdLzoh+i4YgB7SdMgpBVdciEPcYz4OytCeMLs
lEhV49+nj62yac4WljOP8xc2sO9DvwCudFZjSL50jqojSCbeVM+Yy57RqAP+OVcW
i4dUzawdgLfKtY37xhP4e33ux1xe3sSOOw8QQEd4vBD2ESwzzAtkq+ssOME8wwwU
7dKhhYcFkXyXfx2Ao7sv+UrRR/QQza7nnULAlpcFwyHq6JUxjtCe3IxWZ1bd0oRT
U+gMYihCyyW00jv5f3EMdPxkdDXAK0CZQFU8rRn0tYPGo98ZMWxKqLbM7WDkHVic
Fs7OiPgqlUhUl0CYNMIM4Jc5flsQ1INNuVLySeu3Pht+HgnmEGx3ZMXCLtbEwpGr
izogJ/llbv4Cif+bsyY+35HFQ8NtTTB952zmyPUOasxOnQX5jKpA3Diz7WPjDus8
PVzEdNNhof7R3uDXUNfmvWsQMeoSky04Yyjrdl+5jLazZa2pBC93AYPmL2Gz6ZEr
89AkXy6/iiAtmO+NsQ1Px+YjnFbdVHpBMWJf1HIiVrUvHF2rYLHRvoN8hqxukqCu
Fnoth00BaR4TRmsEhpQfOmddK+gbsCs8lsePsYsAV+/nTq3ALGQBECkVwfjANlje
Dt2XpbOaXMPG+ESYjtTEebzi9mLOvPxszQPMnRd5f5qt9h2C9c3f/PC/Gkul/Dro
i0FPYs72y5xcoi1BIV8Kw9XfF4GpFJamgINgs9zfzd2pvGPLAeM1sIz+u7N1atWL
9A8BEMyTdJrFx2zRezotH+eRZlli2J8nDjA0A/EibDTh0zbtwYAn9Fd1fCeZ6OCS
FUqc6wZ06ki8Qh3GVG0ZyuxIlkqlIe5UsNPUg9wEQcq42LicrVF0ur0lkAn1tHPN
ckqnKvm54dYpO2mLuaYUIDFPwu+1Uw5XvZPxACm1Yx8N97YEfLr6M9I9SZlOp77f
XRd1Bby7FnZcMYDr2VRyEdUVFC9Gzym/gaAqXiVbp9QGO09rwoPVvAVv+NDuOjx4
3EY7ahL6Ai+E0IIP8NHoVPgyib7C2xMZMiVlU3wKFPHIAUhTZvf9G+sGsBS4s0H5
gHbivjbPIhf9sKXb4FDs11nrW6rhkGJqXa18U45T4h/HUu7znAyy3m4tO1C3Dw8Z
6TgMh63iYmlUO8sv+sJBGUo70kQpWHYETuEcvN9GDadyAxkBELuk+xfgNKy7/7Ty
f3F5BCZxw/pW9m5jVOuwG0ew3KmUwCcbLVYGn+7wbFiNZhsRDYjDX+H7GTlKdlHm
iiwSb/2dlBsWYudebcV44JuFd5BNSXbi9fbtiW8LLuoW9AskL/azTnz7WFDd2W6C
BNeo8O4IRgimVx31Oqx+5XJOddVj4h83pere+Mk/xCpI8WykbrDgIVxPSvGqA3Yg
nSrhzAIcT3rGZ73FKA8ul3qSxAggn0NC05KRp61svHaSse60uqq1cnifwSnXWtBC
iAL/wbSY4Gnsc58rXFP2MHAXT2Zs2u+cj2eLjQAXUvTfCbEPd29sihjpd2V79uCG
qdIkPKiYUajkwPkFrXMBFwceN8iHKnHCviDqakKulgKIP0sR0XMkaGD8iImNHMzU
zJKQCofPgg0mAE3NZTDN/dozpgaMHV1x0zslyfusLC1mbb6iVGDdn4nFE/nZrQ7h
hO7jsWAhBDapGZ9BuvnZUI1vq+GKsaAZzkXH66QeC1I2WtOon0N9yTty1+ICEa4E
hdzwkACdxfcbZ7JOAoa7wQPCD2Jvnat/3lxHsUqrfGpEwgtlBb/WlGFmgDcscIqt
LXE31KrT2jUO/wYXibFVHediAzSRitUIa9GcUm/glcouZh3mkyExBXpdvrcGxOI4
ZnrI/fU0ycQEu6t4+5mC7CTGo8m5A/YyuOjp/x44OmiskJAHwr9/oAGwBn9MNYWd
e8rTla2RyX5yrPfzGpUc+GwnniVmIczXdhMX07O+EEu75Ff84c2N6hME1pEHjPuI
1g8aEbxQfqMhM4/5+UbCjIgM+8gZsiGvchn8M+QUvkNvz/wodLIICzLkw+RrUB+H
E5w0rWo+F8dRiUkWHXDp09EfhbWCxlCNHilvxd2W8H7belOJ1vC/7sZx2F6UMCba
0iSpJmdsoTJLiVL7bP1OydfrMZcTOmVvWAiDOqCS4NnclZtUPjBY5HcBiQXtt3Fw
0M0yvfpld6teHsC2NzCm4UtA3k19WCuSnFvBW74uZdiQrEu+P2/6+hd+RcMd4p4I
+j15RpM6pYLoJoN/JPukUypaCwSVyDCRBSzAloY8erF0vqkg38laQHdSOPHNkYh/
Yx8cbl6LmFPx+OGTDNm3t7wsdfOu2GzdEWEbZ5RFBzdfZ2St0OszPnUaVcx/Welc
tDqAFMkVxDVBVA3YZdsGgV89jKRnBZjAF/I9jTuXA/CxGcNiNtqj4rRM0Q/Syd/O
wlfuLyDnsfZrM1vIGm9jK/cXs6LpHzXwJh63FdiXC0Y3G+6u4i5ws700P6FATZ9r
bypyLPO0nzIHlRaNnMRtQn3KAA8sRF1oQe62wzapa0v6HBNIM4kjZAxD5A7YCF3v
8iXOf12UxVxvS59s8dCSo1ob/nzgXswW8zs6WLE0+q4LS71nZSs62zaevoBUoXVR
oZfMDK58o53VtQj1RYz3MQTeG9rDt7XX7vllIFzZ5xHHyUaO2tlHtyPcnWmB8j76
dVWYOeoeX+WhvOqjzvqxaXYZ9XBymTFZ8yq3q72ImOWn1vcrGJk29pRr4bcGHD9X
/R4xBtquRWfaJvsUXulDxor3TYIrs3v0Vfxvx/2sNKVG6V8cpyIJEWQvFZx+MQBz
dFbbyW0w11e3WzrigoTq8gymDbjNGYi6yle9CK6PximT/nwUKW9B+Cs2ovFeVWwT
PwqcCBV7ZmdhqIgTGlTS5gIkF9Z4YocIV7tARegDGjIdm5eKPCBNWG3ABAVwcZjs
tLaKRPfVNsg98AiseH7mvT+v0P3Fl1CRXqFgWYHlnkwWqhVsAUYkbFWMm+CIDmBa
Qy7lF3yul4pi6DZQ9ab4lm0Ip3fIr5yHF9RTT6i7tIt+PdVngu6QYTB7EBLS7YCM
Ss1TFYf2qWqgu23rjT2dWiHVxJRMazkzHyk7cIuOr+jLPVXbFjujXYX+d7TQIhiW
0KdcP7MXGNGUn9yFZHs5zXh5IKSeTfAwd/xWeAwjnT/iug8HYYf8PksK2gcHciOU
8CqZZlilJ6w9MgxUhKV0DzUvKsEKSXjd9DNxMOvbs4PKvaj8cVLlkGaaX9STPDNc
/Tz4Q6mP6V8Q6ka2aCCtfZmaf3zdtKpehh+A0H4C6fwb2cSn0GQxjyiR0cubLvCY
F1Udc2brv5A3A8rQptvLBu55FCezVwuXDgWC+Ieo0nau7cHjWOAVfpqor5uRG3k8
drzpUkkyqWyC22u5oYyPEJcET2pziWH/xKYEYTTcyLXZRA8iIoEDKh1EiLDv3wFP
jxaFhY9OJGRPkObw7SyH1J/WRNTHK4rm9hQb89KIu1QuGIaKecuP/jfMf6y3mzzS
0mvQkFVisE9c2ixNe4knf/WoOtFSXUIJMIYAIBKpcOw37AbcTf1OrPt5S8wbwJgp
FILcW5j0sOHQbYmJ7PzF2RRBasn73nLoW6DQf/kkr0vCPDzw9qaYlpitDFN8AYmI
57p0TUcokn13xL2gw/+/+OacP2V7snIADov8G+wqXxrAmWFQnXPbiiRfFuYsXase
A3hqIsKo9u1bpH2Q7lZfa3F+sVZ9Q46bhVeXmGTqetOKKYYYdidpfewAyqOA8BCh
YHgM+soVxqGmCOCtb0G0Dm22F9RI2uLPJHdXYxZpq/ZYIl80pYCfK1yyJgRv86dt
Sxx0CXUlpPvp4x41GPaVYxoBGsKRniCw9CsRUrPZVDJVCbwSQM3L27woxRQr4LzF
pN0+IgmMQaZa853n3PfBxcpSPam4+5KxdcaechoTumvGT9cxgYF5FiduvCvXGINa
xgZDVVnxYHQHooCXf+gjF/hvHRfOERlBkOXMwutRlDAWGUHmj4JHIn1UlPpB2Ul9
BwEcVGDMURg5vqod1EjYTft7DYSeXHCZgZ/eTCugN4xWXDu59vEh5ArN+D+Ye+P8
V7EUr47Y8jAF2IPijIsMCdlfad8Ss8gByuKGh8mi5cvcmgXXqZfeQswloFgfNWim
o5ZzVymzU1ziEi8t1SpUXXcoFPlvmv79DriO6SsMVm3FMTQJ/YHhStLFFKTh29+J
sTEs8OkD3HNrnbq0QHztUVe6LiGS7QeHNmJHEy6RqT4NXxkQB63gbJtxniRMBVpw
z7AVhnYIkwIYrfvU66Z8E4l/ndMV+Iuv1BL2/B1RvLBHTKgZ8QbbH3h1WS46Lexk
g178dWuOZpTHcE4hpdoti76rww5FV8h4Q7ZpEIkVwPVV7njE3MSjswP1ASX5ip9k
bDZG0Dmb8E5fdBlQcLwdFJm5EMehXD80jee0p3LAMHhcA+Hh7SwsGI4eD8n5/Ttc
wrtZS/ZGJjoSoq7bwUOkr4J4NrVTbPYf2S5gXw/ou1zL+XGbhWesTBw/Qi4XysAj
VH+8rzjw3bqzuJKKgxa2z9kyKMzWREpS0RhgAxOgR+992LHGwklW+1UXSR/x2NwE
FYi1AJi0SmdaP5b82AXXIQtQWqbUd8+5KVWuKhIo3fY19HFa3mxKSi2iJPZmUvie
lIV/WUy/zHkSHQBgDai2tFGS2qxB6O4CWQSkQ7A91WramxK/2fUimQdyYisX717d
xJ+ithS0QCTD9XEyHkKcUQVBFtw9OVCkT84VWD7yFxkIAl/PobgItFZ54QNAKLN2
+iXoYHRrIyczc30SyP0j8fNmwigAFXZugUtn5c30n7C8nzzqy0pz0qq3lftDbNCV
Sk6d37oC/4nlxr5dSnfbTMYm6ptB2wHFyV+/6xgIhD4tdR+erssYqDByxCeV4bBs
jNQiz807GNO5K+x+zl/jkcQkTt3W/IIn6BaxwOnLV2dx61IEOxkAP2nFxoZFk3wx
KXR3xbls4aZU7um9zYJSShfxkCPB7eUKb1n1qTv/y12y2flyM0YJTK7g+/D5gT8k
sMh4u3bAWdho7kfBnb7er1naFfQ79IOl78BmoAjD9IQrPZudNf2g8yfGPu3mrJKa
2g+puEZutL3k6MQfJP5oatxPVmRa7Pq6Rfc+BIrnxH++VdoDxUWm7sqT1urJDu3D
aRSIyh1NHUVkPc4izQQ8QgJxDzH+zyfpDfpRyPAdMp4d38eWYhYZHFJc81cTh2Hb
mK/JCCXOoMkGRzTZQSmpYoXLL48w48cBInlogGjiYBncvzmirGwkUTTCzeVGpLRQ
9uTqh3UewwadbEWyjddDjeaOgWbmc38pqUGPtEC8eorfflTF1ynhJbnpFjcZltWO
TEqsfuUO106+3OiVmrTIYAIMerndxgBZ1bw63Vxcmo+LbBzlu7N2R2XoolTCa5x6
V8p8FUMysMbrPhJsF5DuQRBhlEyZheCTwiQr8u+8eAHpmkRKJaSok80MrwX9XxU2
HG6upjqaP62Ew1Y1kup8IArRvNLhipqXgqDaFzKMXRr6TMiSkIk3eJY4JwK5EDGZ
4fPGGUlSB1XTQ0Gd7jv8FEzPZrrmzbithTxgnLd9iHQPTXbux4o353RryI0uEaoQ
o8R1Ap7yoBnxDN6asv7LUf51V9RJDK/ZQh/YytECxllviHua3hWu7PbosRlv1fip
xdF24u3oWaqEtXlZVLctgUeRX3Pv+mE7mKIKPtHUW1RGP6berY+ExKxH07cCHcvo
zBCxXH0vHVrImRbfcGwQNvclUXoED14sU1R9ru5Hzjf/z7V7keYbZ9m6EVUNfGCz
YeMhyBJsJAU2qwvhLVHONyY9GBWVamsxyPVAu31LBh77Z8w2r9QuvERm7E/AUtG+
gN1FzQFBv3wxL/1/B5ElTt3b68OZ0nXCLL3dbV6tcsQmDa8uJQMl3HzP+5wqIuhM
CcARYC5M8ebw2nue1bt/OYKnV9gSKCx+xnaiWeBi2Nmgd18quwUNj6Ctia7AFzsh
8wg9PnPqqxqtOmqK5s3ZQhfNDSJGRVk8WRl7fXWb8L1cH4sZXmdeieRgbMIIjOXz
vMbbaKRab872us+GVbdkfwkRjythmxyNpUXjozjoKDvytTrZ1BZjBGDBUsrJLzeX
ge2MgOptMKRdYVGHX17fQy1DUxokxaq0/HVtm89CRtIKuewTVGWouGLNgbC1L/9J
pbYbBFtfxnxPzvteDdyaMyePLRpQERv+YCinwOZy7ZWBJjgagxIkSrf6kMaN4NFb
Ps1M0VzKx2KPXD3BRNftCigwUc90aEmKVRjv9UmHeyST55Y2O5oRtdVzS5RotNfE
bK9yko13hSZhPDRwTC6qyAJLHo3TXuIBrvWuuRJLbZj1LyBotyhFdOXX4MJJTsw1
wLqISAt6XFCBwuZrcT7ZfTkN74Eq8KsHJ9x5f4/Jqn3+kea5J0sOcqsT1n1jPB56
Gn3N81hY+QQJ7u9RCXMX+h95YUvsqAdlfZfoSxPL264cUXysaYtRfkAZivJY825h
yArl3iIqIDuAMzsTbRsbcrF8dhqb9AcCOUHv1D5dZl5qKdzKp93qLBx4BdSDPYTY
zzVudfYEpg2kF3kETEKguGVfN2iEVXJ7DuFqLkJXoWsNfg5GLoe5y4YVgNUSkKIi
Zfw1Da5zMeCu1TWPXlaxFs/PTQt8jWN6fApSzL3lEKzGZY0djPtyhN4S9cFJcptf
A0dpEj+CNYkd+3QUoqWrfl7tRktjcRnBc8WsKeanOyYEqeofgsMgzM+HOTG5IuAn
wELPuHFu2kdBnNJbzgEz0fZ+T6tyabn6DrejRSRmVmEVE66E4Ami1Z/wUFhxiUzC
Wzj0G8ykq3lMR5yvP3rtjL/BztrrnZg+T7eNrz2k0G3o7lDeDFdVnI//42ea7GGu
OVdqtzjnLUvQlKIVpctzsZLbCX29YouKsx4Uk499M6Im4TbpwAzL0KU8Q5zho337
qsncpjCctjwnbLE5Mi1O9iwuhl7Hn5qsfVdmikDX1JahCxsMTSKVcgWYtgFwG1sy
fV4F6PmCOOIES9dTWFpTZNRBpPFkEGhlDzBE26/XK/HvcVsgolBRiLJ0YEom5AvY
8zFvCHnIrB5iin2TZ79ulwK8C1gBHCRPjEmPzdps4Hhz8DLxoZXa16zgzMsq4m4g
91WFgnmuTXncpaprofO23S7rQyJ4fnFNd9LrYP1XS8a43op8MDBihEDa3VrF8L/2
EjvE4c3nF/P8HKXxBdGJpa6lZcF1kxqECguCyGesDqWH0Co61NB/AEKbOpV6gcy7
NZjPgDi1qLX+YKFuZoU3nbVmDQzeSpU0Jlg+RHHVnxlYOVdtrhhSrvM0cVS25xFl
L8VWHGpUzJy8j24veue+R5VxkjguDuO5HI9K/N5fFAqs+v+vrR7ISvOx0P97yRbu
1di+sgwLHn1rW14fu7cX1TQicSdDdknPbMkIKJwn/CPEN8tPq+ILUnTcxUnFAoZt
UBtT8A9yMjE7rrVyGzUxLNnJNCKmi/sFJbawNSsN0rM4X9YaqvH99hJvg79KZBKd
/N8jDbWBgsI1cAAIC4qBFQjJNkLKzrUKzne/4PD+gpGQ4wgUrtzgrOnlKe6zjnIf
IS0/7Ur07SOdaLe9SsTHxQ3l34n8e3DxFdyTsANizEZBppbpJea1XGlIs6yeST+U
UfX72yhQhokGQCg2NJlo7qV8Ez39mtvDkLmm0ErCOCSz2c5qmgWt1m2T419nPKzv
KxQz3hwpwlYMtgva/kYWxKbudznKOzaFrieMHZfK/Xx+Q/hzFJcSQeDtzQQr0pGb
mQag4r5PqMc4H/C3Z+JYKRSayjTbk1bqQI06R/OyL9jQrjSElbKTdE8wdZJjTHxm
hfAndVW7agDjxyNid/BGpVRByixhiHEv426QCWD2EkJ4zibuF3qAPE7yvJYjbyG6
+T8AslDDTj24tSrqx/i0JedbsvWZANGwJtYFP7X30093j/BZ0z06N368tL+oB54Y
k5j0t2//rhnF5dpnO9OMNxKcXkkZDAY0mOGVjApmPtUCX0DVYSY5fRPkyiJ63GOM
yK9OgGc+sYnJ9cABhXMeLZq2iuaXYQTUBAsCumOkYyZnqZ6WYcKAX5XL2ts0Exuo
j1FB/m60OmBeU4jRVh8JMunsInisEqESinopZeLPY3rNvLR/d9+QVcY9jgh0mN1a
azM9qK2BwMKzE3altzpMDtWXOucEwApDZXbLuYCe6qLgWlB5sJxa50HJsoj3tTSF
RMbbv/hhwPfZlNGX6f2sRe7VAMw31Jfa+Zie/JbinsBuJSXCi6geivkin3jVLM8F
adr13KCOWvGOBjCecUqsMAbJbKSczAhvp9dFqVYSUcYy5Ddfz7/DtU7uFMYzgEqx
7sO9qlshi57PXwsg33/eLv7SmEW+XIKQN51qkM1UbGaTlE8OAv+jHc6kM+y2JiwN
zUbhHSsYF1NqTLwsT2yXEW8FUxurTZLhc4AVFIMYMFytiwiYXYNdGyKTMUUGrSI2
ctKC/lz7LhFVeNJUFogrOSlX/7ZY8GXQMrnuDw+viAPVxzsuqVSKFSwBml3Y7Uv7
4fbTt2OPlscBts7MXWdOCjKg9CqGDHPrL9rxaaa5Tf1hzzbiSssB80QBNRm1B/kG
ENO0VtIxXDNYP2YX2mHcTPzIXb13YWGh80cGodxzMP4IoDNM89Pig+w6Tv9BiZAr
dfNntA8dEJ/04PwNFqSom4txjJgrgrLr2pM3KEv0T50lVA4NtjMFss0iUV+kao/K
F86OMOIawOBQWbtGEn+nUBn3o0aNnewOGyqRSb8DlENjpJa2YVvDebAm/dzrp/I9
TPvF0Jw1ehWfLX6VAIbLmWkpV1niovwQgAxOa2H1u7pXZgql0l51BXdQHBflx8v7
nKPFTGs6WZz8Qxj9ToElZJi/grb18vqTFgq5Cc/w+ALj1YMFbLb5SwYbebzttHKz
ODRZNjO/d2pHtCbFL/GJU+WLrrEzepa8iIuvUTAt1nhAhz5YWuc5bFdj+X2ZMlF9
jrlbrPA4uO1oBOB5e/jTt+aSUgRdkQGNnVAP8mVmhr/93T5XMM5jn3kLzRv1xbZj
0r7/+UWm1EYWUYOGI7xo+RXj1TEcTomZ570fA/Ry5BZhk6FCUvTyrtPxF23P8Se+
oX4HRukieXPxOhfNWZBLULomoeCMZdq9VtiqPkiwFWxPPZKfpe3EMrRbJphobNDx
7brhIYs9bSqqCviMHvs4LZcCRMq41Dr8g/luGpHUR1j6sjpVbq9uJqM4fVIkEUJI
1yf0gDHmSiVJZmwitI0WyYkcx9WR/tExtzVgx6aQvcCG+4WE9i65L7Ry7fRkp02I
3wGbWJ+WMdx61yAGwU4Pdqv4lSPsgCsLrvkLuOVw7PSx9aTTAuGHQoUTseQr1nWK
+/ZsKypmEQYKL5NLY6IEVs4nGCRMjjg8FZ7ytKx44zlzJajAYeFPNlk03r158IdC
euOo+nZ4lcbxAQY7cDAFSNKZIMKAZ57z2AuX1KOFlOWmNrnDh7blbT/oe2jy7QLb
5KT56XM9IRIj24nzpmP+8ij0Kdw90VMgBbahQz+l88Zg4BflUDuzUjaLHWAxnvk8
DcfcjZ0rjmZZj147VK6Li4NzHBKKv9REgbO0Tk+zVsd0ipQomCLxDb6Jq/DHfBjj
Ywm7OqT86KXEDS7d4ggyLrLiQYRphNSa6sMSa9SAY87SQNbcSzFne2kSFbFZCUtj
65Kn/7sO46/53yM1yGZVexwVMOo1kphaLlCsDiIocTxCxfK/PYeioNZL8Wt1badM
Rwt+YH30sOF62eDilD08cRYG9zmGx2aqXE7MJv6N1CuGGRFdX+Rp9PxPy6Zy5j7z
EoCnvBKzwFUtIyXjiiTKJ7ZDS2d1nEl968F9krYF3bs3thlQYKrgv5LcXTUdY0EK
pfEKCp416SGFKCR0rJHUZQ5y8uOuT63o+roFrUzsu9rR7UkJEQ5BrD/NHsBpZ0oX
vwPr469lHj1Myy4ypGIYetWJ45EwdMAVAaKb6y6X0IG37tulqL9biCYka37AV1kC
9KPA1SZmP9VxE1KSyjkfg6Fdxr8rmbUnn5iHHfvH6ddSd+KKV/gHPt68rgJf2CS6
So4Q2FfsFM5eccmYGECgNvHEmgnzEyvgenOxZGiQ/ifTWTJh9EU4RfumdJVzxKsj
3q1ce7XHeeFJSuqAtTLcU+EPYCiJ0J/xH/u1RaD4nl9wTmEt1i2y4EcS/XUPBWWf
lcGNYk9XKNfRboF11uSVmNWQ7pfNZUxGyOnqBMQE9fUyzNBkV+uWPyrcHgkLopLL
6zKLhea3rqcFFFxdO3JrIXOgyIG9ehT+vIpncAcHskCjDP7NFRQGcHeh1xZdzm4X
OcEvQUCUBpZq0EbuBGYNWTe0E5OLUPABeRph3QrK1B54hwlMlLiatS3JbkAS2Few
KBxjSTwk1m7488Etx9ompfqoAZR1lTp5symHl/8dZ81NU3hD4AZ3D/JvHmmT+ZIG
0J3LiyYk6J8eAZq15z1YNPz0YhIR90t8xYFlY/mvQqaUg8ILFex2RwEKr5II0wTl
BVJ4vjQYZnfQmvQ1WsHDEeI/9SV+xN8586HKlaSwGww8huMxQoBQ05Mrdt5+bWVb
419XbPSAjoRr14acd4VRciM5zFSyXFBSM5X82qUmQ0EGA2yqOV+7osbQNjficPkk
jAbvYS/NMkdcJVLZTW+UG/T+mnKOlPFKadCJqmo7Fj7ak2cMo7o0jBhxd5eosu8o
UP8kNivo7OWvoy5wPR+SES02gwvONrvXusqGaJKHT/r75w4HZXlh435jFH87XJeF
cILnyJoZOy0SxjR0j5spN08iWkzFzVzEjWgbohulrsM3tuGwudNRl6R1fxEbNJ3r
hodR2AswrBmDmR0Kv/vLm7VInlQ4ccXWQw1W4KCtw/ZwR4oRfkdFWMa+ve6F+4Yl
lrQb3fhJGGqokjRKSBXVuoiT4FBJ4d08NY8t7cAxaDlDQxtvlu6JRZk0Rjrk8J0r
Qy6J9nfmceI//cMrGqdal3fs3GemK1TK+j92oEb7LZWbBqbfYXAZzIAvz2WofA6J
03/FRWX9krILJmdOhiv36vLDkrXo7gaAzVX+o8Dm8zYEkKXQFFuFSnDIS3MYomup
FEBpl9iyzY7mYc478lLnL0LuqGerysV99y8ndemI/5en0QC25wPAcpBdClsu1gQT
IUR+bC/XwQ66No3Yg/NOKV7IHBBAfIrHZn94FbR5tbhin3nAdSdkdGEhMY47CXAn
D5gh+n0JGUVfamB77OwKs70P6NINYkNdakUOz4XB3LCoE0nTNbo/2XTI+jZPv9oa
gFlklLnA5KwNHZ+nhxateWwXpMOegOJdJ8I4onJLdYNuwcn9zRDAxYGTe3YzOmVk
m8zNtBwsTj1+Go19mpiGkzfj1DWHM6BJacfc5aBSQCZNiZFAK8DPNd1rJgfKS4VM
onAeIDYyTyWYMEM2QkE/yDfm42jzAZ9KCYMA/c/4i4vXXhpi8j0Tm5b0Cu/Qkt5N
GonhVX5YQZx2ovaO5kz2bpPcNl0QtTils6/xA25JHko2sPdUzeilHC3eabGqXjsq
pjHVx/LmI/g21is7YZLfg8CfJLC/t3p5UjcrO586B6axwuFdOi/MDebQXL9n5cPo
hjvHaqq8V8BREGcloP4wR7zdHHx2jfgiWE41/1uJztawBILD/Mw9Hk66aAfuk+r6
uVZUxkWDD95nQ+3lUFsQ1X95VWRHvzvAU8v6x3/IjzRiQxJohLEY/LiGFYuODa58
JT0plnNv30zvkJYHhCg9uaW9MgtTTManeNFTPyf80zTZrf6np5rA5af8xCy116Sc
m6ilx50WeLiy/XM//ujWOfDWq4Deb1+1wXR5W4h7zmHsaIkEeGJpByim9qU2JR4r
CFPflTmSYKIjWZwE1CMCigUjzu6M0xARpRv7yAudLA8KtyL2iKzI/n+ji0npY5vA
fVzxaw1FqJzkdvEuiguLZ2spIUkd7aQqcJ+2Pz6LR73hW7PQuJllY1GImwFgodCm
kamh/bj1GZfhnmS7RNqt+wDlnhBUboyQk2cKISx9Penk+9fhH4eZopzPPcB1YMLY
x8sYjL3RCgheyhsQWOQV7aFXSFag9TW3Z18WkbPk4Y+K9q7u4LIlwdLh1TxMfldH
sD/YivjOGpXbbhsROJQDNGPwu8rADDgFu5fYw05nhG/AMqAOt9FNtHdt+fyAn3td
dVYGY3M8Gl0qWtjiJ4NF/A4abWAW742K/R8B+dXDDiH0wIpkAmKoRs1lo9u+ePt1
sfLDJppcLnoeWdQqtrGGRn1smVjSej/Wb14waps5mSLRDz6MIDiPq0GQe3fjgTsq
L+LSb41vWpDOMGTnVxvAxUkLy2wNn+YKpsT551Dlz1OndjwMVfZ6x5lv5yZ230QQ
hWkM+Rc2Ifyaq0VXB5oQcBV70laorfJDhjO7dY9c+/rRuYusgVANg1vyCugGopjf
6Tqf7F0hLBjUjF4S3DnJTO3WF3iDWHAhIWyDYp2/wY7ouYgAvucG5NG74o7lYhjn
VCc+DlrKXFTcgDlU6taSPGAqgvJK//zE/YFJtnLAsY1lFvMPdf8dXeDGFFOpjJmY
hu3xErfatEC1blj+glixUk2yhZ+lZfYozjkbOsm2qIlD2bAi7vsVT/T1mSdxogI6
FPKb72dBe6k+u6cKl6L/O1IBnELqsEixo3dz1/Xtw+D76m9+pYc67CyP9xwR3rOP
CQ9ah0gryTdutnQhp3zwI7opFExbEzlWYEzFRueYbpBKWWTR+5Uoob+na92+RSld
/F55lNNWGpg1BgRaQW7ygH5zusiA3mucGmlqcu+Czhl2/tg2gL2KLvWScKLSmvf1
IH8XDBhCxSgTlDlOpkq8zy5oyw6jQgiyIB1CzfeR6MxK/+5/pGSUM9lbKdJuKuoE
r+C5q4jN5GygEqAtVS+iAmUCQ/tx9lDSnMpQ8/YRh/nyP21evp5sdaKqJxs9QdyH
rllY7NMEb4AbKqcce8xK3Ups+dGowklA1bmDmDANZ4cXSHCndkvBNfD2kNiP9IRV
gtZbPVtzOocwIhS91F3MnLGCDYWmdb3AAPlaizcljuUhYY7uNufr0yyMaGuZC90m
APJcs00uFGv0Uijtdnv4Q04VaNY1LVXcL593uz3l5TqGjIlWkjqCGWsF2KtVjHcs
IOc7pWL+2K7/5CLcLHiecM0gyYCGpy0mPpDxjfP+nzb8w7VHqJLHiv3e/GxZWDV+
97ikq0hpwzzbdIgvKBUM1W1ksRHelAkKbviN9ODJTZnkWZY5eNWEDr1ccMwDzJwO
jKEZyMslVFJR2AExmL8mUt/R5iTIXHqofIMihDz09xhYHn2EuffSUBPVA11dm+wG
KPM5qmoVypoIZoyxiOQGrefVSXiYGoZRzkJHfWHukfrhgVmK7LuHe2Q+//mXzouy
E6dOCbmBQhE/ERkREntVcaXFYO/y7L+UGKcib60uPrzPbKIUBPVcILaGrFgv2Bax
TLLNlS0onUJEOZel1HokorIrTpFCbFnap5GlrjloQkYf1LbZzjxXENBZiTs3BNsl
fpZ+aa5oHpmqnlpa0YJIJMWf4kreaPWlu1T5L1ZUemvfzzU48litQr/Rc9FG4A0J
P0RurkBI2KsH6KG1/+A4hvALqjdbraRyJLFztAm9AocONCBLTwLVFhcCAYP7vY15
99Gz4RP0tUv+F7ljs8XcjaB5eIVCQIIbJ7dQB5EaHibmAtKDp9Fw6uaYH0hicP1A
dN/MphbyOo6ZsTcaDDHliqxoHwQYlVXo2pjqaAuvJ5VOU2u2bTciSOHcoJTdkVWr
rXimDDoTg5jFO3RokBO/yU+9hbPzRt16D0nrJ8vZmEZWoEZgv30zA5eqQr2p8DJe
Wy19Ir3Ul154a5maVa77IBY/ZwGhBUsA6D0rrpf16K+5KfdeYLQyoA+2oHRYWF2s
aPAidtWiX/aK5zeo2b8gng1xw+rpPH6+WYUGeJd5Sv6maaI+s23/aLwbV6hUEnOX
qwyPildlxZ9s8usAgMKxGS7qnsUMI8zwLuK4XjpDezLNmbo65PsyJT7seQU76Fbg
KX61N+2tGyanE1QjfiHCvW0koqFwURfLjoiPXXMubYReCAu55W2Z25fhCoYgVyYr
yptWrosFO/RxrPQi1j22Ru3n26asKAIVhPknOzGMbKZ7VJ8wuGsAUfp89rGxfuX6
5GDXasctxLVvm8kEujePVvl39D7sGq5e22iocLW724rbCDK8VFLM1umbrKyKThUf
xCvp55NTk39Kx5Jx3ubKiv7NU3w65POdBYductTZXd0S34lGreCSynzT2iQCeW9j
MIscCBZutDkWzSLmrCNEc3a1MwOc3krTJ4b/0N08jELri7NOkB7xk021PhKG3tRl
Oe5ifxYT5r8UYETstj+sVoaVt/+/TDSUZbXs9mc1eLqd1Atga2JY/ZCNVbyrEaT4
BlP5FYEIdLHzWV76fM1A/55GS6lDlTLQKKVXNUOQTsEpH6GpQxKCFjI1JHlG0P/W
Ra2P81mtEqTZPFwefQLKZzf8W65wT3ZTHopOwglZT/r7ZC3dSuj+8I5ZA6Q0SuzF
iJUSbTzKgONcXJmfwDjkq4JsFIpvSq2ZZ1j3ea0lEnhbEAZh9VxDBYXJnWdDt29D
lC1X6CBg0Yr7F8GLLuvkg5Iyiu1ONVTN2XMFUIy8zYcdsN5hbqf5w1Ch3MOUL3oc
vf6gpbWK9XJdN9ZpMtLVJy/hmvQoSiN4AhYTfJW0oZzCjqLZiov+bcdjR9xuQ9Mn
Ql8CiKU8zcdQl7sLNXp+HO+E62/L9/6ikysYMsqN3QN60AlaVrMaoPAB8lrrTQep
iwRP7BnJSKhLiDwg/1avygX864OPOny0/vjRHfF7Qwkb8m2cSXprxlONPDyZ//bP
jeRhtJGUiw5gWx6Nib+PGjNaBVxcTCP+hOYVLdzF0KNopRqXWHDLHkqtSsKdx1mZ
EZNnk/QsmwOj8xpmnATPah6MsDGQt5WARJI1Em0eML3JEWmNXIxHTogEFzi1DAra
XtpZrurTeiH2FBQKW2GPyStGXA5bJcG3i+LD47DxJ8K8GR9MRF9md8ZUVzvkCAax
WuQVoblOx0mUEdXsqKAvEEz2+28CmKpH/5EMTKMBmI7pbTehy7G2eFhS494ZmGCG
ugFEKLjZTKoitBuMs8I5eIk4QWhDSlD8fCwCT3kKiKP6ABaSii50ca9ikKKu+5Im
uvMX8P9/szoqK4fSVDzC66ee9XM/dE7nUHuCtPTMai1NWgwKwiTohLkey+eA92Ug
ibAOQLNKclMp4e+7/C2Hse9gKIWpBtGIgWHrKY30uvAsMcs4L5vT0xR5AsZUoUB6
aY+5FDqF158Or/IaQAW399XAdMqsr0rtSMFmVCIEipLsGNnNAVMv+vNxDDOo/rzG
1/MwzMEB5tgs27iV29sf7c4DfnNxclUmKDyNaRsuj0dfNBvmoNcrtyTSaiFWDoW4
A5i+L1IDUWkfTElgfZ67IzqQJL8IdHO/z34rsHc9XnBQhMJRVzScma+PjEUfRohK
V808vW4CntjuG1482olv4JKH1DlY0xvkglzCUznQKzM4g/OEc6+4xHvd41h38uWW
LilIjeB5rv3cpM17mpqoxZJi/vJlwQOI9Wr5u+cxC9J6B6utCyKdw50535kdtmin
Fw1ZC6fp82YR2gCh9tB5TuCkEfhmGT6LUjfWIAMwLMLQWiYhQRbYzocTG5X8kx1P
JZIuSuUMtVylhk04ENJMbJ/AcQqGJ6DGwzxcDUT0Mzo7FN2o7Kax2tGWhhUrL1At
xqfwWAIbkBlk+vz6j7A+XcGotiKbKGauCZfm1UsFwGeicqVOdUn1t5YWrSA/wPVY
lyq4zf63UNyN+J3XLs7JAXei7uAzkOey3JSheNGa5EBwheFV2NqQ2do1hxqbM6uI
SCQsWj4pCxAGlO0jv2Ta8X8ObVyJB5pSg3rPmUbzuw8RMRr96DXLkjiwDpp3MXgn
KHbrLQBlUjrdJ2Sfkf6kV6Ckguevgoa6GS9H4IbXDzaGuqZk562fYz1tuHiuGV9X
zqr30P/zKA3VWt5oeFIVM3HgnJhgb5/CxcNttLnaATTMDj4OuMUz7MLgAEcYDnIO
3oDG/JNozQDV5eVKvxBqzT0MjSJUVrDeCrW4Kof/v0HBLxzM5YV7DLdHOHrlBzZG
PqTuZszcWHcLqy3Qpw7ZmePdHVAHEe2MzHE16zohmo6ByUxMzHh0T/tJk58AzGgf
qTOEwfbYsXr51PEmXTOOIHDAsdkTfC7npTurPIDn6+sjGljwOOHMYSJNWqGr6Lou
M8n21DHUrgh1SV5QloAl4nnnBGDBekrbZIM224f1KR8Yi+VKw162IWmekWPCppEz
Ce2iEPH6x8cddLIUczUvVRRHrWieuNq1cHX2J3tgXIeqphF4GdyfCj8oyyDX2c2n
+fRZF0M+l+CEzULqEEpkL6DMwnveGhYhn9fvou8uFiaSeQMLQq6RvvYJOqTzFRsB
Yqy7N/DJrrOJnYmkKS5JxRLXrdnlm3EzDSEr97WjjYxwrfrtApnnGipRCMX6Uxtq
o2K5YybXeQiXKk1H3y4M+jy6zrUKjTHMS3gM7ZpI/OideFu05SGPnNwD7+4k7dQe
qVIlN2lf7+UkR8vWOWD1v9Yksxnmt2TTyV7zDw7OhWEhT2y1YA1IPXFWtKFYtL8W
/jWc0rRJ1v4t7VnfLBHyCG0BBnQ2UFl+1eesl4ivvshaBnbkWW/F9hAdFV9TRkI7
6QC8OgeDRCX8lb+tuZe3Uwh6GPEX+JRjQWMvliznVDPOeONLain03MxIj2TDLcFi
n0Q9ewY2YbfwzJyCzp84hGPLC4Dv1T+HubUjjkYfM1AbraaeJ0OlqAG9ZfT7dtu0
6cVc2BVj8dsk+r5T5Rr9B6g/I/MLUErrU5hjrXhe+I2Rc6yF6HNWiPkYkT6ANTJA
bNfIVXAsHtdzhpTVdFPRsK699gWlHNmrSuPN7AQpXWtYhIsolAmIsBlTXbXa0uW7
KuX+Volgd6J053XNNf6Bsz1OtObo8vR6ZByfU9QymHDsfJADdzhXbMXaOn6fF19j
JJ7wIjmFK6OEzpOi3KQNHrtIcrzTWHhK+bDGbv0GfoTpKkM7XzdM2/c5OfODibZx
ri45Z43ih+vz7LG4Bfyuw1pIuZdSfG4DHeT+uTsUdPtX8U+cHdS+RnLuuFDSNHq4
IqGQe9ddFuFMYZb57+AncFSuyMhvbLRZSfJ86qGnMKHMac0yvulXDhtvrBmverdC
F0zKiuZIILa/6PtSNTni/IP94CElietwZGCefW1X3LaoQ/uhvX+e6d0YNLUwtgfS
tC03crYjvJfwNAJypXJv3GiDVjJg5ibKMsU3IyJFR4YT481B6luIhr3GW24YCpJt
hpy07bdhk3cYV70FQtsQMyAyE781NJ89H9EJT2sBbs3EgcOdwY3c3Xdzj0dI63/g
Wq57GeF3m57OqsWE4TQ/PfmOgNdu5lFUwaDwGRWtcX9YJIvv5uxAAcoCixrFSEDw
pN3ubVQU3KOJcJQozTALga6CjU63LrBOmYWgsGLO9Qr71ZEASsUPFf36MluEEkGU
4KkCYqFZ8Nlkpq9rR9+KY8pCJvHtMNaKLTZij1acWQ3FXC20VlzWshtegqccf3en
tcDUZHBWIXuEcxo3wVcKwlpv341l/BdTDJV2wulh8UdfbNlWKqbDzKgenPhkmM0d
4JvRAqm+HVOlk14RLXCvcjW+4p4eIvfSw87hFhMTIV8QPCVWmvIZqjbQcuL1ww/q
FAjqhgx4ILDYOeoRE2pqR5eYtDdZhOl2eJ2kP/3t64Ww59/ivgTdVZOgjpkeWuvM
JEmOpqSD5dlY8xH5k1UVUR0Kbzw6glbnmAEaZmtl/ZU+BIsjUK5ZFBp5x1NciNbv
XfHAj+0J23f2V6mgsINFsoXU3saGnkwburgvLqEKSpDQDYlQsYHTuyhMmPgp9f2B
Eum392SGxNzJS2YDNIxa6OQZwmorpkqVecqDUe38E5YUl4BUqK6/RXlNpzf4jK1W
wY4s0AO0wAIZipnbIas2VvHrdLYn+4gtvfBgnbJ3OO7MjtRMYYA46U/LtAoxhO/W
EiuWEmzMBXsZUeDoo/X8oFu1jXDlJrESm1c7aihXesCwfgW9biO/H2h2bldNDIwT
vlHKVEY00os/yDo0YkXrxBp+WRCWK99d0XvgRtOZiCRlfgoPDH8oWUbu71eZvXNK
4hUfrtcXuELAecJAerJpa218VQUVWqQywgUfdWbj6iGv/9/tS7XwnrCbp+94bKF6
D8SaRacAvNygOBbRy4pPRtoqiD+VWtvm9ZLMep6CNncVHv+ZMM85Tf2TlFkKgJf2
737YMDOI1MsbVu6XwE0ubRJbMLi4gWt5RkU9y78KKNjfy71E+Gl51oHiUT+0N3Ua
5JMwkne5S2b8bqz4Unuo0RaESCfBvFT/i6/hAznct5IPmQz0wnnGLoAsd2DVBi8X
p8ZIP3Ee+Dt9rLdWyHKORn9jf3PzxL7pQlAK20KKAHoLLTzOTROaaJcWIq+2f96x
kKDsxJbOtvVRj+BRR0SBHzuUqiX1bOVMQ4KWPRac4xTViKjAVApVtBz0/4sTZuE4
0/7OX6Aa4f5rJyRgFcaW2jb8doP2Vao1T+RmmCNuTIZ7rneddZT23FTur6/bs9jR
Zm84rZzxbkZqX8/RnujYIFh4DfnQOdjTGqPrYHRWkz3eCYer4CldRaNHhcrjpMwH
fJef/+P6uVZUB7luNB2uAsVXJxxVR8nDXegcMQbS4kNlu/b5tvVBNIOltxyiD7IY
t3QkJJe9b5fi8xzqXjeZarBfPj9JtsLdsF6t2FkERqMtHrRKwELMPD5yFwD+PSJs
e1u9jpjofFoyniHzFd38BYDDeAKc1VV7ychZqplJCGiFc0jeLwnObG3jiIghtzI5
JYTtqt+rKzIz8G+dvEg628odweL1j4Ypyd1zXNELJsjsNEJAAE09lQDxWIKEPLhj
SAsAkkB+DAOjBYkpU09004Z9os5l4p/7nQIYr6V1jMDMmKIJNhBMf9EmSvQoR/bb
wkjSL3N590aWYzg/5Cc/8iHE9O/XwrJcrPY9I07BWXYAVFPiZw7eUIUee0T9gCIt
4ufDtV/G+jWaEyCR/KNZDBsaR0ebhVXjCkINy4zGM+jUq5BJ10lZ0guIJ6zFAOE3
QZLc0uqV9VHlrFkqzew9p7ydCKjLrMYoS5WXDeBLG/ejUPsviqhZMITGE/tnkPyq
CMgdIWyBkuS/OWCun09BkJysPeTbzR2ab+4EAu0XIACMGph8IbM2+jiATIHsScWR
jhSRiwVmpxp8HXmam1T8/Emh13jQ6FxZtsZNZh44552DWtMub6JcJS81VyYb0cZs
Bny5yG5/vNwoxAD/Zcap1KXBVkqvTV1mhF8OdcdyzzAyRcMGUfUeprz/h62ni28O
Q36g0smeM15qBqxakIat9lUaObQRPURNMgJKp0uDdL/kBch99rudomgPTiC3pxk1
XxnP/gEM68QQ97DN6/u3G+ihWuRpDZawx/CPN6IQ+s753GpVtfMpMCNQ/p6PZ5RR
Ly1qL/wTDQN16tp+IjeznpN0AkHBEdyaWEeTkSIgxtNIu6U3D3ZLiaUELRfXHg/n
neFNXF2uLDC5kdYSoei28HwGHeCC/vB9EXabHRP1K5uflhC/UKCLdJsSZaKf+XW1
sj7fVIkIx3t5C0ZHwHItOIob4sAh/dqws5Z5X+TaaDyUciOrYApDjUeg8fH6K02M
ptcKOM6VyYAAasMUV7uootjQpeKy8Gt6Lnr8SJy/YKm1Zj14vI9v+kuvr3GCViBR
FLG0E5vU3EvFHUBOlroGEBHmuE6gLZ1Ocq+GtiqPufYNAIjRZEqasVY7VveFy3oP
/fzFWDYm7beC2FKCub23gS00wywZJgYwJ1nfjFcH07DNtYHBMsehjwWfGLqy1OJL
5p57gwZbjxXYxB/7dKDWR3c27uORbmEwdvekLy2duOuLBl1weetRkEsmpjyeu9Oa
4UHW8GMi8IUs48r3YBo4G5e5heEXm6dXRZFP0yeykUvehbXJb6yq4PnvRZtUJYep
qhUtU72alwjE4Ruu91lCUoRb4MBchFjk1x1+VYehFFOOKqPKBjZCOCMmFcjx0RII
Rg4RVw4tkS/NsRnlh1WOD6q4thu6tVah+DaSG+AUT+07FsfXYCRQIOAmxs/Ze0nV
0QIAsPhGL8LYpgWV0hmN9NUJLMxVoMm7O9jpngC38Z4uis4fEhXbcyq9acWTjbis
AVWEexNHhA5lgNy6ut2P2yZ4mLf3YoVn+5B7B3DravNHuSAms2en2yJYZtge9bPy
ezK4vz50b+IGRqClXX5FQMTlp69T20keSiaLeYQFo5uo9X+m4267/qsEFB0Na+M6
XfUEmBXh8dTuRgQKR7nCT9QdiKG+EXd5+fomsP1ihcFinhTrnqpUWKzc9gRSHZm1
d+F3Y/Aku3CtVDbxfnz5hml7KkBMFzrRbNcI+CtutoGBJu+UH0m0U0VH7FeTNSLp
M3C7W//1jQ/whfi2IB0J3nRbb9174GIyjW1vYjA3jVrVbArmOCFwNJ6rKpAtt0gp
G6EFdCr2n7fb/bx2mblmKMQYVdY8AuZVxo/oyGDBdjEKNN4YMKUw6snL29AtzsB/
+5AYtJkxlktLP3xja0xh5dbdJ/768TKfTubyOQm++FeWZhvRQLs/p/fhlEj/a2N+
L0fensp16oCBxN1uoGuKuqN3H849k2uTUO4b84GClAPfqyWajW3Xza7XwWQKQKrF
/KtKsUVtYC7ZFXP84nmC6+uIfqCQD3yVty+p8zGmxFn2yDA8fUgEMC7/fweSMwI5
IIikjXVBxIYLw3OizkejRWoOCILNt75VZR8aPMH74XWaBi0DysiV+S/pdm0JRyZr
Ehbo5VEgKUHTZubnRD+AcCizmKpkIgE1uQWVSsjgNHFttN7UAbJN80Zy+jLjleL9
k2YAC+I1RMnEFD1Ja5dkxexL1RrLL6nHp0AJ/bF83i3LM34K7bbeUjKfYagaXv00
MznEIesoSAMUlQW3JLvtphsZFdizvtaTcd7fM/ekbFc16Q3fhY3UbP24u2boM3bj
CYa+n+rugqPazFbH1WMRXxJLTPuYjdeGNxfU7Ci3pyZZU5CNm6PhALcB877BRmb9
o8AATDJj4tYBqQwPBCLy7hDXm+PHT4i+3NjdrrgniLL3QmSr3cX8KHFG2FHQVS1g
Bf/nMe9X4zlKlK35K1sNavRAmHKjilexE9/f2dz0Aqi1EipTiydj4ZiFNuZB/1Sf
rUcuDI4UUkSEgZX26iBWJlTEz8jngLyBjuta3BSuCsHbWaygvsGoltpWivBAct3u
cJqZYV9hJ5mnTROAQvDJjo3V225eYdtnJrLPga3wrfRX8+zB07PnxmJAM2tnTX37
HBbOvsHkeFOKFBFlT8sVGwDCLMoumruHX9DVJ13M/tphqdtoqKMx3BmUJXNcS3rZ
ja0V0H12V/Nea7KBoQz2Q7/poyej5KO7mPhT7WlrYQ9S4Zoa6FD3GXXdkudfbaZa
q9QNnlQC2An5WMuHi9Rp7G5gkwg00wxwKSs5C/NERqWXKU9YYTgBumLYzemwmP9P
Z/xBDmxJfT7CoLbbjAP7kt9rd2QHgpFB/Sl26LT6gW7IoemyjgUncG0imeD7iZGx
8KTcGHrtvhtUsxOiOl+k1xXvD8wmP/A2O2G7Ehkk+yp876GYG6ueGjLxJbu+xkJO
ETBCiDVA3sKr82AMHRw8LopUEie+h8ZKzhwAGBZxvOA0Q1RIJm49PJqJu/hTbkkp
GLYqeLgbD9t9VFmJopFJVO4LIKIbZmJXbo1vmwYWLokhLsXh28jVBFIMEwtgzddZ
GxASoT9ztnpJjAvnqYWSAzqpfrUWPc+8RaPzeUBbP7Sy0Z+HLTNE2HQnMpGwOWIu
V4QTy/VSx3hnF9P+P/5EkyX/S9c1jJUhWZKLmpGy4O8FCaApKOiUGsstb9o4/4iJ
3kaKd1xqNhOknRbB3h8Iu63UuVSe/OlLdO4g5GmvxAHiwtYE6QFI1JK1hO6Xce7l
XZ4f3tnFywt5DeH6W8cBDsFhAQOnJKdKiZxpaiVgtJGAN2ED9O+xehKJ3MzG2j3p
07uZGySEVLbJBcRK0Dfq2F1tblKhZxd8Cwki8Eiu4cpbUibVDQ4R1anJV0YcVKSp
Ut+SfYCc265ObvLtIefIPjxu/9LC4otj1uCuJ9y34aheBVRhfLum92RMDTLVFlDF
MfMzxuOn0vfFmVW88Ph39emDiPXXL/GFBK6bZwfgwsAWs6d7nwiSpj1J7YTQzLIN
Ztuf92rqMJZVfQMGuGHXLsfeRSAkRF4yDhujz3nzlUlnij7+jJZylnEdkakXeZF8
+wT/9iCYCDoSLgE9TTcAijVjgw663E2lR4tlOjNo2kePfGGsDau0pH/B5+7PlmJJ
QV5D//O7kClZTUYxcJh6dlHa2Yz+bdu4dBIch+2BHwo0t9fIogBZDuer2Ah0c8VY
dJygjJgidYQC+zdIpr4FWMNHExgnk58Katft/T9veCYt9Wdjv6xMQl66FFdv+1EE
WhIYgVaX8T9I4bB0HgCrzXzDjmsI/1R344pWXHR2IvoJZad0DSNoH0V81BgzIe4I
BmhmNFNVvhL94mqItia8u4Fs7PKtc3cOFBL2vrNQbd09T6MaPKuJTAPgWcZjXrso
fik6kvJD6i4nnw8yP/qXMtUxpT0i9+KHtiNGD9IistTPhzQWCb4yJLCSmow/J1f9
ByVkF0ohpCdOytrfxp3Iq+7kOtKtrLcbYx7vIpyOx6YiRtEKJtepBPGJPo5AFTtC
CYch9hdY/SIHxG/Avb0goDuvIdp2UGRYvUpZA2U7BHAi2XpuaqdXQWSakiW1gM4E
NWuolkDK8wIZimfIowdnte5DV6znDJEQX6eUH6r3y7KCukNSmgJVq6sC8VTu0NEI
NenmEr4ic2ERjTymPzEzWpzYueMr91LC4pTzum2Av2M5qitQwOmgSXEI2bzvA91x
9XcmNRaE6MAw84FDqyny7SkRENefN1ttTXLV1jHG25acXJewJ70S/geLz1SMqkTe
wvpBPWEGP9yhs3yCSL2cSPqfZOJWutXtZZ6rWH0jGsbP4Tf8Mp5H7SAh8kXRhHAz
HxSJWVu6Q2j3wCnGRkNVy6Mo6et4aN70AdgrWqaB40pFHtGdL08/OSaH9QfAM1tG
xc/ZG/OBl9ufkVPlbBtzAx3dP9ZU+lrqF8xJM0qrUP0oCy/U/dlzBD7HHl2FZmyl
JIK64Ls/SmgDiY5cdrIE4owdykjQyYA72ZkiyffH1+uJtm9mBm7Nrk+08kChgvX6
3AaPepW85TVsgbG5rJ28w6pe1EV6GDN6WHcU76uczF+yuPB0Eiey09LH0UXc1veG
ks9wf4UJjvrRhMrzy/nhupZAife6K8ua/+sZWR3Obr1SYF/I7aOlX8NM+Ev0HwWt
svfnSq7VBUdVdvQsGN8xxRXMO88n6KyftCTTGbv5nl11T3kXBfeJo8LtRrTBa+/O
OvkGoAtQlhRttAvYfg1xu7WYJQ4e6xEvtw2WYDG2/p0YR4clzIYHdVmMfP0M5s/h
7dbXqCnumzNfk7SLRdAVgG23lvOQBNOrIXEORaCqqvOfaQPaMM7czzbM5YfbbNcA
4J0zNKPJeqnZzMC+AbS3DWl1ti0GyjDJ/cHCgi8jmOnCMHRKQFUryL48LQTYH9WD
w32O0Z86020VvDIhG1X0hSVtk2jRotswYa5OMehs1GjGxDLbZsu5Nw8bt7ngsEd8
dj3RDCcseiygFacnmYfc42mFVaCb7pkAWnhz9ir50j6jDFaFc9HyRn5mqDEPKo0N
ofY8omUnFqiW6yOt/3tusdUyEjq7XiIukskNafIKstsJ677hHysc1kWc4K5btWBL
zrtxAFadbGYBjTwC+h3y0DaX6k/PqR+FGhLv0yzraTNsiDVWfjuxyUmnmRJ9C2YG
qu1XwpcVJdo5/kElFwioVGFeJlv8VuCEn4Qfq+lbtHQoWckrORSlStQy2eD4+cQA
BgneJ0zgXfMOEvH+j/hfNk0qSq3tTXY8bA1Nmn8RPgZ73dMy8dCOhZWEeLLBFr6u
ifncCvvlZLshhH4u3BvX0Q9dj16DY2bLpmkjH4o0Depf5x/hSo7W+fpCymmH4d+v
wuewhqEohRe65tq0M6ecG2F21+lSF0lMNSmWDg/OL7JrQPjiPbb1wUY1jAPh33NS
C6rvGpzD5nfdg0dFKpH5D58l9V1w0sF41xJBVEGKWvhb6wS6pZH0TO9b5Zpw3rFA
i5Sumz48vWJUAOgHzvMCoaQr20r37s1EVb1zwz2M9UbBVfUGIEq1rrSnSAep/e0b
ajVc5ZF73DgujwFL9XtOPTIaL7VtGsCHQaG/DKz/NLDp32RIu6yVsM0hkwrSvDmx
L008OKe14hdSYD5FscEDSSoHPpSyelKwqKQlRgSYAkcMabFmnOeOkpYC0XfFB0YA
vA5sIGjLIiBhVTiJ/Y4JNw0OYXdv28ya99qQ5IdhifMDRZMumjLXzkFTrTDW0DCt
KMPO5pnIwYbrLco7TYhLChKtAcZ5aZYUJzQtZQsNqol8IyGYBKD/HVYSV548vg8X
vqPm/suhJigq2Fsfttd9uAODq48UWmSisOr/pCuU/dK0PxI5bisDY/C0N9WyYOC6
5irWnrgh7n4LTdDkJFf20fbqkRBxqn6MxV3GXio/mzv99FRhvpqs1fj59/lycO0n
EvN4mg8rrTq5i8WSptSyP713XiiVIOtxM+MvneGo72xXNButGUXeQnMBcnVRleeN
doafCP7TcLD9XZv4FRfYd2N0Jgb3ywt5yZbDHh1N5GFRNlnIs4YdrWPg/YcCe8rE
KU6G3QXdiTjNEoTF5FdoT6Nfve+ZxlE5RpWwU/xCKrkpfH5jW4KB+dV5362kH9yU
XUKcMLTgARDYJqEDqKkVIQZFQrALCZtnQov2laDmc6RyRLPUhPPxOEGi2K+pQf/3
vDZB9bheK4uhRz8eEvLx2MbbTUuwqZH3PqNli7PGHT9ISJoghI52foyvIQRuWYFb
dzyTZ1B1OzxLbE5A3xzUAsdBOKieokERcmHtz1BFWfOekAfZA5Sp7j4NQJORs7RG
50f706S98en3Sc72Gdgrc5kehD9kgzzC9snHBGuTw0BmCoWbGRAXGtG4VqVBy/Ng
05+/ZLoqpX1/ykkY1vyCfdnYN4z9rv4ZmAzeN6l6K0nEctPTBAU+T7mio9jwyokj
FBHcP1ePjvjGPTNrJsFlQOfKp3aEMFYPw672lXcCp9tPabuE0k3RnQ53WiICrzcD
FTedccx1YBQiOmAt6Yy3607ZlTQlh1CfV5hQ/Cous6jD7KvUlYogLa55f2DNdxuV
EuqIFWUmBzOg9B3ZdgfWtORhR9yWFgJIClW7NIirf6bR1ENpstRJ1RXNab+inqfY
WoCO/sz7SxoqmMzn0h8U9AVD7uu2eL7OPriDkA8W7RtiIxItwu3rWHATy4izo+kq
rqnLRHuiwlHngPnIwplzCAxLzDf1yafgXjjg0KJUEXtaRiIuMJMqW0uU1XqWT4gJ
S0Brm1WvlE2BA0QYKTQ/zPcTNxeLJWeqCrsZjXJ4xEuougrNrqpNgJ2QFrJ+/9nY
FyTBdrvwuip26OlRo7DGNafXrkdNxuZALL4rsjmhFHa+KMXGICRYApTD2eFgwhUw
OQWWPGR15eevNA1m2F+mrniMjIuvrjPQihsd/NUuGfZXFDcjdESdQW2W6zuIhv/g
FcnpuoRT/TN4oBrsSdCsgydk1rSv2LznK2UdDwHSdM+74Sa1HHDZahWpO2wgdszL
h0P28802hmUzPDJ0RPjPNsnnhEvyI5YRxQdR+C/pnciQV8nzv7lTzVQ18hNKBZrq
0XjEMuHZhWNM7thcGH4DoYinm98n0NK0BGIrlY3xISHnBVC4NGwVakUET1In9aN8
QvdzKCeKo1HqD9SwHPlNvW4B+YZaeW+Y+t6E72cromUrR2p9nt5Y7ooid0OWXUhH
OMqGMXjnypxM4O9ln3lqSK9lW3QMqUxaPuf9iVt/bmP3SVmLMCOXLqT/0slYuvOg
cQhuKF7TIxodQXQ9McwIgp5Qlc/EbS8DneijyNGp0ZnU6/VOZ+CMkPYRvKWEz8un
tm/6DwwJ6a73f8D4OjoB5+7BV4snOHAuX4FMDxy+sUHhwSvsrM1q22cIfD46EVoB
OFp42+m3k/IZUYPCVSKBViDLoP/Ko8P8oMNRJYBTSkqv0Hdt0Q+KMPSg/v9ftk+c
+aiw0sjZa+PvXnCybhwH0hlkBpKB8gWjmFuWaHzZxBmaK6EYGAMeKruBc4Xbca/J
HK24UvrdBrVJ8odOM2adXuj9FZJcfAzJlmkFXlcgkKoLYQ56sTBq2/JMwJ+JG+a3
N68NQPJC/NuvD/johZkhAnLiSu0xdSoa0FZSGRogVy7R0BQpnm/lZpCfPUV+bZPF
0Lr+0lxxOGIlWpIh/3oRPesDeAjSKPE2hySuZYHCsfp9dTsHNxCA6+q9jXXz04tJ
YN22A6ByWPp4qEODYuqihqCWllQz4rcxKh5RRNSF2WrRdhUCn7XzxBdXWXEIfCDH
EPTzl2MQ1rXEESZV7x9T2RNAOpH7XxuewPuxB9a/0XvBdDzEnxcFdfhuGZ/DR+Te
tMpxCLSRxg7yu8RnzwCcED73c0Uqy87e6TYznSZ4T9INaEBuTvgB2sjGBZMlTdA5
FtICwtiK5hhQtePaKpRl292RHHOh37puqkFt41FWAv8aD9anfNTn42V/XGHLu6gE
KAULBDmtNEplP4IFonkboImGkx4JY0UNKbuJQ2BmXSkXmZKZC+JmoqpQmg0NqgZJ
kCSSlBeZh8aYga6Sg1fcWUTQNpyAvkkHllaty4P9gtbmgw/G5hepu6Z3CcJwPY9t
I+2XwabPyqyZ+lIBnfaVARSCdWiXWMBpn4uv6xI9chE9jTP+3LkBNfGtuM6Q+XdH
5VI4qK5Lx5n/a/ulw3gp/jwwifusLNPuY8mVrT/joHY+8bse0k+NdUDkHx5RDXBg
FAK+xstBloNWlQqze0osmvcdK7N62VVf52L2hImaEQ1/TJw+01Q1pUD3zXEY5Iv1
wBtmhnXXhu2Z3shaaK+UY3sAKSmt7CP6Gi7V86J7lb6lHgTlfvRK3ktTe3oF2zuM
Sw5w4HQmIuTwbrmn6tlTWUf/I+qlB/uUgHw0D5lwL+EI/Usxn0drkuNWjSOMWFIA
7u0XrnrfyvK6d/Kb9foHf6p3E26tJFoYDx8sU0MoYHErsuO6VSsoxu0wtKziIipt
jLmEEU95iGVhF6AFr9v3gtSFd+waukDhJWYbUwKL4Z77YC+ElCkIW2xEOvol3TCH
YyO0M5mjpHnT4B8wluTg03TY6ASnnsiFwYvurIIxqrMbyCA9bCf5VHDM5gYOwEaE
v+6tJCwCBP2v4tGtKKCKuefDC3aXY4EaOks2TvPr61Fho+iFPuca64G7157G57Jv
pJVU5zNXXovEHb167NaMNNpMMv6djMRx4kj7NLEgsNfW3ZuDkI+kb3yZQ++d04j9
fH955jamrC8NTw0J9lHTCHKPXBghxuDC6SemXBUIv1yEy/UTu3jJDsSh4UHcLdA6
isQYqV0LMi0hB0P2EqU4iyGrCtJe1NxRrfWau1kjUHr80WZCMmw1HiSTESVY1AKc
eGXEPG/cBKTC8Me18G5pufN6F4cNoD9LBocE9VRPI5ucm+GMNaQlXJmOAHa08daK
q0ETMVum44foHuEZeReju27iHdl3ulCJAiHSa5GGIVJKht8NCHwzDwWLPO82Yfsr
D0/4zJxK1C49TRZwHrMNve2Wg+ghpa7y9f0un7Obgqh0dA2WxTeu7zP2dzC61yw6
RGo7GWf/G6MQ0P7+67BxgeaNs6VuwMX0W55/AZtDBJxLE+xpKo3holZcj19oatTr
j5TxO47DUUMQZjZTasz6d7T6yvSdWrpYgbwfIfQJ5zQan7zRzBIRrXyAz/bwnobQ
sm3K2QFZE4wEjDZ6iJmEE8InWpJdxhV4C8E3r+lLZhD//RTdYcuVEdGMZxrKEhOw
OEdJkADGLvbrQJGkPT2nlzdqfHpPb/3jcPRjIIxdqDtROyhG+TZFIPQZ12CByfW+
XNbBP9ePg189fftHNxjU5a0yEHCCUeVAw2DiEtjrdSOeh8saboV45WA1QUV5GEfl
e8/a4/1zbRPUNeZe691uiiX8gncgQfY1ei5o8I7vqvvOK0KVvapl3vqSz9QdWfjz
TPXJTuMPXfBsIykDrEutQSIxeHpvlY/bM0yLTGE1g6Rxc8xLD8j2RyGe8OHdexQ+
WfGTvVictko2kMBicNONdy3wXhKeJcEBB0BhR5oKC2C0UbmIWv7HtxGgmQva7lQ4
ojElSDUtbAoLit+3+hVk3ioWDo6zUCwIMURLLHdn3Br05/4/g1ZDMVsL8/H7zsFU
zABo6dv7PzuXtNE4ar5ErkS06WXxJImBOqAbymO2AP05NVrkioRsvcYVI97SYIwf
cDRtJYQtGI2tge9q1iAwkEths3SAxUgB1Zv0tInVjZCOufTNmHnKLLYxk/7wxs+9
fjEOlC+SVsy5hwF7SKL7T/kn/tcZ0xzdrIjHvgmNYlEn23jmro/SXo0EUUnb+POw
R/rbXAv04tDAVdyuIz5ngbh/N2TiEgYL+rqYcjOa4N+kpK6Z0KNNTrmQdbjpEJsV
wA9V8+Rfh8OxQ1nPKgf4CQRHirqh+ASv0WAkBVKnxlhjzeDrvd80qk9OvcJaGSTD
6HMqCITz2cz+C+kFwrdi55kpB0KiMxIiql2LR/nvsagYiV4bkW/5C61N8zp9B228
DwhNthSb/Szz3EcJkobjknqaPQ7bqQ3NXbXszMaCxIY4J4tL5+cBaUbXSq73WKXN
nnR9WwXyUc577Z5PC8s38FRhQfvRCp78MMOynhUNPh2L/UHALyabodzGI39/DehT
hVZ33LmM3ub8RrhvWx03+K4Gs2LswzA362GtNzAj0SLHiIXzzevWC/kROJsS4W21
7cip6P/FlhA8vxSCPHJEBIsjopWMm/5MDaT8/3kGeV7AJoHu/0LfYVUYvVLdEdoB
orTjJEnEXi4Aga0ovFRBJSO5BMuqhIUBZDIPly9NDyhKB+1/isaJ9qddwemI8XVK
I0svzKK1i4fFiKc+yhRHAZ29xrsfVpvKK52ZG0o1aw80vOM5IkOdR0X2RVoZIMjG
r/hDEmNFUAXgoekwigMc8xK94rXzK2YaxYpL8/64eoINAfWjwE+1v4cn9iiztbQA
SJaL4mcmxUmk6TA8r67n22OPtYXC8P8+VeRHtcxhaXdJP6bC5tdd3ZuuUlUKdFar
FcmSusq47oI2E9MpZlDWmwFJeZeGau0sLVJA3Dsi1tG/2mz7qXJ7ysel9FgA3tp9
ZlWk4tv5n3pL10ledoeFxR461XQD+kQuI2pKwLqDFSKl0PmcXbDYjCka8gYQST1K
DF2yMLcC1q38P8t2k8MTBiiA9ut/wFN4JsR25DRuRC1BvcQCP2X0OoeeYSp7kEja
sZFhZgoqe+6qhmX+QYTxAMg1s0KEzCMkF+BlX3+cd5LHlVnHTqcJu5dBasU5t5u9
AHsjI14kFdvRq6brTwJFN+lrRdfH01U9D3fpOwUuoosnR6vriBN1O+5jnx/JwC/9
+EMmwc3hbADj2irBN87qmnxIB8tKpzfNrblSoUFEdw6MRTOT5s5IpgKMWX6ddmwl
842gYbxBr3taLR/U3s8QA7q3f98E+ePF4Fb7Sow2fpsdh8POf89UU1KenfEFEKFn
GuaJ55eF7sN9pZmWr86DXBIG15ZuerRmYtTaRTGdvu92NDMtDlgPJ3X2bUJBxYGL
9m7I6N5QY+fjsNc/dQnJ2b/nd41CZhq0/bFWGLEj3JBVNNaiFAX4612wo+XWjBGW
X07SpFe7lM6U9unJaPKyKfIg1d9bd52RrdRnBh9GdPqVIMrW7/pUoOUt/N/x/DWr
ZxM4GPMkbxJUtczpq6M3bsFAhiXzgJHz/yl0crJgRF++y7X73rutozn4lODDafmf
tYPBsfjWC4xr2yePPtZ1uE/XrJ+vGoSFHj9Ga9/MS7kn09sxjjLgslIzXhRay1lL
Pr7/+HsNUleqqUwgRb9yBAMPgi/viHqaFFIhjj8JSzIqU4CNiLi7Vl/6xaVJN5CZ
86W5DVPRmnMek2C6+Q9zC39VR/NjctlK3/yCW0ZFQTHTeck7u+qOOx5kjfKrWKFc
GauiaqMirSI1QXg6Cx+cLUXjzgEhOC2Mh+7IDo3nXhQDEBYfB4amexsYMyojD+z4
1x/+s3ML20pDhYaW3zmfCr86f6oEHp+NUI8+NR4jThOUd5AQZ2+YeNaKxNkIZIN2
TH3CrnLSoHSp5Bp8kTMAwDP/eJxYN00rsdFssUNE1FwALjrOPqYceleEzZx/XnTV
YF4Xn5r54OqL7kesdq4ng9DyCj1TMfAo+evNE+9kU2MxSqtpQJWrszG+gHm5K879
Og+jvllykgTSBAcFJJ3yhmNyg068nPT4VXQI4mnwS5l5TuSx4whb69I3fwmPjUVN
0AtdXe7LduEvrmmvWxyj0+ucZ22IOp9YiNuTIoTpjHaUi38Hxkb3jEOG0hXHyFAj
QCDESz/zLhBPUY2x+qvQWKYQUqRPISuO5GYeidPam1NLHL2Q+entEX8Gc+qhHoai
1BOcCrCHZQIqesZzWgvaOXYyCtjfnNCvd6BD0CyJKxWxJNagzr6G3o77E0CEkW/3
EYW+aEV00W2kutNqRSnHQtptP8hmIvmRzVHVOrHg7VmHoVGqDqvHF9f/RlqOgsRt
HF/f5XBHJelbPmmvFBFt+bef84+6mfJ+kE8uSjDXnz1OqtWJEN4gQR1KcDUJf2Lx
tXJz0U3JWu59941ibGVti8SkX6JyW7QSNZtfBkeYh5mS+Vzz6l0HfJBANSmu+1HO
D5odkYi3QoKSI+S1G9o4CgMkm/J/5Ql7drvB+H+QYJDTtiNKgtUTOlS+CP3n2TsD
cAMNX2nZkG0anHBs6HS0FeI3DL7Sk9GSXM+MXyvo2IXeT6p4Xa1kuu5AJDj1Xlqe
V/CNkvFkR7XKI1QvEZtZavuPdPI9FCr3qn4pHDxXpon9OeQBeDdFpyHY3PiaAp9b
pOAEQF+3sqT0OtIYgWj6aimia/3o+kHMjUbJcCVVJHMoucXC7XxnjWVFfa+6MmEi
FGDFcLUXYByDFJWg4DJ17Cx9OQHoWpYCQQQDhiR2JqnyiFLJVukAJqV0YBXnQ++S
1W3jS2JtZGJ6AianpsBFsjL7c3oVqkUXLwHnGk5whRtiOCTaU7hXVuAjI7fi+YdX
2A/JFvroKTePHQS2lsmIiByGnySj0o2R9d+p1NvELQTIUEa2e/SqDTEXTw+flqsH
dKnoDS7eBmw40qqud5OacTt4L3V3/qmsu7HslG04wGP89EUQ/bmM9OYwMrVn/FpA
1svujv+Asm6VQEy6PQHT7vgN+y3ITivFNbhDetUjgUWt3iOqy8uAxKwKsvN+F0q8
xWSKdo2GEhKlhJksU62EdAbQpYlVD1onS8PlDz67M54FYVb44h0UWnDwFAok9xTW
jb7/uegOPV1S8gJ+yqBca51nkSSzEHj8LM1cLI7ZBZlJZpbRBVaHos0ZnsKoRcHX
lTAK26zMYdEa62ocsmPpBa8HEUbcxr4tnTwj5debjelBuKH90elOihqeZ7p/gqSK
J9iwf/QF34wZTb7zbbUhrj4uYY3sQWSnXnGVVHSan8i0I3XQaNVv9MbZXiaVHEAw
SVAqcl20M1haZEI6X8tTb2a0yj3+puqMpM3EHSmKQZvCOXzo5cjgid4bvZjfvBg8
xegt6BHVwJ+uwH3XFNMzziO82LvGoYylyXyvl/BqF9hs0Fu24BrcN32Gh3eSohM4
1ZzLfc3Z/nwgQEGapo6oC1c7m5taCyACFQphZ122XV21y8siX+qPeK37RRbXdG62
dDX0Dgnw172K9w5b6c4HkPdgZyqEeH43dMLTYeOLXS2rdXP9cm21A99yE4i3GY9b
RBien9lAxZPyxeiiWRokWNB+V5j3Kj6pMd6YI2bl8dHIoLiX1MNoEWMH20cUDcXv
mkfTNqh92FqXWNYUH2+vpkAkl7NJQ4H+dDrtB/7Quuff/S5C/ecGyLqs1gbJph3h
9pDAcK/wg6RuimErzXPbsKqyHy1+QlFZeWSPgYgjFL7zblFkmaGlF7btEwMkYG19
jNc3flASZo3j/hDeglVikxenOIC1M7+XX98idj1/CBEHIFjYtqs1xLx7LCZv4UQG
R6xarpoBQ/WipGMSvXumo8hfAzXGTddgsJXUqaPTlQDOf+sZrUWZJNxokkGc9ar3
q1L1SspnhOw+nAbe+RyFia2pgc1QttAjdOx0oE5xB9wvpoYS1+k6kAthLqfXbkV0
PGd8OiudN4g3kvXxfC6vZGHu5+Xoxj2Zpq1kvAlfSn4aeJ+McxFa6sBMTEjxoUZD
wrwL7dpsIUmgKpegtyXpyMABHTDnnnQLKGp6W8swuPfEPqjbTWIlADGCIHRSCXOz
oMDf0SbF4DOUvmnGAtWlR7atU3sX6pNM9uzY55+B8mOB9WlaGbycL3z0a5mGureI
JpQb7M8oSWk3VOyEgL3HdQv0JHwIedh5G/fq/UsZTgB5PIt7Ox1KxOeLl6I5LplV
rUK0NrpzT+3QBSXLxMrc2Q4UYk9asZZzuJGIEc7NnBcOFuXXN6tu76e1HVXZ+uI6
M0pRsW/hXA56mFBDbh91fzImt5q7rpOPLYLZyCQvtprRY/0oEghB5TY4rd9TZm/e
M9q4/UjjRV7/ABjWC/mLMTxxZ+TVMnOdq5jrvepS6uK3TSaKh3DPGItdjRyGQKAW
A04KDzrRFkwr4ux9IUCYnklAzh5neImdJps+PbdhkyfXyxVs1+SmPod+vSRSYeNi
fUwFH3cJF7a5377UAP5uvT3oF/qDXQG0LHzXhAtzuEuRvd/Fl44b6v7HEWtVxs2M
NFMxUQiw37+ZIzOrcYrKlRqr1fAscieFO8NkPGzyg79D5xBwJwDrQyIUdZs9yi72
qL7r+m298N8HlLgB879RthtaH+5Mvl0KLiAMqbIXnewLlMXcRYqy1G1Fxe7WM78B
NbwN02eYmU+6E4VXdw4r2I7yxYaIAGrXZ7PmNh1AfssfTEPzPIj/mgobCfriP/AO
S83wIC0vcXi6MXTHBICc7S4DwV+xuLTDPS5Vfm2c7awMvofKkBn3Okwz5ov+fUG7
wfAEvxDbkmqpvK/JVypQ2l6UdQCIextTi0GwtqsmGMOCKzaBw/oo4tX3HdC4i6HH
KE5rHrIa/zWg/MXRATcNRiLlXqMhXYV+b8nedZhHVPO+UOYHzU9ZmvDoadYRgTG/
`protect END_PROTECTED
