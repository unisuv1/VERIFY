`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LARkf+7wAREOjKkP/rldyAJCR4mhk4KM9E3QNTyQ63WgxtUlQ5oG62a65j/4RsvB
4OtPUJt+zBvzvCBq5rbQ1ueLfC/X0n18964Q4KQIL9PB3dI+V7g9TWZVOgGZY+9X
jehBckavY0NVzeZKIATeUc+owrCJnVXD+YsIAxdGYpnvbN7h5ElkwFbBJ4NJh3nS
LV/4zxRSbBjj9gi7uHjmKclxCeJGW4SE9w525Yb2x+dsH5VqV54mry52BLtTK4Gk
U82H0G+NWOgkmR5VvEbmCZts7LImK9x7Eex7g8H1bGqG8IIKBcRf4xlIbO0MsZTE
vMGRxIKM5oemnifmRevG6T4ymp2dGGsJBVSWLt60hGhXS4I6oXYnXzg0WFpGknH+
1IRLnto4W8LcgLg+uTc0450BKn+wFXXlr/Q3jGsraeQCrAijnaH1SqDqnSLHKpOf
nNduZ+Kcn+1DDYm4aOMqOrtGoEbhxWYe/zeI9NE1F1BHzwKvluQ1/yZtKaAO7h7d
Odh6vKAyWh4djiZRWAAE+rskq6kQeD83UYGMcGPSSMqudoCPGwLZ8TNsta8zp9Tj
zj+0sAAJjsoAiZlDOAptRY3mavoIzfYfu9YIh7S1MODzsE717wggI+iu1BL6I4Py
U9LPmbmP6HgflW7mUNZ1cMbVjW7J25HyDytPiJQlje6GcUVb3mYvFj8eSB0DMIYD
2A8kbFXJvJrJhCS4KXD4bCnQHnXxDgYvn2wYSs9BhTyFY+LZTPFS9gtI62PE7tm2
MpmZtvEVchyExehB1QtZoLcuzIW2E/ruuTa0XOwOzdyU7ssyAiVy5SS3pGgg5W07
PPF0THWafgvO5PQmjSwMPec7qoXyd6kICA00mQ1Q+FEzshB2kBlugrJHk7ZdOnfi
LkIu5p3MF1kbjEwij9jIUoFiEx7o3+nCmfLKgHAc0Uo66b5k+dwR/fr+uO2ZvlVl
H21Bfx1xLdl9AAOsjdO7w+wHsLs4/8jln7zd1ITBw1EqE6cxYTuLzG0BO6p7oorn
FhkS31MEo/riWvObkRPOiCcYcjVq0Ecfw+icDeIpdOvO9iUdKtnBVcjgwdC5Png4
E2dUe4HlP98trl16y8iEEGDTqXN7IEOqcOzd+R+Hfl6kWtI7ofbWxvtGLhSCGymI
quyge4XMqsLgtp5iw3vYM6PHRRDwKNFGZDpuRsf3o4kQ3tNlOYnRauR6nA//rYIe
5srYbq23vbBrlFsFzw1pFwbzouaX1/O6s/4dyjeKpD7dVv3zLno9tg/9NtCy0qUC
xBBpOU6I9yHXMU6mfAfT+jcI7iy5rxfJwjZL7JPU2nr9ZjbEPuGA7BHNOQ0EXd8w
doZjMWbvWEmVE5yj9jrrI/DZCBzXnYohDuvVvfJFXwVOLUZSJohzPp5Rdk78XxCD
j9sky+E7ycH8G3bJVsnKTgBTxtOyCNyb5g2w1LZs8Vg3AHR46t9XU3iObrQ/8pUs
x67nrBIHgMzcSBo8ejWf7jP2Ahk8yXKm4pQaBGbhWqpEahepOfip6YzpuFYrjFV/
DRGgFBO+UeJy+NyJDEPEtdezBflSvkIByPCFHlLJu2S/Hon1jWkwY7GW/O7W0V/N
qIc4A1R9/JxAKOqNEr/iozP5ZtTwEALRja2uYRVIImpawnRw7npQe4J5JQ5UbLK/
tj5lPANUA6KtU1QAu9YbEw4bFmMm2q47FIafiBy4h3j+WcGQtmuMIKFsj1TCCFbR
q9Gwm+u/PnAauFpoY0gXIS5Cf2DdVdMRfrGrgyI0ngW6Vv9eRocIVe6BMhq7jCWL
XhH/zjA1DjXA5dvp74YYPOdf/RvX4BtY3JslAqsXhW8N+OKo0t3hxD9d+3+vnJWk
WO25grvKeuDkQBrP6IRIvDgTk8jQmLvu1KG98hR6/ezKtJLa5AQW1VeUVakTE/JK
4Wvv7KveZvf130Ze/kFRUCAHnZxCIgjuXrg9YHqmkt/VDWP9hJSYKyM+mLFWLsTZ
G5pvRKworUyh5jbLlKvGTp2G5zjtVh1WvUeDXtEYc0g0ZG/PR7YNvgGNjKoORT6v
ua3gr0kxHjcjXO2+72SmvxtP9Ia0QKtB4D/jNIaIN3dwJUCEeB63YZ9Feglbx/Tp
ifrK9Vw0KHKtkj2xgKyxYoCq1l+xAeha/pCWpKOrYDMS0DvD2Cc6J+VS4E84aiif
m64LOqVFsWDTv9OI3pIgtHfEqDunsqO1jymgV2eaEmHpRwUSAC36Zx9Fdr9TP/KB
udu37MWLn29yjuAauGS7CP1C/zaU2cJ52YfyNCLlLqKGGOlVf2beaerDfGq59Avu
pHkbRxZjQio6KuYgjEdkqNtwlXXEVIHE0HE7VXVnEI4ZGbshH4/N7mqyzmWRmt3d
aCEvl9etyXlO5vCMrOgoxluVg8+09jnKSgN8mNOjTyLyNyl658yQFek2QdmowhZx
FCjJxBPFoOBx5BDM7NxPis7U8UDXe0V71jvP86JUgsq4UnD0xJmwMReX3JhDbZdr
KsUwnhIKSOaK2hX1H8/zIro3ZxIgy5IiN5Jx6I6rediKtpRZWmyyDkru3wg+I3Va
7k2oHs80tUYSpi9Upd4DTic7EzGhgiNfxFPHsaF2SQshjvOjcnTPKqOUJDaCOegg
g6nylyZ+PBRBAqx+H4rK4pgy2Va6jaChjwz+MVeAXc3q9kSYp2kNrNOQ7ebBbWms
3xSeOTiCagQc431zT58q3EYLf8j64FZYaO4/t9el7OsIW5hXUFv7voHlVr0/Ty13
xlqLydLtvreuLpmr/eHA2iBmFbR1NZ2rGBcHRBnQN/t/oEMaml+JfHl4lBvCrgvI
fE6IREdH7zKjyxCTFG7zAhWSqz6AW2M7h8L06XMnoszyAOmAinfHyx5I0XCaFWKx
ieDL8IHZoN0u53op/74/aLHvNok4ZA52gDdUlNmNvsOHnue/fIQww1/nTruVwdI+
7VtfLxmG/KxAyo8FiSgZy8RjoFCZUgcqRDz8E1pn8/qaErQMLa3yyelpi02WMMEa
mmEvUrd9VtdY9ByFUbuNK1wApf50e3jwxIauh09mEORSYx6jsNWsuBOvzMkYqn+M
cWI/Sn8b2EbCPwyYedWKgCR1vM27o3F0pJzxUTaeqwBy/a5rJi6lJ1wPINkEAL50
RpnbncfC59CJqtp+Nfya45w0oir1bVp371z5W0r/U32m1KVRuLWPl5o3dB1TUbis
wBW6x0TK3P/aHZRcQxOM+/dKHo+OuF04mZzO0gBsxlHTwjwc9bJf2f+e4ZdpL22z
9u3FNixbazY/j+uR/FPMPn0XIMiMtjcIsiG9dr5YjCV2UdpGUfiwJitevH9nJoX+
BaURiLL+wIVZzE1QTIxzFHiYwMZXUf8RUdD6L0tusuBl/IOaO37CnyDUEz7RKcrV
Ksm+Uc2jAzsPdSU87Fl6pWZhoTCUER+GHpAizpNyBjM/duCep+qaKWWob+64nrnz
0vepvotLSBRPv5S89I7wnP0Ymk5NRMiBU7GLuY+ZvvSIDflMZm86TX9qq4eYz+yC
9N1MQ0ySiWa/GXB3Tg4hzzxRWGts/yLad6GUi/2pmA0f3gjICYAinOYsP4d11r1J
N6q9S0eNTTdyVOcadI12FNF+U1Sj80wCWuHVb8g6n0T/rMa/IM3R0LzPxeW0wCuK
P4c149C2WCsYQEVN1JITTCWQfH/Q606PLxHJLul53r85kHeH8NOuBLz3ND+b+dNA
9vHg/9KPS9Fcth0obcNGLgJA87saeoTt6d2eaBKFALZtYMwLkH2wpn440yQL2GKe
YKhyh9N196/YjebBV8W49RzKo0GDO/d0+btcOHeaigjIjic2o1QkZpU0dy821Wnj
+8cGdtveicPvnxONA/z2BiV1rFkaXeAHNmvLMG0A/rzoLbPYOcq0id9h59mTAYSb
6LLHkMHUKc2vF2f+5TGcfKg6FqVtvLad7E9pbxKn5loxmv2NYC9bytobIjwkjw84
5qczi+B9gFKYwwkSmvp/8davv1M95a8zU6uq7ue8Qi4NZuCOPAgNqugEGnHv2xi/
utD4ZI5kvzZ8ThcMwtgVnfLVNHRR6qY9ZAyHs5GTX91drXZ4CIYpQy9vrRamEJbA
aDtr0uWAfPSi3V7xva1loXr3eFXGIvBfEpEwxtl/4OWvcMIh1f1LLb2RyKq5t2zc
PUZcdenhshaX1nc16Y7/sEhzdHwAMBfrTos15LkU6Os3o2SIG93kPwmf32EUAYZd
K6Z5Uc6IzS0cIFEtw7ywDZ2QSLbypkDVaR9iY/+W7udadcK2ReKqTUn0x62Mkjnd
KKcUr/n9iQ3YLrVRhXq1Yjpdz4DMeLP27HNNfM2NHpMTPQzXnW+tWMMzRo1r7AOT
zzl+8qwHotuTOuMKgmsEPAZFRit4rvUiHvLj2H/UqxuK+gJNgGS6dCy89nrlAQFe
VEzZO2x7qNzU3bLXVK/NkV9yIqwaAoQ2X1HAZ5gMLWKBFTSk5MgWDfspi4wnkdbl
pAgzjRYVz6JUU8RXADZCNFbJmbismsMhH9iVnLEtMPDZow79FEldBdG+zxUhCYJZ
LJxgV1DQm5JhNLdcNwRSM9R7fo7GXn7eyCIpAMmDoEW9GeMIY7R/XgIORoJGphH5
sT+NqIqqBcPCxBoVC9FGKAH1Qi475GBMrlAPMliCuAYMYdfLP8/NXgIzGO7eelKa
y/eF5XeFZDxtbyNmLaarCgycPhIltOGX0Q53i8yqRV3EWDYY3dFuJ5kqYCDkoU5G
C30FF+R1GUUPoQeQRNs0UliSi/B1uQBXEUqMtPCJXB99mdRta2U0th586eAabM0J
4Ql3vHQWYxTK9meHVZKdrvB6PoU9x4kHLRQetXfTA3xIBSOTxk/h+ISop+aZe+aI
QgIWxZjgJmrnlTDkjoBQkxAHApWT2Xeg3nBrNJIe1gqeDfOVM4Hv2qxWdnfM6x5V
257H1VvdyEb8SQzQ0dUOlCcK06yFxegBTm894x3et6CBt5+w4OVIpUudrhlf74Ni
7xjw7qz59YTUiWnAN2OZBpkXaDnGcshtrXeinxZtGUlvsFGpRz96MZxVqVTcDgYX
DSxUt4cCKTGSC6Tm3zMrsC1VUbLV+HFwKstA/Oy7k37xAOgEvpyIkImEY7DphgPt
8qcyy//xNwb64i5xlDXFabCyf0hNg0IY1PohNbMaylHTKFSxEv6hbfqFAcalXIEW
Rkr1qyi20rD5oBTgdAbEZmKCPWrNUPF0LGEkQiX4++0FBz9lyf1ULe/vR/N6BImo
CLva3CXvibWG3sA7gzVHyDhA8AQhAUQZAD9bO9TaAvaBwU9lOVClDcdEKSkHKbV3
T4EgsuQ6GRbHVZa+TBXp/x7RuQgRV5hSovxrl8P7cck/h/eZT9R8r8n1Qjq72Vwu
R9cMStUHC5+DLEuh1+HgvXg2iR8RXGt4aN6YBcRv8HC04uhRkwVzZ4jcIqatjQLV
lUuUIKO5Sy2qVO2jbyCXTvcdQdPLCemMcromL9zWdIZDZ2B2yNcg7CjPVrkLja6A
cgND7sOvkY4n0YsCuk52q3eQqHpW7AZf8UDbEjOPEpEukvHOxgGiEnJiWn7WZIc3
xqgapSAFPTeD21hRVTJZYEdizwj0QmRTg+UMzR564dk5DEmp1RN8KVgEfrXN9njK
B41krNskemGuFDIAen4LQsRuuV8HuaJBES5pXnRJYfktlgn+kQZKIrgKs0AOXlSR
aOKg5/BL17EcBAP5iRV9wDwx2uUacjFCWiaKptkhUdu4Nmuh/+P/3etxr8M+TQFO
hPOzYVfVNxG7/KmVcAnsm372vAQ57JhyaPnQi+n8rTktwBpbsY9TtEp0vcLQE1fV
qUIoR+6zBsvflH3pNNMBjWzgr7fdDXDm+TzMnEASaldTlbm40+07Ox+WZPco9Ps/
gD6Iv0ongSWwIsiAKSmsSIpjA40tV9QNrYyUw4YfvR8vbiAwV/r0CQo/jz3McCXk
DtSh2VwnKvUsdEKtgWZdIAjEvhdKmiFACxIvcLRU0awXfme2Y1MXYoUTHxsQgP2W
HDzvQHJhmWtCyZ8hERrXR93E9Jr1hp1dr4nILsQdRWdWJ9XyINbRbT4LUJ9wOzqI
Oi6vSvJ73XoUU/HZlU/7OeCvLsqdN3Fg+0KlnNXAJybLvnPnyPsNasUuqXECmE5q
yzcPk4VXCF1mhWXDrZrZG4Bo7ZqXdOURe1id+6gTgpgAIer3FjrPm89Os4AN3Nrj
tUF0cEVOYBZgoY6NFxH6SHxJPSF4XSzg2skEiIwSTLELEDjSfNZFkgNYLQgyd7jX
6dyGadaBTlGVHdkoZUMNxqxqJeIt6C8Uu6pULZyYKQP5ZLBpRwM2VAY5PJAcz58b
+FLv1TIf2TZBs9HJWiBuU8eGaGAcccK+XXaW5X0zV8W9wMPexzCWuB6qGkeQCVf3
dqMcQCe3G+SBw1chznjqw9SQ2SdGSkJsXQydB9Tofv4FY3XjfJh2CGj5QagZ9ad4
vX03EEw+RIb2lJRExKUQR4y1bSyf9cTXpgP5yOhOVaoR2cMZIcaIILga5EAK/OHd
LKfI+1W1skBIrhVcbDbKKZY/xRg0CnifvvpuSmSmiTVUOUpL+xZ/GhNRC7haB96w
W4FpqTjllcgRLYXN/G4SGRxiRE1wPb3+2551U4ZjKSW1SI7mtrJz0cY9ntGMRpBC
eVoFSJcGyG15zv7z9E0oObmSRXpskDpJPoyv7Fi8oAZRqNK3R9U1amVlKfYnn4fG
HS+B7Or7+TY8sl8uWb6eSh97OyRtQWMc2sC58EpdKY/tYyEP46QlJOgPW5nrZiZ4
Wt/9one4w2C8E1gnJKaAF8W615lkfCsOAOoeP0oy31fvDI60PARtv/nTJ56WiP3j
TQHv7ZRPZHZsNsS6ZoF7LdLrAceMtWMrE1aifijLGNVwGC+agzSS+kRgBaJivVJJ
VjRPghcDy1p/mbTqz5wYy2djdk7RBDpLfr6+LSG0L3vz90oK78pNnzmtmcBVsoZY
flPjUWKBpVBzHAfFCyswFf4QfEMp2VUFdor4etis0JV+gzWGeEIOYbPiNu4+YqWa
ZiztZMquUOZhd1PRAOFDHPB8knHP4moQpYPbqnsU9cdRhkIE8nbIMV6f5OniA3Wk
EDoycBxGFav/QEeOpfcE5o2Tyzqxcz6oXBoRciBl/RHxUGr6MTyGFH3M6TCFIwaC
t0Qfuja1ihm0K0i6RezrybtcDyYYU5HYAsnaimMri/h07aAD84fmH3FqDMn6OtWt
hpi6/PP/1wigQmI21FtwMH31qHw7GveOLyV3lBgIamXvEvOGPxf223J5fPWtScGl
f9q2GO8GIcaOoSDgyjhGGYZ23wN38qJcrVwaGv0rpWIMeM79P5qWG6zM2xxitWGv
seGWQlNKZA/sSyRJattmoyiQzB5HkVt+DpM7Psd68mnS+AVdqHLH8Ogv3IZ893Kq
bNtvJJtBvvvRbGkiNcZKrY+5M21R42241WoRk1M+jNdDhIAmv5pgH3oLbxkparDc
1iGv6GGwfSXaNS+9ra84ncrWOXGkXya8uKpE8l2DxYCoZNyT8rgrNsvPjwSTykYY
3wwW7IrWFLF2olcR6c3Jm8ZWpoDds8T74Vt83O3MQ0frZA/lvVsnC9pCKKd8Vi8m
1/gnIpiBofE6UBgACi7csu2SVZ/lH+Zi6aLRdsBK6WRxCno7vkYIjgEOPswgH+sn
qbBSHclfWgjaMiHT87f12mi3nuZdZ95yu/RIGYnX8X+wQGYRFF3W9PB5Vt5LV+wm
vfDP5HI0BU+ZQGnW5WA2QKg2aOpt94hcu6B943jNed1ZofjjJ9VxWqsumIt4DqdQ
buC9ukUyHSUJnetP2Y09BHe9C8l7PFe4rSHAK635LdGY+1+ORMAqwZyRIUiTOerF
dHrmi7la6ua/yk0hNcBUWn71ohkIyQ/8Ysfg75y/UrSJEpFxO9Jr6pIUkKJYVwkA
PUcQIC2lY9hbfQSasNQAj6NqTW/LhGAZsKHuKV8u37kElZhVelh+fOJ6X1fxIBKt
7SnMMckMA8oCgSqssfKVO1VI59Of3cksmr19l4Qn1Y2p+Xi9fn0LgNSDmYwAG2xL
bztcL9zfLrWztKu94gfUMmjpjJh3xnvdiRnyKo+qi88ArUAoAX/6L+isBL6zoIjx
y6s4H0WpkXCGeVlr8B6jm84Q2ymeA6ja8zWdi3+FtZCCuoUsb0eRD+Ywm5mkHBEo
Q2eUiBEYkjM97djOkjisdaRMUHKUYvD3Lad8wpvYYbwoKCncwv3MCK0xiULKtkca
8dDnn0s9hwHdeWhxT7dDct2gJJ+BgUNue126qs5sh8w7bFkPTqs6VHUP7DVfJDye
McyID9wcU8MSseYrEf8+94GCXKRPEnP4RET13V4Qcybc0LTUc+svrX6oGUkoNpVo
7Pg4q1llRSAVHlZ+7bRLVlPclA5VqYzkOy7XBwhk4y/IZhGzqgUj/o3Im37iVISC
WJdOewmzYjxfJ/DuGhWUHwZUECptR4OTrUljgffvBUsqtBhSSq2nnlWaLcHYgHov
FdT+SAt7lfjIf0GcwOdx1ri+a5e4Rjs92TqLkXDE9RVr8OtTeqvgXUxHghx511ZK
s7RvuDuIemYt/i2hxxWcCA12QukM72zYUEs9hqHG7U1Q5K5UcfCtkhiaxx0BFiO1
gYX/LWqYja080De2P7QgwQG6l2dHf674iRZgZIdmqiRLBd/YD6dW3hXPWEdPfD3y
McPiGSEGMPAm4YkFucjJM/sXKbQ0CHt35UGUJEujDBoG3PxFTs9fQ7Zls42vG8yx
9wafoDpT17WMTVUgQEEV4rNnuVsFohw+fuPP831VhyfT2F3cSDMU6mkR+F79oyXX
j4RVfj1OS30R9drZi3OqaWoHiggVCHItKAnDUdvEujA9GHscRMECnY5d0Mts79PD
/EahaAMPmfxSibgZsyH8VoFvje9WLuXEbqXQm3qw5dOynkHUpGDbggmFFaFBfve9
IvxAJ78qZQdDtyq9tbmgvxOGg5ycISkjYAMoMGZXj/uWYiRGYcNFkrqVhhuLZFfZ
v7Sryh5nvy0tXlA1KlILyEiEAJYKS0uJ83PwUfwGbrfupdy+PeYe/qMDzH/b/jk+
+o5xNghw9clak8bG6iTpVB3UEkblDdk1nANHaXY0aY/c1ujHGVxRQpTUu95+EGz9
rNajoS0qfJHNF9NpqsJqluzmYYaA+lEPwQgE+ApeTyUi24wRYwDeNaS5X7/375d5
AXnn1iR5hV72N4dkoMRh2xu2Gv5B8FcOuCZR/6SAdYAoLgPcMCaDWOJnfVj3xzIb
257k/xRJXc49ZvMzL3h7q0hNWVvIdm2ub35r/TKu8Ug4Rf9Tu8OnygPKRx5unEcl
mhKSxJkshcEhumWZoXNt+welmObR2IAAS7XbTp9pxNC9rgFr23ldnRGnQAcX4jsG
nfKhPy1GFJy2YVnNoMShE1u6c+XjYgL4OGIp3WZzjiWGen0xIvejdhyif2lCvDKL
N0qAtzXVQC9/CgXRDDiKIzkjJpxvxJtqsM8vMsaWIe305ROQ//W1Md/3h8TrKP3L
H5p8/if5yrmJnYVQ2UEjFG1F4CewfjJr/4z3CrTsD9fUfX/NVaeIN/1BdJKE5l+B
d8qSMJpuAQ7L78fi+J2FXzWtyU0W6fY53R0t+YhKvddquJ9h/Z0f1czHMa7TJ8F6
WRaJqwHAVCNv5UtwwLC3ZJGFDtjX5FVlQhHb7LpMlyx4s7DntBhqYiOi5fmY0cx4
JrZmkf4ksLMF1/GseEJVfveuHr1S8TSPiH8XU4gVu9x8vc7fO9HkxYAqhpXkCDBd
21VML6nKV4GtXv+Ifl2tkrrgIXliSWYmnDBmzBJqsDmLoqbMlqvri0e54tNibJ7A
4mF8djRL9fGx3cqZ4om7OaQgzNdAJoqezXCxgUEyruHzreh7Sdx99VuF/RkC3Nrr
YQRP1SfxUzExMf8wBes+s/dOC/NWbvfE0ygliBxUZkgzZs/1SHyneUiZ7MNopBmQ
pKq5psgDe5xEepEKkVOFhWY1XJhD1i8kHgwZz2rdO+RBeVqJjxSZ/XSbBmeBz6NW
6mNE0asAOS9mQMDT723JyFXA7E7M0w61fxfNmAvniJ8MCMrzHcVdblUVvrDuegX0
DPLHSUJviuBbzrG6oWIHeBzBEfphuT984GHFm6J6Et0XsDlpl06AFMbNtszdtxQh
ya4f8NVKh+9PMFjNXiS6RnMyKdPR++GLlbzB0dFmDk9ZoThVhI7scOYgKosqxgoi
o5v6DVcJgxa//G0cPsfXryNabU64EAMncPnnm5rAvNlp93aWDGDpfnskni6vWYY6
f0QtXm/yWoH8VWccqkk883VIkoE5QIFHp2dHC3WVW1Ch2ldW6zTuimfYlmv7jNhL
N9ZtjgKSlc4PEPhCRgtDmNpYfPiZvbbsWSyEHiEpsOBGz9OLroyKzCDFxF0ATmjp
rZtBjflBDPKc4zsRSNRMZy8YGrOKK2Axgqnp3DWjtgJc5Slx5SCahfeqo1Ba9lur
fMlu4THaA84xbpoez4xmk3atSQYEHaFkj5x8jpG+GLxu7OD8z41lUd4MdQvNdg0c
HtUCGn/y1kcCHilzHKq+JEKfifVNt9mAhIsic8iFIgKdXp8pj8BhJeU2aBM+aYCA
a3S5PYqY6j44GihdeEFvhSBK+C8dNXcr0Ogqxuycm7+7Zi7FKEUWbgdsglttrZnN
mRrcxB+hHWqmIUoUFvpEd6xVRsQ0RsV82I3Nw+C3uf2ysSb9cUMBcpQWnxatybxo
tz8JYZBgL+DV+vVtF6rVyVz7TPBlrliVYIojaeZoGsQ1RMXDTgWvr7tFjr5YK8hA
YW7qR5CbqBZwK489LipYX6+uvag70tTH7igN+YiHm5Jq4RIjkVpfpVN1IxZIWfnu
9HKzYWztoBXaR93XurE3bgutH3AXrkrxyUrN7PaY4g4Rpkvg72mSyqwmM8Ns3DOJ
wxpbXGDTnXmU2Gi/P8Qk54bo8fOwnOwATMZ8RrBcFPY5oQKTpY8OYLCxxE/0R81v
L7dUVTMqhHEctwXad5+JAQ8dgRsRI4nmaBl36czMV7+83Ye0Dv46Ate69YJ5SvtW
90DQhujmFQr2j++i2uOv7Fb9xIwx3+iIY97IHLTURJxjzKZ+PpWULUxmBarTqhaN
owGot54EX1MNNvrCIhIGnUMAVGgmVAOIRC4nst8OPI3YF+XHmVYoB21GdTSDjO0f
WgPutm7YfiA9ZKRepK331V4kct0XuZlK5+QRInLNOqtgdokaPUHXx9D5vn1mEbSA
HcUvRz+bUuOiX0m0UALH612ICzrC2U3dC56VsZ9X6uI7O8U9Mre/qZZt+GoTKa6w
gWiJVXOmj/WUUYutfcD5AP/3q/wqmfepVICEpZY2LXpwbYFPNJH5YiYg5RZkVPlg
qNZYCsCY4SWmg5YPAQJAhOjYB+5D5mENek7yb33WdtCUlXrm5UD9a0xQ0FCftwZO
GDHPQ0+tUmjTBrejG/OKgMd0WTzqNRqh5/oWRwK6TuuXhOguw3N6DDklvFb2MYQp
HC4oZK/XPOWraxBft/8aThdFpu7rU6VcpRsl5vDys9IDI7mVu/VzC7d9NVdZ9hat
7LTBCh/TjPGVRE7mGuiCu/orXG9GM/jXooquwlthqac5KbJ6YLUT70ZEu1A3NIsl
5TbKp8iTgtRCOqBZkt4pDDeqcYuI4N1zgoS2Qjsz4K3I5XTZ5MV2dwynS2xy7N2F
lRPS9fs4aC/4G4xCoX6N/XSCfHOen0VaOgdeNQOAxLdzPWZ6Bj+mQ2WxzCTxWxUL
h4lKFbOSSv649cCh6Rd7KPTas+GVBHcc49zxh6Sj1jDMthbWP4/3JqeUuIOa5DsZ
2lLi3F2/PNSg5eR1CD6xaYXI9mHM+9udpvsoUiGyUM09gUvAH2EYmr6w5gEVjgIa
6rVNNXp3ov8VE3D0FiRsPMYq783UZNqXz6jXySQBnD5f/CJjusGEaSAMbG+qTqXN
ykqOFuCZToLN+jCNg0aw8GIRxeeow4dqcVA2dSRODy3v4QvTmLaIjhtPz5iQtsUs
QW+EnVwp1pmYYxE1qeBEsJu8qarJ2DSHvHrRYNL1o5CWt6ne6yCj1C0VMR13cNjS
tHJuATChkxqEsBAAzga4eSb4E38UZA1DNCH2rAjUBmBA3EzPpQe0qHBXKiybFtKp
FVnJqn5uDCDl7sfgQNgOPWcV54iGYRmNM94fAfg5ivmlpF+HJMFKD5cO+klmS6dN
5SQvwyxxJEPLomBMLri4jqvs7qq1/9t8ThGfQ5PTXuvLUhRS9HOVAX8Zafc1oj6l
Pi8bOy93CQHVhkQLls0XVGA8tzcdyeRwqvC1z1avobovejN0X6NoAnBIklpcLXku
t7+w/Yku3YlGEBG2lqfFju2qrhxs7qk3xq0u6O3keXthxP6bVbRDFc168GFytAa9
us94QXlufBnywR0+vikSFVTTsHnUWzxMe+HiPtRSlgwg3o2yjtMiH1hRb7iz+Df9
nrGtRhSrlptH3y6C4IK5Fq3gxSWrKjMpTlHkGECVJDnTrdwxxfYNFCKXxqAQ6yLl
sAj1KI2aRCKtK0SZmiE29bgmf3UE9d7KpwJ/blvHNYSsq1/sp+6upRN+ohXniVIh
cOKLQUT8eT7/Pdd13ynDVZHx+ZVytddIjvbuhrnP2sagKgPDWdaDigYcnnjker6M
Yd08CRHss4kKdTRxLbvE3IrXWBncGFJ1KnYuF/cjEzYMvtDyHHaeG/2GePgiWoxb
6ex1D6Q3j3kIXrn7m4xmr7XtxkdTQF/k+9XezpO+SPiBSAOfW3XEOiCOEFesfWwm
HF5Tf85mhzzqLRwSyKbKfaWTVdpgo18IHXe7F4IutUPHuRN6Maq2neeV28KTjqaj
pYU6S2QGDuHbCGFimP9vlh4Ur5k5afbgI/dYJTRJnWLloiwyN8FJ5+1zPQY/qjS2
+n03NKhkvEbALEqA5rim5X0hBYvffUamtzm3fwf2A0ltTzOTraVRQ+3oboieFi3d
PlqEtNsCOYpRlRhaOxZGGjDHeSjXEiISKmbY7djSFB0+Ylkh+8rYGIhGX/bhtbns
YfeBslrke3Q41wLcsjNtDBEKXUPtRIrvxSg/H+TbHwwJvPuLWLcSjCcw8ZN7Lo19
BOBXscRz0m1AZzuTnYIwmLC1gN/LiM4Y3MIXKfZv9vjfLf69ncgzg8VlAwN6Carb
QMSQh1ue+NuPzMY9ulM60FbMBWKsQXhkwtWmpCGE5ulJFl118Cbo8PSPROtT9efr
`protect END_PROTECTED
