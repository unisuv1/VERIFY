`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
6a5LauLrZO7rUtgRaBCyLg6nDPvnVAk/pzKdfB9sgV0uqsgyWJOF6fUgq2KHWGiv
KFmvh3tNdXiKIKnDmG2ILQWIL6LgAB6m8ryy1KpX/tsibtVELK0liA5MsGIiUlYc
rDcaqUFDYAOdPIQpI53Gkj7C1+Co6Es8Xxr+Ud5ixalRj5r4E/8vceizjizhGSnp
BZWdfY8tcYn/umJt5rCXkq0nO9Fm4xfAwnaHDorMkenOAeo19lLYaJMFz1jsV6WE
gybdvfLXEvbv9TyhX/HUpNgJ/Dq1SvUvfmZwIvZpCZpYuT8m1HnBTYkqwdOoaShA
SvGjcxS2dAl7hgFXD/G9WuhHi6e0/KGIoj46/YUtwKHRIB7d59r57pUcOtNkk6fu
NTEYtkoIofgZytIo7NqgUlYvXXtXJPUYEqEFojO6exMo1uNuDlFJh+U0fqdfjIta
UKFYXIUKXJTiNxsd+10LUgXj1gaLefWrLWS+I58P/bzgNawDbIzpluTZDMCpc1+O
7jGRpBnH50eY7hPVG21KAZOgGC5tJ3n7QLLJjqdLjs28TVn2Pj0GHZI74ALyM1oT
w31iwID0RHYcufO9g7WTyFE8nRhH3XkW8fyKP0D3XCYiW6p8lLUbRRE6ru6a2fQu
+5bXhzl73xa58lqK29/6SeMlr7CcDrpUXulQ1BMEQfz49aQOvgPjEt7PJHK/cHJN
JIRBjtKMnmXx+uX5oj/7LWql6fnR/lU1TzQoMNzxrIuqSIGmTp/8ff6KKhCjVZdH
syGO0/O6ez7FVVIfVJyLIt5mmT465UCGcvi9NhHVkcyPXOXjgmvEz/hZncVaZkma
hIAWau8ZH9LkfXjAuIgC0LP9lc22PMj6ZvyzMgNttzf+n2j6131yBvWwj2Xo9SHs
Sz6mcGEKoh/gadQwrB/GyA8jjvBuRP7CxV0MJ5AB2Z2yZzsAK8Zt51xMOS1Ufpfn
Ay4AIUiZE5xdAmuBeJdKOuKnlxJJUQQPqzzjNHEQB4WvvKRrstfl4kUjTkLLPRiY
EcABnibzySSTRrTZqHBz6CZE4YwwOjsP89QiX3UGU6ACaBHsn6VDvTJ9C8X2eiZZ
Nmld0yCRNTuttAZzihWYvlVy63od0pQhuteE+odFxQvPW9nJ+oM9J73q8+FSFvfK
kzVU6A5CVxpUCWG4ZAf4ev36kb/lfLqdO+EA3BK0oZCuHMiO6IibkbV2R05RSMGv
8YtkdEP98D8UXKAvZ7FgpACQ22dKLiTW2kVo1hd4Mpifw2PiTr/5J9U/qDsW5cfO
be/eHcQrzQOoq7Do7FSGy2qIdEuH7pHDQFBBzFeRatDwMvwzFeDfjohjAStAr6nB
TXHaxGE9OkXsVQmxaV3vYicdZ/ozGj5JKqZUAaRylr/tS2+8c56SHjHJe9gRTUub
4WvhCl8/y7WPpQadmXlvbkDmWveC+Drj2MlBUmufzAygLsmoZ+RcE7cCVk/GrDar
6m4aTUIwIZITDuOi+v+VnxY6Fiqqydug53VFrPaeSHFO74sNu/aRaKQ/B6EQQvq4
bMCtCaLjwkM25NH1BCNm1XMKGcqjhrLocFGxLm4WG/gW083x04hOleZYKQAqtjG4
wEwz7W9Fftq4kW9kPYCPyuVigXdWMJnBvPBgP2e8REkhWW3659xEen5/fqi4MyT+
oHCVZxqeJ680Q84oTo3PB5rpJIW5z35U+THssLc3i/svkJtfxOKIViumCv/XK9IW
u0TjXI+6pOW6jL5wLOBGA5Z6dRVyTwqUoYts61miwACEoEA1RNGm88rlabPkCUDj
UvNF5N1qZ7fMxf+ZADfUky2F56bfXOj8/7WHHgUBNiekkakBUjlN0zoRmIJje8sN
0cJoV/hq27P1gCvEJ5dRHgwXSq/N+ZQ/+ZiwL1LhH3XalnzFoU+6jAwe2xNznDIJ
5z8owjepQDoLFwRFB1H4iSgepHGsUolPUjOWeD4BhJ3dokOLQ8LNq1rxtZiHFTjQ
Df3ueZz0zIf9+h96E8YfknTdTk/h8NHFsHgA0fXyETuRHaitH1J7C52y7NMk0NEq
vZhk+1bCNd7Fq77XEBSMkeNT82Bfy1HXDWwq2KZDV0OHU3UdZgQ8oPbjf00x+7Qm
87w9IUaWo+fc04nBeBYS1lbriQ3PEO9UdIDpO1SHwz/QOUusAEj/Jvc+VdRjiFs8
1xyDx5PfBZ7hzJGKkJSyGyg30xXw9O7u41OrvO9TrOyXBi+7gWyWwLghVrE7fl++
1CvVzQtD2CZWRUWdC2M7pcW0yspovU9GSrMSwyl36kRf7pOTVw+za2dB3UxZsWsg
IFr/UrXmzOT773JrrgC4veSBPnUJ3+0DyVs3kdreXMwQF8TvIQaWRKXt6Uj/g89M
WUc2BH22nA8Oc2qeEkMEMmxJuUcid5nWc4vstmk0fzsrrpxqDNxbHH9cOzOvgqqk
WCq9wNp+rPidBA8UJiEAnLPJgZtuTnLOIeMyDasE1Ygn9OtD9LlGt82HiXXxNtDi
8Nj9qqkQycN5YPv0Hlp1M3Ox5J5zrG/CyYX+aSmjCkQnfvGm3x1RthFrUfoeEQHW
rNbDE+jFmT+rTEJfxcYgo16lZDzS5EDJ9F2pAQUlkPUzaCMo/Ueg3+qFLa/4Kthg
wsxISLD8B3e2mGiW3HOiKQXXdaXV4yEa56H87HVpmEDeVovbkg9qu9m75Xzmciyd
n+LIfr/qgUMyy7+d9OGDUQli3nQdrUhuQmPmH8ar7IZqVVVRJRsrtzQsuE7WHqA1
qpoHzI7tZpYCMGgjmnbjzi7F/R2an9+3eLSUvq3nI7EuqHrtqgSVk5ZQlSvQFMqd
njPn5J58SlaZDfBSipzlk7Uc5qdQbqMEYQCzO9BAS0QzohhwCqdUu7uDre7ORvVD
Or+7qZoZL/gH5nRIv6p2/K8s1lTymE+QHBTui6AIe78F3Ef1EMYI4FaMEHlgzW15
edbpd88sIVCLe0h4ZNJ4H60Fvc1GdOKb20BNYJQ9qKMSucoIlOCX20mj/5+LFapq
WrIw5iObW15nKJsqJ8F5HtSr2+aWEpzM14QrIH1WafJdVw59gBxMo7FI4SvHl22H
6jY3s1+FxQurYODQ6sp71B+U2T2ad8Z8Wezz+/BHGbGFbKhE13VLxhwGdy/R7Ve7
lomhIXCrY/otcqv1nDsb/VRfovM+XDY83ySW3jpIMDdY0dnxjm9WQ4HEleAhi0ST
psjsUOjU3anDMSUqmSSrjdOk/o3rzOERlunafXDNW8rlpntz2u71vqzIJ2wc1OQO
MCy6hCf2sndin75WzZzValiyzD3fSroqsn/I/Qf8cZPXS8ftDdvqXkP5vFtiOsbB
d5PLo0d8xqEGLJ4xJQwRltbLMFHCaoJY0sDZUc0qLrGmh8+Y1JovkvftHIZsdA67
VwToS0hZgBnKstYHgdUTM2e9FscU8binkBpkL6JcEdekSQ4hwxZFAsnA3rQXdM5z
bYPHW8+oj9BojbQrTvnIvvpq4JoAF32YQMUHXb9xtSfKIjnPFbOo+j7vbt0bAPh0
T5w2ab0xlO74ECHB+/KWxcoEkLmJ4saGsEpmD8mIFp4paleF5MT+n7qSlcnQ8rw7
igEgFs7t7X9+DI/Z46nKGFDKq85M7PH3SSoWZVDD6GoVHNmmftsDuSGj7Az9Dd/m
XD3sxTybh34Qcc7JzR8Jxb7bEqSS8MLd9qRyM17XWSJpAIlAh0TWZ/NPxEwHL0rx
ylVH6WH5rNDBK0+OyEeRU1ax3Jt7cFlHa9gA9UxTRFVFE51WbEhT88EW7vZtO7xW
dk9tbdUVWao3BSescO7C+kbjg2mLlgsLHqa72TV3WuwvGkWmSd8bK+DbCK2QTGnt
wM8f2FU3vIpccYLBEaCG+97Lnoo8PljOrsHC4SEEdFT+PGt3NYAQTlTE0OpWEzHy
qPSv3Y4oKBIMfPgIhdaM+0TV6r+4rn31JkdUGo/OhqaATOdjIlAUTU1TY/r8O6Zh
OIn2yO3tZTQVEEB5meOCJ+UzKC88coQCs/kw8i5TiTYT1KK7fv92W2CCSyw8vj+c
eN/Ln5iLNhqotiMx0LiZrIx8fNVTmizULy9GVRrk2UsWFc3bv1RR7uLkbWm0yMR+
1NJe8/+ye5xL1i6NHZTW5ZWY+o/VZSGMZPrjGqE+I0O42MxOUrXwxzFIXou634qJ
UiOnSzkV7KfuwabCkqu7Dm4HIp4gvJwpZoo/4R7f1D67XbM+jlsrKb01elKHo6S7
MBoBKDfk8zkbpcqRfViMg0TUtJ9et/9GBxJkzSiQY0TQSKT+jZ8w0YkO5R6LsSuu
hZSuOmV3ESC/IAqIRwqDthzsaPRJDV0uuQ4GB3mwAYSnvCj5G9JHS+JQbp4GFRJi
dgjwsAqJjD2McaPlI70WzpuqYess1203/7n3mFpDsKRYivPkLhEXPrAl6vdIclWN
bW1aQgr/Ma0MFhGIuq7hTI1LCk6uwmTRhieY6t7sQreTuTmJgD3oN1HQXkmY0lRH
uXvb0H6cH1p15aejYmzHUMZdHF57h3gksAIdl65YygRKo94SitIrFKGmzcIZmQzx
i/NrMhg/R6AzaEaACKk7V0u1gIK8AIFFpGB3T6lJHY+kLSs30AUuulVTt0uKTzbb
O6qVJrvYzHYvnLiPmzY5k+2Y1mRUlh+4Af07EF1Id3u23Ihxc8roGP6vyhgkX5+s
4QuM3B25xBzubnPLBsuI0pSvjiZfwAuDfBnA9RggEcb5TYtKDICs0+1a7pBJLT6c
3HZtZeF0djfJB3KuGBxjNWDcbJc8OSVGd9JfTr1ei+6n9vzxbVKTd6fbTeg+MpZl
ZLtjF5dIN3gBTpgG0Js9dH6zeto0fUWQ3xu9tMGrd2eoiz2RyPv7h9BBcVXQY88r
hhkt9n9BTB6AmKI3sGCQx/C4vCZ4R8TKId1ybwPrY5qq1ZEOayWuShoTfj0SiRKV
nnehRqf1K+/G5kGu/5XoiOQDub4ZA5Fkt9zijcOnS/gY692tLef5tvmzYWUsqViY
yoXaZcI7819ASriHR2lZ5DovkHD1y/YGXR7a3a0pTWlctWtWbn40PYCR37+eVMW8
BgHfoyBAW4iz4yA55oXULZmWYnBrdwiDEdP5I5Y6HP2ciaCT50S5yB0KTp1jRGf5
A0e3oyFLPQLA6bQ/CCfKXlIAYfZUo2212trCsmVT5cLEitOzEiAENcDRq8JyLpS5
TZX5rpgEzf0lCEP7KdZ2VhNHZtVYIlrinGO0axaKP0JXRohC21+yeCwAXq7c8mYY
pnWtx6QL1bPmrY5zvQZmIpPFA0J1kIsKVSFwhr8nE2qfiz76Y2q0CRkSNuz4br0N
cstv3iZ8UUzSrO1el41T9LOMLLoixRF4jXJHkQaEfu058R3iIK3sVLAUU/pdjzgf
yitrwzgmmliA2hf++E2xJqEPAz6RsMrbx/DGnLKd4jbGh1am7Q5+3EBgXIEbXYqV
WPyRpSA9KjlAxwZ6ojk+Oumb0k2DaPI6SXQKkh46YESn4T3WixG/QqJpwdJcV4Pi
fOCUI8vMif/spTKqA4WGRgGKuTG7I1R/0TYQ5Ckv0YFQ3Mznnj3gtemKmzt17XBm
XhnXFXHd8tIJI0qeuEhQ1TNxOBE1YVyW4HLVe+RgdbpVtTrlSysR/FZdVvSu9BUd
5MeKs+Pyt2NphxhqOJqLFxbK+aDha0FibT9Qs+LA8sZzyuAciGmp40U3/lzalPeg
xnlUVtIDjYSjDZwlBkujWX0oRv6Mm2DK9AL37Uj9zTbQHFSd8Oc7oPaMiLskSr4m
3wHlI+wlOevycBdAz/PkeqsZbG6Te22maNBA8gkehGlFpWmn7c712W3ZXdBEI3wJ
8uFNK8RyrvqACJXvven61hsMgS2idhNsGBlWT1fIYe8FmOreovCR3UBdqVvv13bj
1OeWRd5bB2DaUu8NHlwY8UOZ3MXZfZbsr2d5QXcMwbnn+rfG4gIzRpzI3gSqmt4D
EppPXtPo5ff2tQ16342O2W+hdRFnROHpAwhDkI8fo3Kh7Kb/WXDaPMg4t828vRhJ
8jJFNCWU7Oj/4HR9lrpwfgFYh5lHKZaGAnudR6xE30xvWiIvzPhSuiOS9lUKSPse
XHyWu6zNzIYTtH8wcTLX1PAkteRguOdgnHxe+3761BV1GaTVWweRXyPG4rh4E+7f
d7l3DbWJXzRSjxSshurIQvMYr1UDjffu8DpxMIy7CyBMxQizqi0PmFlUQ42sKQwH
EMTDjCknzRSIgdjhLoVbgWoVeigNvos9h8hzNesY0t/DiNYKYts3IT2Vk5DN4U37
m/tTu3riFxQUzNlpAihaqUwnULcPKnIxB5A3XTmQYAYXJ4oMN4WS6EE1EO6CsEYx
9FUtBgyne5Lux+8numm8ySoy+SJAZlawnSfRaFxdxLupIf2I0DvVpyCBzWCN99BE
XHtFc16nCW5z+wdgCpOKDZFFdlrC3bqwk4HmqGRMw2ttnRI0DhUmrg/OVsAZsMOI
XhBLpZ+2lvixEmV3XU2XXRW6ASycXjPY6pJJJiaUe6qkMb2br5sjiuxpCx/Hcrrr
BUV+zqeCOV7u3WpYXT4Z1geKPSdLX3EHl4LK/fSGGmdamuWMGEln2JneAZGBb+OH
/DF+yLDvjO6ZGf/zLpuRgxJIxoGe/tH0TkGv+nGuHL06OyX4FVu3oFZ6erg12ZdV
zXfRMSP9TLXEjkqdwXWMTm0R9ksoPLucnAhC42WtLRXR9Y6o/PYL777P3g9saYJo
v59aFSg8rZp328VfIcQCA4ilw/TnlbK1g9qjlKQkrecpOBhIHeetho7FZtsMPUIp
fhFrdCPs9KeIdzACj/f0npbxFnAA9/3kDZ1OwRIOYdcQBb6X6KARNsWols46QdSG
WZBMNMdXXD8V5p3jbLzibkMA6nZr5AE+0bFGKTOPq6UrW2J1vq7AltvPK+KnvAe3
Z6p2mh9M+tn/mEyrf1xBjmJMnYA4n7Nj2rJCK67zOxjKnqVlxhR6OMG+rGrlcLZk
Euvg22WFKRpqUUYWJjoyjSH8XhgpUNeuJ+44HRJxVODzE8BZ3wid1h3u0zq4wyH0
f4ugQDeDv8yrod7HtSFcFZHy4h82Qn69RB5WW9Mhd6f55pTudBMUyafyIhqKZ6Bk
kKTKCPuLN5CL2GL8J8QsxDbXNQJOMbzzZDvP7ZKEDpk7q5cq9ibiTesP8/NGwZ4V
rtyfDUaG0NSSkIjrvbR4gxWhAfEg+z6VkZeSI+LyZzb410nbI7mgwiT+CjudMGQv
IdGORTq+nKIlKdy+xFShMFk0Gz3nOZm0/vUHe2mRc4F2kfIxdQ6SlHIoYAY0Ya9i
bGjKC7afxQvyV8WM4Cgitc8VJyJW3G8V7d/fIg5I7jUjoKuczaVpVEA30vX6QiSj
0BDzYXFMYMiJvUIv2Sl+0QOC1nD6D1FZnQF6IIoBPM/GDSVBmzi3XnE0cy/I4t3O
71AsAv0IwKbQ9E/2XPI1avFkMrdLDZs3bz+PHvT98KoQlnsC8mOq31dcZ0U8WlDx
ANKWa2UztATbZm3qY+C+yhVusLgecO7ptV9VjEbiPDlSqy/nUv7VtpAQR1xqriUX
Y49Xfw7rtkVnpCBbG5jaJwNSweylQehn3Nc/o/sMMduE0BB1mPI4kFOirXJ9+GsV
+q+4a1RJ9KSd+fY3pRXia52I2TBAVnsf3ArMgglUAVDnA6qU4PSBEpuiuhgz0Ix2
7RGQZwWdP/dGb1BeLW+e8IhzrerUN0YfmskJsT/EbuzL2DvzePjGv8f+HM1K9sbx
3e3xILdivjPyDH4OK1cNpv4n0hPUD7VAm8BfyCgGOyMql6qA9qgw61aCS+3/LMzd
nFd37PE5qc9ZIcvyzpo8j6gerJqRhI8ZhMMzgRfFOlX2aSiYZnxOs90YPOHlxfrv
zZvuD5TM4St3tJiKKJ2qnjd+uZOXMtagz7Tdh8oPcAkQ0UauqebiCW2HmyqoK3vx
XRSHkdoRlmiasfeqq3vzYYnU60yHD5tQABuwK0v+edIo5kWGqeK7vSAK4KswkKBF
aaGeurqp4MArPyC+b1+p1AvciAJfB+2yGotCDCmdL62HXlBhaJKbOljCaf+iDneC
4h7gy2lMkptqbRo+FhGuYMk0lInwT3nr2tqV5nznsw+OuJKGRDoStDrr4iZTo/Ww
KdGOWzjBrX+cgVJbfEb85JDUTbbzuid7mJ/djyYQzVH8Nk2ASa3SZSfBwURT6S+Y
9JxlXyQ9tD+Z+GK4DhPJPXNXq9o3ZuamI9j8W3sfLaHdQ7FwKOCf/NjGbfOtaN1g
e/87X2SCGZLGluQeLHNEouk0dewOWx6Qm7tQh+GOC9lUUKJMMRh6HUwRc9z2EOok
l4yMDNiPukz8RpyVDiLQltRiGKwFFXLSGfEJ9BkPmF5yIYG4mAuZpphZNyMBLBGO
x9Aj1r+EsrjF0wx5Wl9tZol2l4ULl8MYX5mFvhoHHmuYhFf0Ml8REiE7hbxWEgvX
uusl6nm5kuWJHV2K2dcAiYIkLIWYfTGgJr7+9nzZC2+9Fgf05jWueL9HL26gJ+LH
WhM6aFgfEvE2w4nEbbSApz1r6NLkOJTlXwgClwiHQIzUtYiLdU69SEssxoBvr0UZ
KnPAq9ci3sGE2Fxi46JSqkko28biJL/RgAv12pPKDFNZP92aLOn5cv7eGnUAAY5o
z7UbyFhnnZrcX6xQvRJZ8DGFNWDT9QBejLhoYz7xPGYckbTyb7x6P1HyZ2qFNXpw
EWX6un7mt54/a8O6+QWRVx5nLVUvvWv1oICnTmdhgEZwCF59QGGQ+TP7OhZaW5K8
Nl8pkhQHBN5Vctzte2CA2PJzj0nDxnZt0h6aI6PiSelUvY+P5mGfvvYgaimHamF0
jefObhgcAKzv8sw0EjaqkCCqdM9DQddU7TsQvGychZpjTbxMHNS1Eubchlz9sThi
2QSqMqPuV+GWS5AkrlqLxUOKpQJ2DR/1nxhAx9zgOPevzjqXBozs8V1TydSiq9Ob
7tPosNv7kuK7HI+qJydefTzVqynzeTTGCGfXxh3PXfR+CPBywq4KZ/H1x79K5SrW
g533nyBJPPXMJjBfNrOM+uQR1oaBS3vjDLcJrg2Ot0LkOjLlz2xe5nJIM+zGGwNo
Ho69X+bJyZM35/sZUjVUzrzkWNSD9ItpApccEFMgbdkDQbWv5Ub1/7/PLCkOQ34L
9T4LcXppUUHcDp4leXLRoHVOWLGrNXqvebbsoVLzca67CCTDp9bkOvkK1xgEN/H8
W+G+G7kfVFIenkwD8Ar+N+HdhT+gRWgY0bPsrjON+OWtwXcP3lPGNNjmYBUrrhsF
ZB6YzqmwJbKsd82DDTD4Ld4ho2Is4Jt9dGV1PPhYjC4nqylKyWLT29o8YklbI8sR
r+CmLgvK3k+zFWywSNfSuU7FVdb/6CBrK2Ev1IaCAMlahoehjNvnE8ntundywLUB
mrNJdY1Z0OiKFTWsvkITZQnhgEqUncy+k2gUby4k4p0wwzvUIPdywCERTzv1pCl5
Q6mld1YBvbBKg2raItHQJR5muOxvLCA5MV95tjDaOg3qxFBSGqLK3DsHJCKLftCb
KLislLnLBRaYlEr+/sSsfJTR2H1pqDeVzc25m2uZ6K8XLRDgIvlzGNHN1hWT285C
511MqHSFSjJWoA3bWeAdWVM31exiBVq6216YQANS4dugPnBOISchhy/u5m4vGJi9
iD9bkeqSECz3tgPUYEXWWb88eto3DH+N+3ENg3E/DJ7IlhAG+ZBnLle5aIfOPVzr
TsdodLz5KkqEpkOeaBFC0ylNxAWTVK6U68HhHU6q67tIzfNxXwVJBHS7ijH6HsY3
2vCvvZEj449PEqOduyLBBuyv05ISW6JEsRmv840sQCCoiqbRrzvg+mS/2UInNYUV
60DFUbk54AppJmR/QzlhJWtMUJiXKxlxodvsOwqAJoLT1rEQxMrm+eQhAolsmx75
t+tcUwJiX7P3LeCBdrn46HuKKEN9TxWKF6RD85v6JQ12eeOMNbsMOuZgha2dewaG
Fp7G/AenoFe+HCSM7wRiQmZh+w5XLOsXIvUQLDeOwo8yELbN2CgEXdpFWvfCmspf
RUMXuzX5vsNyIRqu5CVjLVoK7K1zRCkmV0Q6ft3bOGL+UPZnok7u9Oe5QbeWY2xf
XGWTbVzjNkkQLTPwWVGzGs8fS5pyx0Vky5q/OIZ65UP/XfCys7VGlpZJKkkPgRG3
fFvfOtiQBNzY0oyFsiHT+rvLu73plzD+oOb9gpFRNavAybj0eYEVqABkXHbgm2d6
X/B18lZOy36iEWbnOFemBEeILX4cvgmk3OYGbrkO97BUuJ0UYWXtHFu2kfFu4wKo
cV5ykTaAO0R9qj6ymQp6h13gvRslifKIyW+hyH2YZTzbnk3zlxFVu0iw35dwRLly
gisfFFw4wyj5176i+H1Y9wjXzfpECZs9ysK7KznY2OMVo4kP7Veqr/wsoS7XrELd
/PmOGFpE7nTEvmA5UDQ7mHFC9xBWlXQ59KJ53Nyp50fZNB8wXUQ5hZOKZ7sEcLT8
d9DcyhKlYhp80RDcLg6fUqbqE3Tyn7EfKBx+aEvVrK8jc4Kb4RRv5JFNiV9qqIMY
U/Egu4p1UhFU83YVIrooMVdIbWzUeSwMBk12wGW5qwrzjLiGy4mEziqWJGadm3ft
GcDsLfyDhdj4ciJeN+8kSgqSzdM9L1YGu1DSIrgasISpXt/PCApNm8PLyn6KoLhp
sZ1g0yCE7IMAW06X70Uo+osTiE64x8O4/yKguSdUwRgYH+DkM5wcxZ3O9sNIgVQ5
1tuMfufHLD0xQoLVUTImSd1hHp3xkCxFWzjSkpMCcXE95XgHBbYvf6InnjIJQEte
fT8elYiVKTHeP+UFz6qCfsrtRcyWnw27WH7uJjZnK9bm8CQsCWZhYhvUgHP8Eb00
TVBpCVXU/5vEtPLtcDpJepWpeSJsppVcKH0+H+7eYH6/+eLp9x9Bd91I/GWwTIOR
OYGMWqn9j1+622PyYrrIq2ciJkUuRm/bT7O93hvqUpQd2GrtFS9rBuMhseZ/Xz8b
zrYWwwijtdEmYayxuDetxP6ZPz5GSde7nnKE+qntjestqYyIwsVecrZq5ZLm4u4t
K3lDT//CSgHkBon0JMCEwqJItAIsrUxna7ZazXfgQaiVRq9F8HWMCWrLroPegLs5
5lW/h+moYzCqwLXZQMlw+UQzAqIkSM8THt8vntRI8WU3+GtYbjY1071V9CYxxcik
KRUfmnq5JhiR+EvInBasO8dTtqOsCjlegSdCqO+GnzAuFnLUVPRBf5nx46D20ETl
9qwHJBiYSaz64bDIgeYJiSPYpLwQzUDoqeTu1fIGy8iR6DyQI/6UzYQUpnOfwr74
uMzbL8BtG3F+dvk0XYH91P/1kC9ehmvkJvDr66ewXH+403VlMKe6RhEEh0tdAMfy
KlObU92gZniVxZidL2ku/1J1gTS4ZFKQk1/1i/uvlNjmZtDrgMnjsZlWjIXhIudV
+E72/Jp9KIpIkaAhBicPitJ8qzceNrvv5IDqz9AAGMM2MFgt9rxq6Zj9LtzvtqB2
VkjHbBbFZJrXBWmIZqQ3yfdNKu8JQC4ld3HGiZe/3pkJwiSMbAf++5JNdPJgI4zw
1m0XkdDmRCBH7EIz3pLYbKy+ULpNOd0KVTwjSIuH9ASrHIvObd0CHgGPZTphlZHk
OsQ8ulgsDpEX7luikUrHul+PbDSBnJ+9QcUrGB9RY2cvhwtsTU7zqbbySoK/PRIL
Wc+ZCEwWZFsiFbBU2hqJ3GCocoNVtaoPYMo4Fh+uavNFl2gFjCY3C+t2/YTuqPGu
DMR/m5gL256LQ8egJur1ee0gBEjP2AbcEk/g/o0sQ/wMeAF2MZyQ19ENyPweKMep
LKSTH18kJyuhVQtRLAeSBIZHlTcM2bJZeRtQ1FoktNSTD/P4Weqf8Y7lYQtF82H7
duv2yU0ES5PWGt5WORgA/vupDNYunCfyHP29sl34I3Z3ykdvLFKrguuuw/C/hXVZ
9T2tCSu/nYAR+ZiwEQSgErle7ccZk0Ubk0BsvINQ1KqKYECYsAsnDLXucNv7hG7g
N6Z+f6IoX17Ig9AEVfPXRvWfOOGKOyjUKuxX5y/ziI68hWKBEYRPD0fr7unAU7vh
FjiJYyt1LmWJ7VEaSnRwjdYxChAiv850Zjxv6/E/AHGlhBxcM90b6p+OSczCvAAk
o6NPvtowKsS6gS0ftPAsZkvI7zHPOZmAIlqcWm4/N/vHvgWCZhOQPyZDB7ZP+a8Q
4z5J46gXrnvIWI6KITtNkjJF6ZEUqnyiSRmL2kzJd45xR5W7HH1dNwz9FvGzJrOe
iHOyUxP5zPEiYGvuHa/C58uPgMiQX+qn5LVyqWVch/oC5JrI8B49LDPOLbiTPhYJ
ASwoXIvwo9EPa5Kko8YIhNNVCgxBRdlDgyIpE6kd2yQwYk15KDp1kyKaQMtlP8fc
9Wo9F/h/b/TZaYpUnKJYt7IR0h+OehtGKFUSU9PsRVhK7vardZcbA3H1KWDfHFDM
cMYlcwdAuO9xaciqWHlReqotJNQBr1TKyPczAn38tDv4Cdjg9FGRQNUcRT9qQLYm
jOLIXYcU1yoMjqtg2g0OBWKsv/xQn7/jTaUTFvDMYk9hXwph0+sRT9aego5FXnYX
jxopvGSIC6J4gSAeb9kl5dsju7w9ii5+fe5npynUL+4QIYrOGOyxAhr4w/CgyssQ
+2YEzYb17oIuy5s4MmolLPmqBCwHOAjA8S6Swyh/9b3YRcoB2z2DRKv5ZnDnkW/I
pI53L8Js1S10jpsr6wup3bQZ+mRguBqvBBb2i4gt9rsSrKlGfJQq1Jh2XOovvfi4
Z00fTB1iSBCfQmSNWN46V1/zuFrjMvK0Cdyy9nL7aoRFTFTBDx6OHukmvGEb58zQ
fwTLpvZwAZd8OTRijnWioc+m3r6XfK/33svB3TVZkHFnXka/QRkXBrzS8J9Fy4Bl
lpAKtgPUdJ8F3U8KHdIPFVdxpj7xS1gWHFYte+okXLsPEAmOTNawgOywDc7v8Vxf
GYjhhuJNrnzA7qr0L5bJIzRycRhZ1th0fzg5NM9YKbykVa1Wla+YedEfXBV68/FQ
sdzRUYpUiVqfulbinoAK4ASeICwc1IFdQJc+gHZ3pt31RHTQDM6mNzVw9ykJ+WIp
7OwSJmZHJu0zpuuZsqIiqwJlQTiHQLUzu94IZ6FWrErd8HdCrVaQa3YWYIj4f0BQ
dZ2u9HX1I0VhZr/RUj76XN7ttNB4/ozMVZOcZ/PcPMlOOv0OJXSCYhD6teNFTXCJ
zE7+L+nPfxnp48aUjPF4M8CFTdH/yPV/F/P6QPL+an1D+8vHjPJ1YF7xI/ytYETG
/Yja3kEPc2C7rR5BdFkzo4oiFVfi49AYXDvCvgOGkQ3WumhKGRkKiH/T9R9+q94X
jb0mhjb4nWEVPskwXMpwklxsxwKKLfdtl9V5jxBoYf5pZuHurRnEH8W9Up+6dB/q
P/aLqOp2ax58eRG4iq9f0FMqXpPrlqiXlxWn/4Hf6ORW6yi3fK5F9ndFtp3oDD5m
zVKAYestlqOl0zZ1tsJLNkQHzyubRlvKclPcT+fNI8C14m+FZbbryQYTr0XmpAlK
Yz4Jk93nxGb0qRcTJuiIS1gdDJ4iQ7b2TPzoAnJ+mOCGdEw+CLp+RDyTksFqT8YP
4fcRnN6pw5kTuQyFQm3c8WhFhl5COvmwTxfU78ki++SRzR0ongt3rF3bLKSCnmqz
C5OsUx23vhwvvMn2kVuNGjmp1KBmXKxtgsLDfvCskK7q/JV5sc/khwQzh9pZclKU
yPv1KFAYzeETIMJg93xoxYA9eaATpjZMaZOe4THGNqwSo4lBRLgOq2pqIZqKE+91
8Yl2RR1YVe3JIj2iGXjGtbkAaNoah46Q6p3sRoWzlx9+h9nMJTzM12BQBir7yzPB
7vtLZewtvwRdErV46B4iZu4/4GOpWdjnlB8IGolfHMbdGpXdPlti2P7zNczWbmAa
+fIbBrie6CcTGa5Qi6b0KZ8W9z1lFHi2Kot1o/ZIco1o5wf0jvi71OcDyDpL+Jsb
EPAOXFg0hJ6uLppodeDQ0l/kBflskVvkOs/ING3D/dbi8XEDvwY3bhtR7uVebRGe
W3nqrAE3dobpsAc1JVj+r+XL83qSP9ZyQP74JEE6wnPD5K2zSqhS3cBRPCAqbCah
ha+QRjeAtZm+klumtG92dhjXR7M0TDxVYtu6/bfqirA4I6VITDW5vHe0evmNajEG
n+RzWueSsLspB+XnTopdCwn6y924DzfgkcmYdZvazPVkx5m2j8PBSAJM8CtjHm4R
JIJOIC9SgCh2+oBN8TSJpvi/mX1G1wWDXLFcVZQw/fGtjxVKtObXS91q3+YVSg44
ST64VWIIGElL/zGB/mZGoJibSrQDDnhYg7RjObia8hKqxkWGjTDv6hC3Da4IRNib
OcjOSKUzIeEeosBbfXhNIsqiVkjo3EMChotoFEy7UmZD8Pm8zYQ/zK4eaCVZNuer
ZZG92Vk7+a6P2aPITssVTGtJAiwqXAGflpWnjpYIdWFDTCSSFrQxQs/fFp7jI8w2
egCxqEJSEl8eNrm6ITgWACImE9qfTYV/Obyk3XrZt3vTgbUEy67h/xoTw1n9hVka
Kb2fW/4reZ8zxfDUFMogv17dOgXbvPJou+XmiqdPlEO/9iOz8ipvmTycYxC/7nzW
qQDGMhJj2hR1+Z4Uw1oqKubybxOu6bSjLgWW5pLKfkxa+0kSV61S8L/9IsmkbBwa
9YKMl1usNol3oxGZ3ndUq+DlF+R+Xkqy3e9v2xbpbXaD2QtELQYKqDjCSokM31uu
itU3anX86RhHHdgqwNUb9uJYP1RA7UUfsYTMelEeplqo1dgOkpopF5CHLgKqsVWC
NkySEw3ctRDb6pvr8ABi3kkqBHmhJ9EEUKDBhBmYYj8l1de1F06KjOR9057mo4Cn
reGgxsX99fwP5odlBkPur3RVaVJeEBO2SCzJWjNVp7Sg8Tdl6QsfAd1QuE1bDLEb
UGiblCQNLdMeMyTZG6LVwU274jk/vbduFa96i82886KyvujxH5VcbhksyKufJetm
ymsQn2IubOcbzjC+8Jkt0ZPZv0L7zkAocVGB9dFk4DKPMzkmEF6GLpQ+CxLuan7d
WXGEAvCb7DKUR1N3imgVCf9u3x4LpCjeWWZbAxulgZwhnTcQLwCI0Fq2BTMg3ZYd
Ptxi0krna+1QbvNcvN07na7FImkleGbs7ltTJekO5GEYkEHAe5ke5fuZMMez5hlY
C6GCESBD8DSlQICFoQ9ajUslj01Vp0IwiHRER+olmPdBqGn+DdfAaMciLIbvErmg
Ry/FGRa11EbaFnqTIOm3ttbq1p3kd/JQDEzSZF7nP1DGF+VgnU8xuRuDffxzDegR
KJrk8Tmg9oZsHvi0R2NRxLSbRr8DgZtHP2L/aFe6tmsMv5wXmmM/bMpfmjZ0zLBi
yxV0Dvi3UY1ko5C/Oj4GPKmwJ2CCiavUmXI8uFY2UP9r8mREyLxy5SxCix3rU2Pl
ZbA+xcOPg0F9pRgYAAZ8QSMrOK15VSBm9CqmBolAMStXvQmmFv7UJe1cjFeotPDO
RdXBQdSiHNFTJL3JpAakLMiTc5AJfj4NDqoIUDI8EdKnbu99Wv0rnpw5+kF3wqlE
tWvgIub9zJYwlKlmqiA7msJvNOPSVpCSX90ZGGoo4GHYtRL1zlRa8wjqHBg2TiEE
WvMC6s1mflJKPYXUj86Cmr5OlHcBDfEjd7iTADln0KGSFX+UdmPjLpbBfB3B3jjl
piQ27WMRcqw1Q1KrLIsbsnEQpCUwE7mIeh9Fv86i7YH6MjJaUofjwMTfnWFiJUg1
NDYkj9CNpuuOwPSCtl/0kMnOqGsEYtbDw96RikSgD5W1raJgNz5+BHzOR8OrqC4A
RSSplukPZ+oNZ93Ge0rk0qTHd7djtg5BX4C4SSFUhOgS07FUqx5H1Feqc9jWSW0K
rfil2tCNlw2WuxXUxIJb3KOvDEQRdnXWcglNTUYVzzNE+wmKrkinkBAyobqv4eqF
PmN4BXCzBz+rpF6FuDnxLZZqZFvgopLAnNm4aKp+IQHtqx9nku7quboRKGF/2CR9
VWUVty5ESB94ultLS+n9UAH4FKakOH+erAJUFLWkfJxpa/eSyp6JNk2YHuLivRYB
L2wOIeD47n1SxlyU140X9MUlbfpMHFnMaIILEg3ATsJaWpe9VJr+aN0RGhcqdnY1
rBsdpL8RZJ0EGjDPdSSWJOJpYXzwX+si8bma2f5WBNMhb0hXc88DGRnYZK1Tl74E
hUZgiYLZtYEy2/qWQd2zKK/lCkdMvfbmdEb9vaGUnlZNVUIH872A9C0nfsd+Cfy6
HN9OBmIIYzUdxS1acee5mR02gYOHWxZjyUkD5FDRIk0v50UUVefWbyrXPXQnxNwW
dvvF+lBbwhG1KsBLoRVkfvEDkNXBETuTi3/2l/RCQ5doKeOB8T8lcD5i8sxy0eKr
WqXGCAvFgSmHoElmEfjldmdqhn+L33AyILJNNsj5HaBc6Du9JjH7C4+ElQSHsXnK
sTegr7P+7A6TZfz2hgPP4awo2JUELZQeXijHsdVN7WOD1Uyc70BVHU7PbFnqo3iM
YOTsKg1HHavW6hwTtbXK77QzeuEmfiLVukup/HGu8fqF8mWutL2gQgKP0VB+fkba
hYQ1m/qgkvdgpa2rj+0fGKn7oRFIXr9fUaUBvnlh9qDIlCCJOoQayL3MD13hx0Ux
QsWuUsIveOpPlOL9qOdegYBn3tBLKx53clXwYM47ylSt9ZutDSQE0ehPSrJdQq1m
aBXZVubPGVLfVtQ3w+wNky1AM6DC9ynvfZZzOjht9/avrnz4Rok0plnoI+z9ZKVA
xJMXi4Dxh48PVGjw2cuox9OR6dkfVyTIbQ1D1ak0YBaX+sJE4xLIIQDSGTRTN/OL
NUvCstOhLfiV4sY7vbf1wUNacEuQP/9TmSZ5DvEGVgimLXYfL44kMXm6+nIqYn6O
p0ug6OCE3Rdj2FXoujm+7AC/g1FT13LwiZQFojJ5DlYwRDQ1RqeNUr622Vm9pJQc
TGAJmQxR5GgvhLWqoZK66kkbcX1SknZtVzBLMlF+b2SFStoNz0bbMbx5UpxNdgjX
/m/6Ikz6NC9aK6qhS5NEm1cduEj+394rJi21COmN+5nyRfpSvLQ26eAo8zL79z0A
iWSzZCuPAFe7RTZy14KL6y3NIczgR8rexr6qvkBwOUtJZKbmX7ZESkl324SxLUII
XfljYNgbLOXuPeGeHy3XNySNEEt2LWGwBbP3OL9S7mmoyCT8LM76ZIEQHSgfCnLw
XojXHA1bdHlZHwCjXv6AgNw0aMqgD5nUhDJ+wyb4zQB2XpeSuh+rY2cDcFe1j2gs
HvkhK646oiXRMGkuWRhPNNiUj4T96beSLHamswmBxWwwKpgvEFeUqxfdB8nVlq8x
HCoLqs///ghAqmXFtP9ll2t1fOvngN1mnxX3XdneHjNCXxUIx8jimOFNaGD53yrQ
3jnIiPUCTPaijLhXcWncsw7/CD2BOKHyWMKZ5FUcvzDfPMJzWVfZ19Nl1RnX+Izi
oqO0jsQDrnPeIkQQy8N2sfIOiJdWxCXVoDnkW4kXMR2fRL+tWFGDoc0xEM9kd9E2
LpGsBCHnoNihy1xAmfzU+KBgrvvf7dXg+AwkS+JRv6U9FFn/Aihul9AzBbeQSw3d
kzZgAKZQ8K8vJnlm26Ma/HrGgSdYvb5gQNhmLzBYV0TbcInl9Dwu/QSlP6mnFLsE
2rPpuZw2atWTRxexJ4PvzVNVK6/l3ngQiDYdo+pR+5q+lAlZbDP87Gy5Ro6rYFLC
kL298TxA4hZxEr4FYymDOLifbYD9OXHO/wnKT0kr0jzhvQDwInhhwfPAJEl3unNG
A8Ho62E5ONtob76NOVDz3n9ZF8glwHdyyaG+iu/HHksaTzQ/y0oUXeogtyb3qcNI
+eEP+fqbOJtxNoo+0IULAeXvykh68ef27MmgmM0aiYgq8Oftf4p0e/f3Q/MqVRp0
tOCwHuKZMitans0MttPVZWJYQDQG6d3EFmG9HCCLGOnsJfG0FFj6+ptguTUUHgqe
SLMCj1tvf6OwU2BZGGFcEZr2Avt4lB5ndzV7H4qmYOGbdJgYNvSqwtyc06tZvR8Z
PuFV5bQrD1BgfhjRpJkbmi8nAOPOILfj1iRiw2jk+fnTGWiZznwUDNDIhQ7rS5YU
zcsj0fRjyHIkCaBcAASTh3kPnX/vZmoNLE/U/V/+ktHkFY8xQZXzdxEdp9U+FIjT
Z233YO/SuhLQpi7CazIjFIhrRUDvhnGb6INRg9o2miaH2QbvMA3G55wdR+r+6mdP
BCX1RJzOuxXdWIXKhORecgxuvJjFystQ9jkjIhfjzhuJt6o9KjYSn+ZCDK2eONqq
fDQrw1cHH8sm7jVpkx/+ffsrpYDCS2oe5hTL2j8vW+rmluMlgjlf568aq7U/ej5/
qSwMh/LL2eRmFuQoJ9gtZIj0PH1lEGfuwjCEIEfjDJ7M1n8v91bKc7BlOIMfJWLM
ufYyp2+ZPcvXgZAP9ql1pnwumUfRpwlY1KLfynbQQwD9LAUj6G+1HHbOVmhrcaAJ
+Zu1QWc5hpIlQviC+gUX/xxZWKegTeJrlyhIZQCe2os3NmoqOSWu0s4BZOjcVJUU
rU9PwXfJDErrYGkE6AV1qine3qkgFOEw+sTXSud4C1gfCVLnVVz9PnZ9q+NVmN7q
e4sDuLqpqSioWAGSRgnybZt4bft7trBBUD7BP/WBphPvFXSfa1gSv+ecG+Cvmeau
t7/JoL4M/uE4wakLThl28YH1tjV/Q6xljeN4psBvKKQY+ze3GVyPhtdzVuqtgNeb
VTrPeIEbwWevJ3A+QIzQBuet2yjz0G/aLmfcIXigYTUpGJsPoKi7x8GivxpnpWrq
0Rji2cowzp4lz86cehLzK+2Nvl0+NU5G+5J10Bit256NvfAtBf50OFjghcMa0eCv
4thS6CozXXmqZNPBbFCzkSuxMl0CaQk+162JY+oDncHqck2Xw45gUG3IXdhqZhPv
x3eY3g30dNePqVP16FcP4kQzgC5scpkcyp9xrSJHPUQstEPeVvcAY9aO1K2iNEI6
UHDmQd4xZxnr8jZFPjVlTv1I68dDiuYYwvVwRslDwbgpe//w1hmU8tsz3QbqPJ4M
ZkJk1GWY1txR2Q7TItx99h6BW80UJN9YShc6+butkYEP8lTPKva1Gq9m2R3Z3gqb
ddWsKwGIATz+0FRppZ0GIjKfzkUrh3WaQKFI3q+gHBxXTo3nRDHrF3I5n34xxG0L
LD08jdBoam8rav1WYtzBVjT0BZbaP+9mcINaTz2UUjxeWQAoCpnmX32eDhNnMuxy
ZOhYIidS2xGuKvG+09O0Ic2rezuIcTKNntwEKfnh1q2AwZYHRep/Uwr6hdUki7jo
E6de29vhe9ZEbI8jzpTh44ZuI61BBtB7NwDOQmSFyhXE/dP1KiduflEXhDY1qGVN
yKITx4wnYJa+3LNW5shjgpJ6fgwxsZZZvwG6iOZQksUAhhhXvNbMCdQ/IKSw8YUt
hy3AIq8v+g7o94u4I/F7rXaEZrWfudiEcOcSIpNB/wALL8oEojmTab3Np1utiIob
m+LInYjaU+itwiQR4vZgli33q5hDj/ZJ89oqvJ5P5tlxg2PD3EqMKxsSPX9eCJYt
CojI6JeBg/UQcZObbHNC4mp3FiJgvwR1FVSuIAGNcIY7LJg1nq8zdw6pqdokR5A0
LRnCS/rrPUR4YxSqsxvm/H/0h049kU3uVNCf6fawzoQBa6nH57CiaT5dOEzGn0bC
EzVJQ+SobCTwXPgrqrH9qsl19w7ehTgQbF6j2AXRzpLqaQF7dWM0PSzFfI/VWIrV
C2FKY1QqiE9XD1YkfTOsvnm/CauwauhZJCy9jj0RPXZKdnJD2iFsBODSmlXykj9J
Mo7YQIXltxK7DiH3FWUCNM2mxKGEPNMtlkisxtrsg1xbHCBGoGYOuHp9GVMCYZbp
aFM19Ikn5sKtcSLoorgnEU2qCJsf50H2KwUKaMTBNXfTz8ESeI1eeJz2jfux40jE
pO+/8aTx6VziWFiiJ26DwOtmeOGF1AeQthjPpDCsnSPGz7u6xehzsZz5a66REhCP
wlA8/4QuzYmxUa7A1E2NVbFr5M+Ye8P9QZ9Vx5r+SJTl1xQNAbbPx/HOT0BbqWGp
VYfY8u7wZ100cI/qRfw0xwSCVmaPKJWU4NzhIvfbLChYM6TNgAbgt4EiC4w2jZST
0ya6GgGswqv+5cS58kVMQAg+tzq+jj+oFm04+Ytdw/PqkM44ki5c6jc+rKVgZBpf
+B8wqjeWAWktEdrP2rqgwFniw5bK8KIaIb2k+3ot/BCzAKMfYYuqYWonWSyJrRga
L26RR9Jf3zCvAd+0VgyvjBmqkJCU/jy7GYxaB2FshTmXmmehH8w8bjdiP85ZuC6I
YNs+AeVumj299Ql7e1IACDJkP/rP5x2HesBe1/iBRSQ88Wz3mWgokWTH5eASXQU8
/Uc+20A32VVp7HIZuBvSDr/J8f3JBENERb1pk00q6Hoft6xsRKlJ4UGEnQr/1nKm
szF4o0a+ecxL0UfFXnz7IALTGFUyVSWx3bZNK3J0HD9EfoFcMJmJCN7mSe8/QdFQ
k6HAsOUmRay6I3un1rJMDtfBPOdvlJc8YsrQ9M6QD+wDu0Ggti4DXcKbgTogT7Gi
2XIEvZS+x424W9vmYFLcX5/b2JzVDdFoULPqgGe05bwH+5RXvYLcb7i5hPHNtpF3
vAq/UJ5BYt3QPe9pXHSCByEHXcPLHAiVPXn6NAWuuF2cd1UrdfnjT6EYBFYjRfFr
S+MeUjrZt4MY2JiJPEoLj62w7IHVR91ELR3pFnR/grcJ34sntzIBX+caMUtDe63C
8XTOTHtFnPUE2BHVE8M0JbW99zr5BFjwqNOJPWqcnZ/oE3u2a/yA07/hnSAaN2aj
4BDox8e/OJmqTR6D2GcQfCGdqJfhCn2TgxpHc7Yih/J98xcdtsfkWeXbn5ssByt4
lxpdpL6JgrXeARL8WfMII5TScP+wKwGqXjwRfdEjABHUdemlh1P4TzD+sQ3tjHgV
JV6E8qCvrNyojcNfnXbxqugmwKOUNiQCtNwGSV+pr6lCy5lKEXkEhkVxsIFIkEc3
/FqCsEdC8bOOXhCaC6QjZWkQrh89fOCTfJ0Bd6d/oEasJsV9uRMnGcFR8rCZ9o8r
RUs+Q1IX7dutkHcHv2olc46zanLbhFx4AzyriDtOWyteuwFHX+dFqWEpPFHSME/z
Dz9IFQfRtjQQdwM5S6/FCiViKcu/WRKmmDdwLmrcRoQMLTBmYhKmVKZRf8yK3+CQ
UXOCOoUvSFQNG8QJFZYbADQcQVfcCeECdMQ8CVHs8QFUhKVHDUjeZhS8T6E9DVjl
y3yfEnyFx4Q3CGSJK4j1Z9NVB7DTY2o3On4FPopHOb2kMTtwqawBIODEqJ3ctDWN
HQog+U7+BqaT1i5EO06AnSliv+bJIRfvio5B1eYiQteBj4tTzjloAqF83jxBDjQh
hnsWWd2I9bJPg8VP+P96BCbdzn87xklmiETra22Wr/aqzzZ+krqNeIrsfTO4fVx9
XVoex/ruBO+IN7DACUInOcbBoHkkjPXpiKLpm/h1mqSsSVzFq6XYOJHhZH4E2GKj
RyKvScZvs4P8uGSxjX1ooDkIqzbq2Nb9L/pzUF5vQQReTbcplpG7lbsi5pwp0+jY
Gvrd7RM/OCDRf64xaTa3zKSJFOWbiaexLrU7ejIae/Uhmaqz6SEpGFmpn6pO66tN
EkhwlZbFPOTQ6aSVMYKDae0g6z0pgXoMXdCEWNt0NFIIPs3gODjeLAA/wxyTX0Sx
qiQae2bhAjffdU6YLk0XYDBdyHKCsn/a/KYOyrgHFjyrTdG/TIt/Jt6ayQOnZVGA
02ekPL+f1w/8bBNY7Q/LCIX8Sb7PRHRSQfb/zqH1ccvkb/CU6viSIwe+Sj/ix2uG
rIz4P7uwa9n+f32C8K2Nkx+AYwMHulUl0W741mRz2L/K5LUUb3Ou/gi/e8MbEY8R
SIIRKDuhxl2yAWKlr+L7Te6Hpht6vs+5FetCTzIZh9+2EzjGDQvKTaDWCaOeRWPu
ywuWKUPszfcd7ahSpqgQ23XjQR9mBrUEdyAUj/fkLBNR3eu2VTYr2sHH/Ug8YZub
SnpK09+zcsraDFwN+07QfyEoJNYBNNGdRDZAeSSRkQxUJyN/lSC1ea3j+fIeNiin
UuwiZMN21dB1S3SOAHo3ww/tHfCiK1Z5ewiBTLNufgKCasWQOaIPbHiuC+xIcIMm
gnP9Q89BU5Mu9vSpQqSfSnhIwFsk6ppnZGT0zrICQqgkne2OiDCNRlfJ2tmo36nz
Zld3xu52rGY8ztvoxikNVObnSTwoJTvbLtkjDNFRw0meQxXO4Aeloo85m1sySU7i
pEe+qpUt0dsSFM6xq5daknhRcuZVpqhImx7jHTLU9jTzrWlUhNJfqjGFQF+gq3mR
ftq9lYdnl3QRemFHuajr/bACuLVzWCHsuBgZA44hCDrwaRbPYgYG8X9/H8M9ykHx
zmvJ0pCSme1nqjnxaAre7j8FrBDV8C08Ezshpzz60RtDg5HT+45oF3/I6yV2UOiu
lafM2Wd567MXsJxocir6UdMdeoprmmGVR3SYzs5CyyXJlLTWDC+fMSweSEPO5/tY
qqtnvH7f5IbQpGwxJQNXnfQ5q+O2YM8DfTOeRPM+5Mf7VzhHjcwjs/VmWucKjlAj
wwoXMYStiB7LyX7B25qKG6pOufuB5NswzDxPnvg3rGUbj6JxFcE7T/9nXF33MsJQ
nnkBxGtunj7+J+MIU9F2gMWc03yDTgZB7iEDp9QHX048Kxl1HAovw1R089X+5H9q
PfJlp+SZqZPmAjxZodjF9ZKBL0QafhluT9M4ZY3fBZeEO6b9fCCiYkAJTrmGtNQ0
Qy+C2/nfBdCSp5K4/7EbgfGnyTwL2gE/yOAdoqTSDesgrZ0SouA+CrbldqWEM5IG
Boi5buZjoLk9db7esxz1koN6v9tuqjsw0KURIVxhtJLT0nkqx4KORpZzeS2Vvzbb
zcU6mvqcEOC/6fPqjLfk8uN51u+rd6qlY4tJK1qdgJiZPde7dKaZL40S/sC6EMbQ
Ve3GxEo8K2myUwbpkMyvW26gKTCZq5QXVk1RfxIdZoXT9wceRqyS4olecSROiUZT
O441AmVNMNcX64S9gQGa3Qn7Jb8nCMQ67zV1m0dczzW0dG4LU8Id5TJt7isnJ0C4
6EFhpK2El6jUMC5/5kfLE4+AHJWsVGZezmioX6UgA55QDSiLGys0+dcVk0liYuvs
1LzM8tfStsQuDZb2kOW1qIrS0zo/sesXQrwfDuluBkCZmy8aPZlEbeufivRpig2S
5C5valU0aFDcXZskz/eYEUHf/l//LYezJk9fibAQviv3YAoS6jSW3UmweNZs2RqN
N4F2Sl6QcyT4Yrz7rya90rFjOVkdRBL5atQJUY3Ar0sQgMuS3mRcYUv8G/C3qCEC
iKUMhjepSTrOi0Ns+wZtB9zo96StnIkQ2UAKMjWAbwz4vEAx7oLU/2h1z946UB8L
UUUb2TF0TJ9xTsxn5am3ojr0JjrVH8Kr0O485PbxphWg7rIcxG5aTm5GiAyBaAGJ
a51y/6g5FxsHUI9Xxa6toxBiApB3G8pDz5LX54bwiaIlnc0uFSD7q0dKPRy49fJc
WwRfr6dd0UdZvhcZbgPOjMxoT1nsPucNum8Ucv1qxw9yI/OjjRKa9wNB83FYrJiz
ZCgi3xxNSWLhMcUVAP1KLdLM8rMUKgRk8XeFYovopcM8e/RskeCPCgNozJ2/Tytp
RJVoepZ08cmTQE7Ldg0y2S0n+TwJ86aNvk/RTZn4bBsnXYNKqF7Dhhs/3WChleXp
4YCMO/im7r8QyP96IKhIUjbriEEB7O/nuwTKiva9ySSGPFEksChbGTiHy2aGR37t
3yA4+c4FthiMaKYDyEVDN9uN4/a0x9/aRjq899YLgZfFaCqFadFkix8juEk0nUqJ
rsIDFmIVL9YmBqcsUQ6mSh9xjZvHt8DYqM2SMcAcipPxi1m/KkFJYRYyLa1I2zG0
/3LhtDiWYDux0rMxk/bh6OpVuMD5O0H7J9dmZ4VZUbgor60tRMxur2FJ8GrOXy7i
w9zICNHtKJ/Dnbc7/5LXOReQBqgYQpHYeUqag9Gxrk9uuPk6HIkMbICJ1GUm7h9a
RqlO+IxQ+rvIkEDQApYijC0p1ojQ6R4qHn6uN9ccifoxuIDmYUcR667iT3ePg0aO
MgwP7PwYNpYjmt+b7k0+bDWIHzwPbMoL8AAtG88Lh//SriMQl2v3JPN+52nNCAqU
wvz9boNH31c7uD2AGUh/cpqdRmTkhQ6/QWywkSKO6eE8SeKlQke4/5b1hCvnGPYe
/K3NBrPq7rW5LLMKclftTSlPlfyqsFxHV+Qd+VQ62WfvSHT8+iy7pxqiDqQItCkH
hAtSvbHOUBj1waRWVbBPmGExNDwv24vVb5iXt3VNfDqbJwBlC/y77mhXzTEcp2fw
4cxytUC7GlPwF0y1khRfIeK7CO0dVFbohB9BRxQOF2FwS1xghvyCePDsSrBW5kgk
1qXfBlcfn3Q/ezB9pwOnhmgp3fF+s0q7EFKfSg4WaG+gWhu0gmA4sqrzUawTCKXf
zbqD8vg5/neBiLKnJ7fZq597FzqLL2bLxOcCvttoxSRj8h+lBiCbl+t/3Kw3z6iT
S29qhy858OTSoO7k18sQ4kvfdQMkIm/MrLh7K/9apySDBkRxssRUcRimQrOgjS8x
8LB/xT/3f6zG7Eglkw9wTmfN6dTCXDhwxUerNlkiPbk9TS9RItCzDW6TPjbCyyjS
SD53CP+wQ+hWOonxGgc9MnO158WP+83OY5lhgu75bEkM0tSE8BpOC4tb2/ZccNt8
w9QesBkKkRgGyZI20UOh7EyBofJyWgWHY7uXY3JGf5w9JP+2xEvQTurc046qJdcK
z9cia6gF0S3r32kEtfFSRc9iTSUk/quWjMISLB6gtQFiJZHICdCZ+7MlG2GeZtLO
Uykf3me0D5UVAxNNYZzR94RZcXjwG/IG8xQ8UGUvWclyjTflUGel2YEAiDaV0jg1
5U6LpO8toCmeXevuWhBZd58/AbGlNTGv7iVHQ3mni047Bf6sN8Mfa+TsOKA5jgxX
DkHsUHxlDlYQlLYzKGqarqriaBincZb1HHvX59Dv11i1dUrv4eKU+EPFTVrXrfPf
GO+o60cPp4n+2GQ1aYMqI3/NJXYNjFdF4D/u8JTUUf4dmUrQoPFT+7E42k+gveP1
gR5/xCQy0tuilCW6WrpZFclcdOzDiL79v0DQWuZpr+R8+AuA9NH6MV7MxEZURyEA
NAVarn7wMqq6Mjzk/ecwGa7YHwULEposGN/TMx2M5+yzwku/JAOY1roAe82QxRZW
SX4w1p9rMSz4xSQY668khQJYiEkf8pFlWj6/wil5lFIQLnGYzvPspMkgbYZzXr3f
2IeVK5olVIK68Pp1/PQNgunMVzMVMm1Nj0/+XTOaiuTCQ4MkUTaeESso1Hf83+zG
cCg0+at1nqg5WtGx7M8/DTlFYUx6TENc5hiMn3uum7QRg+Fen4ofxfW8oAgzi19h
8kLI87WTGxy4TAT1Eb+BWCW4UV9lkf+Uw15wtzK+WkCx3B2MsvWNtduVQItlAZ9S
XueCi/SeBmfkcyQOs+TyY7WjschC43qle4XNUuXc/hyEaGgjEeCVSFqN05VzCnHh
NDR3H0d0ZlQQJ9V9wGppKHmBIuRm0FCdXek6UBaolnGk8ce3C44KGFT9GMUS6PSM
jv7bBHLDoPDjOUqy0oBT6Wxv/jtboKzRK/slFn/6whZbN4bRy4zUAqjLoP6aS7Kt
y97ura4ndBIbXtL/XJ4Y2aWlJ0kVXK7Lvdg3Z+XeRGfjCRm9eVyQhgCbIwSEx1Cu
CmfNGXgw5CfBR4Hf3fIj92LceCa/7emjcVsEIaM059UOCnMgn/BlUN//DHBQS+5F
mT4ABB7L9KJE37WaJdMN4jgz67dI23zIF+7OGA8W2VZMi5xr31d8MzXheLdtX3aL
5wc14MQqZMJptsadBvMk4LVEIOAkjuaTztabllzQnTr1tHDARLiM6xL9p8fqQuI1
qw0mn01V6OXUW2rqyci1n7My7aG4fnkFrdeZI8cKa7iYvZuofN9He8HjEqMtPXP/
2WLASf0ftEIgXrWr3G1xOAYLMGVZkBEcPJv3REnjKfoZrJPvdd2c+0rbjHubMSus
mR2OKYuCCnKCepHNcO3aR+MOx7myvQbuK9jGDMf8+7v8rVpcGFP9X002fBK6gYQ/
nYsFedG0E9F2i+1rx8sGA2/UntWbtoJ89hAZzhokhlqHqv/wFI5akmsgCmzof4k9
b/nc7Gmo1PojL/nqYUf+xC2TLa4HoHr08e9ZiWuhVA3ur5Fngpsd8MwkzB08bQXO
ofeHE5vIMd0pQZzp4MGu7szK4qpzSbXB0BcG3o/ZHQeOGGbowUphqKED7Y8F8MTr
wmW8TEz/A2H2b55S3XI0s8XukPpplG0ijBThTk/qPwvab5qpQR7ZFZyZ/zg/5tei
KmTjY+WJzF2tIVfBg6Ku+J48heeT2i8cqKFM3+AhCLCzEsOLKkwda/K6vrX60Rco
f59t4VUaTYJv8vuW7/qca1LPhDvVO1dReSza9G1KqYnDncvlvkPY87PCzKHKGEW8
YSDmWUyELOBo+xU1tpq4z7xuNThZS2D+igk7uELezoDbgUHP2iVu4rxKq8ChhI5A
wJtLAg52XqW7DWA1r+B2deaZ4VoqUSFuMU+njizcmEfdaPMh0ddvf++v+DRGzO1a
6DgSWXxNO0EdgxA1XDqFGfWtmw51bWPuVqn9MUgg4iefIWUx7aiI7KnraYs/esCD
wYAdHsXm0MJGn8i+jPlCHkalXaUGCOCyDcTjzdzNE7dnlXee8+/zc5RDIj55LR1z
u5AIBPNbMSNPXSU6+feH8JCF63Lqrd+djknq4qAfpZV0BzAWQZUYfamdNLixUN6i
K161joTlymFiYMfFSkXWIvLx90Vs6s4y8nWI0QDcbSrVlyNQJQVyOk6kXnQpur8G
UWDcBrlngm5n1zEOSYV8dJQouDQXvRcR38XE951dIuKQx9J4FFBRBKEOkhesOKli
Yr10ZbtTIMxM7+RUesJNYmEjnIY0d2tyoeaGABl8otk/jxHq+9SpAarDmKGdRrt+
UKZaWmn3q2MsfTk51vCB4VSt5mFuPr48+0OidRMhB5GD2Bu164Xc90pfFgmQYIEr
6nNtw5qoJWIk/xxlDxYJHG5nzrrM4c/AmyOWSajmlcaY1pkM7UFxy556eSfWBrTQ
BC1kz1/2aYJxIi/VsEsLqnBriUv+jnU3enlQBgdjardMqIzLtk1H+xIGT7q4dnvB
vVKB6GnF8mWMQru90o/LadClvQE8H3KrpS1t9ORJjLjWm3vwZ+yUx71ddtnQVZCS
k9r/Gt4IcE/Mp7H6K82TltNFDvyZI2oEBQq92shTR/uBRYObxeD2cUw6196jHBa9
rhvBroFGRKwjVR1kX2tIKBryKdFj6lC55f3BSnU5acBPJ44I8HpYg5+w/OqFWHMv
0i5mNKFSZz/W/RV4cv7HXQkOhv2TzYiVDsySHgiCtRInK2K3tKUIFDmFGg9FIkE3
tpZ6GueJ5kkMSZDTZTDmHDhs6Yg71TIu4u/JwI2CvW4jKH8kI+K8HayVmXMM1D8r
QX14X8spYhphZeFMGgPnn2Pnrs6uHQgviIGIgWoiFkqcTS0Apv4WhX7LzQIqI+9a
HMM1LAjZT6yJy2pmOhDz/skgQp+kFnkYQf7cM2v1uyFcOuARB3d4GbAKzblGS8pu
LR7Gpy/F+ksf7mTomuUzFkidZOtVbnoVHylKRhahMpS/F/RHejnJLsRd1VK+36iq
VaGfDvLdMX1CXA8WgPp1Bub3drbkwJ2E8yiaREwLwNKYAaB7fFoN7mXoKn5Oqxaj
t6bdAjRVChDL3SqnScTx9sdlqd6+3lRdanXhEe7gb9uqZ8g8Dy/SA58pXa2YMMaM
BSjinQU7ygwPcEPQYYlGr7KcW2nholB+Onv/WDw+2cHt5NF918IUuzWJquKlMSi5
qd+EL1GB7i5UZurRgJDFeFS1kr5IpTKJDq4yt/I3bMvTRzYfBMGsJNRSvxp9uJx4
8WwW+tccSsCqeAdvFCXzjoFeeTJuRe1vgiMnWT4kkZUOBq6Iv/PA0IbQp5srhvG9
0Gb8z+CqYWYkUEd3EIcIrjcwqnjmCTS7Sv/7c8vyyRqZyUxenF6XxiUoEILVjR6h
efM32ZTcSFY1a39ydLKnBX86Y5i2L0EazsZZf/7aLf7iVUkILhMVRhDD59c2KIIU
kadKp6C1DY41Y/pkwmYNIexhY4T/Ljl7Z7D3ld2CVF8VhL4Id0RUZLC7KFNcnaHY
HD66qoYUVN19bhaDRUYo4L4lKKC5KgzWvpMED6t+9t3aUT2SMfEbQ1ql8S7ZEohA
OaI8uqX1MaQdWhP9vTHOOoNIjL5tPjXEe6Q3pkhoG50S6uq1UXfyr+LlrUt1K3ul
Aq3T8joQyw6PzhAB4jdPli/xQyetO+7pPKSA/1Sj5ePU+nYKNJG0dw6OSTsId7Dw
rvg3dIa0xHjouMwseAMIBqePMLVhjupDWMQSxfbjhsxQ6Hsn5eJozAtCS7R+lePB
k2xfpF8YJSqrcXda+UYUsJdjTAjbY0DabdxWX3CFv16rvQrtkoWKrBCDG9GBuLk2
S77elDuhgkbyFEbBtJA7gaUikLXOgVP23qsnQdgsr1eBXj3nulRnZLzgLnilVO8d
89StnyuyeeueeHYSCiX0dJoV8y+3rO2v7uh6PiuG1lsGtAAGCrwxu7Sc4wNtX4hx
n9obDCO7wY0xOEq5pPUlp5RSu3EnDrk/QwenNpJdYj2BKtOuTOZyiJA25oJ0AG4x
i1J50VXcaHYPAggkzA7Jpn2Ihxaqk0GN8AfAXav1TckLD3f/Uk9app1F7FhKXGU2
fY5IQWURZ5JhzRwI+m5vjbFARK5dGCHuf1M3LhlwoB7CkKnCdXvdsy1+1WrzaG3k
394XUVcAz3fCTH9WFEjHPkaH07JsFsHHQ0LqQJS0u1DnXXIq3d/AaxytkbatX47i
EmKO3cnJ7z1hWUa8BrSCBsuP1SKmY/TIkLGsg3+btpj7b6FygCBRLhTeUxlg95Ix
amhNanAps4m8nXqIAwNP+jE7NqaS5Wg6wiyd7N51ygSEVcg5pbCbhece6ktsnJnl
cSIVbRY0Li8gLnVR+EAUrHtrrbqEqHJj8u3XR8asc4ConRf6+7e3AUHMRbuSWDPw
acjFxg6UqVCT5lHineyW57mNHDa7wG1fWGglX1JPuhhqCkkgPvWbu62tQfAFphjm
x88IZp2b56UfT2nhQjFS1uaZ/1Oy+h+LjHBwNWNSu0Ki6jNLnB9HCZ0Yd/ak7sa3
noyOJMW/N3MPU1rMis7JgK9m5DvSwl9rAxpDXzSCg7TiOkl7axu64eUFgybXAHr6
UA+HZz8qarj8Wvs6fqFa7Gscur9LlKDcu71xCVDI5ZgPHYtgmHHlxZY/5+PnhdL6
hBhyKDtU/Ug6qLdpsWb2gmdej4fPuwAjMI4UhqVueJFDRttsa69lnI3huhWhMX68
iq8yOLXvUTKpUXtpsoKJ0PIDCS3I/37hSeRA1PrIGuggRgB//alxmv6WROkxoWsx
1gOfBe5KzlX16ExuKdJN6RjcYOqnvnACPitIijwFUMGnIEWaHmLloZS9TbG97rCj
IXEYBtWJbRN3b4G7vigzAqeXj2bp+dilumstPC6IQmsi5FR1VLhkevJdDC2oeN38
kxCXPwIToYDi6fV1oxfGq/cPbUJYPNI7M/oosBh8m6dNz+ZYD0lyfy3TFqv5oQGv
wuziT2qc0Gapl3aIGptkEPwPxGffqtJR5XgBlvO8krbLW7fkcHkmHCEPPnmtRlbs
CH9F0GQwaHGRWvRtBLgH+T4qmQ4G4UWzE7vsr5JHCBfKPb/6fH8+XzDScxFvBIIw
8/DBJUzoX/wuLhxQCu/dnF0NHpE5KLpVxoewAoJFNCz4XqRQb327n2z+5dHV7MG7
eLy+XkwTbtUfgiYDJiS/UW3rVIjSsDyEg0794SZ93m80Hje2mE06WiIKVZO9uLIu
2ZqTfQsjr4CbnE8PeC2SiCxtGhB6zNaAV3332BL2coAs0TDxHo40My9prnnHT9jz
zfFvP3RFeH/oc8grZxGxDrA0Bng5VjKX0H5KZjuSHUCWHcu0f0KsMMpDVx/Qn33P
vCGx6kUUe3DK6lUOz1Qdik2gb2YM4HE5GwqNmukAvGJ38vzGNJBR9uY0KJYgq0eh
qDCBE4hm6Qy53yrjkY9JKyaxrNreB+vh3DNWsCr+Wq6B57nJIQqcMsTPyoaLCIYS
pd/HuEAX984ZIsfkbTLgCrbvtZUN/y3bbS6naDmNi8fzbFn81S5vM8oCde5yBxOP
chzLSjRNg6FYKkHB/77w9/Hll4sTZp0DLs7CU6l7Ki3S22gNasQgo4NunKEeMYAH
CC1SCT9qvJi8YS8awvDXrgKblBoEOcmxPq6U5wFjKiAfAOIT2QcxaNSAAzXD1FzM
fCy4+3a5srRtdffAc9LzMz4XHLZvrgt0AntAfn7sorWdtAc1iK9qTNxZNEGnFLB7
U5ty3LgcM0Gky6GRb39LiZ1xhlCdX8C5JnMmELiLV8b9NJHc9xWWtnhE9y6gmnst
RZPAVS/iWWyWa3lY9+Ile52Xib2R7uhzRrMY8FatbQohXsgoIZrwLikMHBZbzdxD
dU6LcO9lhYeCr1dX9JGWreiFfMUQW7PDsLf8reFE6ttaPcqMxGZgaM5ebKQPqxp6
eKcfE8WuUQT7Yp5iSn1MWJQNL9KMk/cMt5pblJ7Ss7bFjDEgg/h7pj0NEhabSoEx
RQlw9IiioeZ9wU6VwaecKUcQdxTYk2uqSjKUCTfL/4TtK3UuTbyMdk4Mor2Uf0LL
YoIEhCW3Inbn8UEa2lHISdCATQnHVPs+D/zhvuOnwwNzwffpUvKLFCX7+RvB4nvE
tfa8rLTt7v+0+2/V8mVxN10IdITi9ejRnvGH6JP07EfHYN8oGlY2riDxtGbH9mAw
jEBo0//a/VwNG2rnq5HdtTx/OcFSDpIIaToUPNW/QSJOHJRP9ntljcjA/WvigaKC
Qpzm854FwjD0urNR7aOhSwnX4nN/JFKL620YTlSMDa4ZFdJYVMonOU5Lel+MQh0P
/OxK3d6rLzFeOh2yamYlDQDR/QtB8u4peah3cgcEO2OnNkrPzb087sNCDMkbF5FR
R6shJZIsAR6KnZP2DLs4Y8cOpc0JMa+amPJLA+FsP/SuAQbhqpR//FZ3dz1NP6B9
SwrdnkRLfant/YiL+ILZLDi2re3pN+W+ZVwCQjHXarbeWcOwU7EKXjBfDaRYhZ2h
OUEgfEi4rO79cuD7dM5rVMZvA14TIqmcpqE8oKE6I7aIeP96xqPTWGF4aHwhzRmJ
r3xSPeiLjDkTd7Fqci/AM9wWKFAvXhYfr8ejot4SaeOVuF0mOu0xqkBif1+mulYl
3iz03MzooBGsd3CRwx5y0079PdowdMXCYkXDqjQqDlrKFLNoU4Sz51G0kCdcpFfo
bcz0hDe2OOm38BamdjsRm9KrNx+Zdq04jCwUDXUpGK860GvPGDaJ2evD69IDX+Nd
Rt1Fzk+TS0OLWxThjcA9k3QkfA68H9vPMdTpSrRz4HFYnnJI1hSvNmhiAvFtVSL7
shJKesQ/z5CG1MpPNNFhSFByELsQvSK+cNyIPQVgDgK9dZiZ1r4KNCcNAFj5gr6Z
CF3ls+N1LZso4I5sAXs4UCqA+xivHHa7reheov9BQo84gFsMf2XQzxOaYeK9qF9x
tiINhQelvnlJIhlLa+WFfHu6EQBPc7T49CTKeEDVnLkWG2AN2HsJfsbh5/EMu4qL
9OV/QE6Yn1mdWIUhaB3i8433Hpv8PrL40Pv0b3vsy2IDolpLgVNhgVroYapovBNV
dxul7zxWaSI3gYgURdXbafhQe9vG1mH/zFgG52yLXqaeQin7JHt8c8ePZNnWs2Qr
wQ7sDgK5YMvk9DQZOZGD9SrNBAT2cIlcG0qGssvxhkmuNzBmfvjyf3+haI/FzzmT
Ftc2XbidMh9u45OwY99IE0yRBSzhZ3wZORhqF4zRAlirCwIMwdAbXyInFf3ibahJ
+u536Col82F9CPrOwJIE7kS9Fc/blsTjxoeAEts9As8EUEtUisownwD72BxK5JtS
Ad9gscm36L/zm2GHiJ0sLxhBPtuePqlVjmKANdySQoOPfnGbgCVU28Q2TNnGwFlV
WM+gmpDz333bhVYTXZzD3aYrMER1OmMYwiuQYMAs9ul4CkIwgB/j/Jx9KoEfoqG4
1H6vO8aNW6PlvexYzdGx6DSJXvRDBZnXsPRd+G2oycY+lOAdrWRuuuojDpBa/Ur5
HMzs7CRG+f0oUudeyN9lAYteRdBRkBAYAIJMkEuzNEirb50HEP6eCfhaUiEkKOfo
AEeRZ8bWijPUiNxZFj9aIauWID18+2guTO6Rz9EwZkf2rCccOCRTe+8EeRj2ySIW
ZmLJ40Jo2NVzGcibtrUm9v003zbtZ2LKpygPoIS7pnnMRkGDuOcQfxmROB/Hb+y6
EhlUPc5EhRzmq37dJ5St91UrvxWk7SyjAZyaTOzATW88l1R+m6OqAbKn420Zd0gi
shvGkrMeXv8t04YI+viaojyKDt5aHMkfTNAwAszgn4nvhF7qwrkfGoZEZ59mh3iA
ApkbmRmdfYk98X3em/MmPirL7SXtW39pq4xfuxfNzXkIrGdEWGk+8uibxRnGdsYM
Mp828fLX4xux+Idz9pdfUVXH4Wv2eo4ifhdw4fUmHGRzKHor6ofM7IsTW+oHa2qu
M0bjbOpyhWtjBctcEqrBmJihLD3fVwCka2HN1VZv2EobV4NpCsqdQd3UbhCFB7KK
pYE96jLJp8PWNPUdIy4I2PI0BDx2vkl079b31Lj2jAdKcP7gi6hUTYNH00CFXWGW
7WIXa38hwAK7PUOzmQxeyJP8UWJwI3AW1P/vE9sVcgaUyfUz4u3LXenmj34+kRla
o0UC7SL1MhGCgeT409oC7eMbKarwma6mteoTGAccMg2Gf+P3R3U4FuIRBcEFx7mT
Dm8yOOSrEvAJbmHo+UoUu4L0k62mhxyW8bx5ZPdN+2fh+ZhaAPsmEAjEj2Pl5aiw
8yx+tZLz7m2AKikh62Qy/XfQdiAdrbJOIvnSyTSoUQtygJgiJKCIhJvS4rP6xwct
kp+g2h5Cy1PsTBQCzwtlYiVo2dbTwG5mcDbg7MC1ktBNg0cslFQBpOIbgXcpnGdS
EjQaHnruJd1pWIiC+QsA12z866sUJyBnEygSZwOvUhUqCRBaNWTzmZNgjcgAJiB6
XpW4P6FGfw2wfpQBUBWony4+1iWN9DfYwKXXsI+h9J52LFWpKSmvz5BcXGlBvPQD
a5gfOfWVD2eW1jXfOmNYCdeWyuivXKGa6Dj1BPG2EWt+D2XvdyQ+NbnKHsM0GYNF
2unXIrS8uCE4H/6aE1znFl8mzjXEPCfzatWKxkt4F/r35FCD8QiNPsjWmpIzFbK3
t6eM7HQAd/1Uv8jm7/l5oez5U91brAr62C8QLjNSylfKWTGcdxdy2NrO7ldNl//2
V+laIZuFgpMEn2WBVzqnlvXteFqrLWFw7sZgwV0cR6ybWgXGTDISX1WqZvYyCjnh
LQQdk0euD88AUh/ZJgY0kajiKzTDibuRufdoPqabZdCjCy5N+Zc13oqrxE+nT3qI
p0WnALc+QZJLrVz5wZP5ZvlsUK5TPkz3XYd2YrwVA4P+mI0D6/oI4WvuwSZRuu8B
V0IDILt87YJfUEcJ4IlTzvmefA8+zCoRUeVmnLbDASltXQ6mMHGdQfSPTfRBunaA
i1uBWoUM4s2pA/M6BeS1l+5mG/lYwiSPAq4ogxnvDgnruKXFFZuk3c/smgL/Ew3d
RHQwOYNfFayXaJo1cfgqR/jDIlgDrAHJ7Fi2AQNq4Lna9cWi7EQ92PyiNsAJY4+2
iszQ/R6KKTxiYMMiXZ5h1dZaUXt6dNysnQcLO0NnYptnJfUFdT4Tv8qZRnJguXD7
vy6cMok1Z19rkXptxVVpE+fKB/trSiU7MpfMvzDk/FmLjq38ez8Xe38RJMeXEDvu
6Gazfh4MrdNqCtY4TBXe8ODucGOuHtoE67o75SZ1U+moMlrMSSb8FejUbpJbr4m7
9VvefdKQPsBmaZqncG1Nn9c+GC8oXUPelxa3JzqMwZWNorOZOl3rHVVaKIG4hJVH
ENbA8uKDUEwceF7FMilCMcWIxPUeJUTEpBBXwIi9Ik68FGb2hzQ7ZAoIa+n01sR5
qZoiGlM5nApKi+3FyQS1AzXn5DPL+xF2FyCc3ydIsCzOdW81gTSpFvh6YI99iq7X
8Qw4Y+sZo+dzVp5iHOSGHndPaoYslc1PnQuVEX6sThvKTN5ZYvh0Rzby3vP+Kwji
K6qPIbnVlbYuMpX/JRiaNLIgASczgQvztfmfrstBhn/FtTyYpKRNrw4FAWS1IRBK
7jWN99B+vDc3wZeyahAZWRtWf5GBCsT+1wKNhjyeFwt4WRAUZaiQQ2rOlI/9TpAX
4BljIF3Xv51x9ixQAJ1PFGy82wK/ZkybitBMstJhjyF4P2k9z7yYfKYGufwiCuoO
wu7teXP7BmQ8IlmfTUF7IfpHkzxgbRtpC3pWYAjS6nIdhpI21LemupeWx0OpPYCx
c5FzybZEHJLn8+W5y4cxeQURmr2lo1ZU2uYJc+M226+UpOmQgK0K6zp/5PnJqeHr
CvrKya/SFKP3S2QcN2Pf4lbgJx0Kp8qKZ++2Yp6CmYDVEMSrY/5TV6UZ9RjCOJ4q
tIQmmXRoe0WCKL2xiFp7EfeI7JKchfVj01kWN1APV2wCn//6NA3WyU6dFWj6Ey1v
ABKL13zTjAhixaO9EKvzNx5Sb7+AG2QbWumYFcCZVqyeLth2n5oyAlhooqeoUJp5
3nYF4zC18ZFAZQ5abM7+3bzMJGGPtkI7cpywqsAcqgebJcoyAfNuGO5/aCZrNyUu
N9buDARPj8fM7PZqB1cPKACffcH1JkNFwjOh/4qfulalTNQsctPu/6Yk6s3u29cs
8YevOZzLEZGPSVtI8WTcflf4bNamiZipuqsSQop836anfikUTD20oXmIBCTW7wKC
NOk5iaOw0XcB95M3v8yvx9usv/ySMF46SzkxYB2CTtwM8b5QyoWCaGld9R9Gcayg
qyna4fq7FaHaQ1imMOrSIRA1vPELDWlIT7/OKubwtNyL6IfB3teU+acD7AhcJbrj
Pq9JDDAZEKZz3Pxb9ZJuVOLPiAGMucmcEyu9cBQWOcKf9TO3Qu1Tbf8oY3FtaZr8
kycOVu/J+oIcZVWamcRynhSwuqyTDlMNQG2rxmaI90MrsSBhuYt42emFMrvJKE2H
yWH5/t3n4/1jrJiOrSU45G28m6IK3VjoNMC4u51L9jot5cd9zw7vLM2NGNKSTijI
sivGHinLIV4mTc3dFauIpQqsGo9LHiN2Ow4Ad+YUgn+uwPbbvQfdRGnh4ve9Il1S
NjBulyIXhUbmtCjSHKvh759B5xgPzc0ye6mJy609Un2ZuBnMA7xKTSppnx41PiaB
Me+Kq17JhSWjEoagkQC0ws8zX0tghtHluUWCsJHHYZnPdj7Npbw3IpLyoXeWtUPQ
wSE71lHObkgjvhpBciK+O0OXWNRgjD+4tgpNcX1M601OoC9mlkYwzid2Wr2X0aK5
AUA4jT9YAkorDDN2YovDqqklFsThPpZ5uLbVVFZcvFMrNOvRIvYuL2Gf4cJN40zy
plVBmUNB+/zP+Q+fA0ahfwcOKFNNfTWnY9gurUwb7Gfzmp4DKhd0oeqOZr/Lrz0z
Sj2c0YXwmhUitjJAl0cigzpyQHDGXtQx9v6KwjnKRpen+aF9Ja7D4cpJZln995B2
5Mh0Vf3bvJwTcxhd8T/udao8B+qE07oIBX2DFGxIQRDUbfZbS45359cjKcfULKlF
vtJz7PHX4LYJMchdrekKTUEon49y0Wquli/m8p2yiafWcOUbRIfNddfWEqLRXfRr
MmFV/0S6Q6tajugei5exskR+WjAeSkAM73L6iliUrP6Y2YAxlfF/wxraGN5TmDr/
QdeA9gnHpOWlRbf5el/6LWK2HVlyy4kyIPzzLd/yMWuPGibY7D3niWKruFK637Na
Jx2Utk1a278uADIw6GTr6c5jFbug5uBybmbmhwPKYdFi3mZTc3jr2kzcwta3Ig+Z
NHI/C++yCYZU8Nacsf3iSpvYvePzKRCJfgWrPZ/0YJdTyxgw8jHCjvL75A0P8EKU
DkuvPT2wHAXFC1UKHfWCzjEX5K3uQvqxDgtCJzyUnwerK+dAe6jwsZq8DzM+4klJ
XNwwyAVY/S/ngvtWOsNp52C9B/McQOPKyhduMrC19GhifxEkeacbuInW6LHXfsAA
en2sRPwDNuBfv4eOssTv21gk4nD1/sF7eGBr+kgFEgzqZgkfJSvvGS1Rr5tIZb8b
g7dNPARKVMOeFoP/rTczORq6syfQSmbqfVZOyNCharjysh3qjbnrRIvavWQB32Kn
mEJP+BzVpfmbehdRoy1nb6TCK0tgAO0GihxaMLRIpQ10qHjODT0wNZYseQ21g9mn
skOTnbW7FhoGtCumvh8xLTHJ9XKKw8jQ+jzEqcp0VLJ2vhegi3p9/9Wj/d9LWnwk
JsJ2TUDefIMf3U0HHMhCgxnX5loJyZbKaaASVqqDZHsKEdByrLXcctAxuzPOBEQD
+hsCNOJnVzf09ZUhFHr3IlfgG5wFm5tN1hFPpkKicNvDZhqM0GntzZ1AGxSGcUPX
nNSu97vLaFvZEJvmCiBPxOGucb8vfxJK+tBA/CaqBbtH8iuh8dqG+j6Y3F+i/ClN
clP92hXgZ4wVWv88cH9/xpXhQCH4P/wvlcqblXaYy2+uyjYfCUokHGAjbIAh8Qx7
TQv1FdUrhwwdZNriSFMG+aMBJ0PCTiXTqhzCKvInwenGZe7JkIRkyUTKm3M6fpSA
VVc0RgHTzmL58WviQK9QWHm8qgr1+yLNMbfYJSZcu4D7VD2h3WQ1YfpQn6xwpnUW
52awKnYmws89jXazooiRSGg18T6Ny6S3N2E8lYuCHTOP6wkzaxs08C1W4s1rEIpP
0aGBrJ3AbQfelrY44ucG62pNT+aWcvSIVXLS0IHIB7wOFt1wRl0exFf1UuKazq3K
5L7hOS7UHi47cW5zH8EIah+1WtzDUGm/ZphheBgZZZJjLygsWwtMVYBP70Ng4QqB
oiox159x7E4hPW5Jfn8cXZl+sRI/JKtDe9rDR59acrwaVLdlKM1uxLHV6UrnSNfF
a94CpjDHz+mRo5w5M9n70vhC3yE6s/0PJjkSEkjEFLTGQ7/VlrqFYuz2f7ctmvrO
M75CFMSmfWt3CJeBehnbhs7FuZHIn9eiIOHYFE63OCthZXBU9w0DpSWIcRxzcRdR
mO6hshSksqkobvyvx5H/cfd7CRriuQXgFnj3cq3g9KNKIphxK4sskejnIYPLvq57
o9PowipsvpgSAdwwrJ0fOJPmnhvMMAIP0ys/OAKWmQ6e4YtN66fHA3jWkIvI+gB6
kgty3oE4DaS6Z7L/S/p+vCmgwr3Y651txvFkf5eTarjRVdzPsPDY1q+ufLQ49y/i
pzJ0w0S6ot3FtIJMkVSf7piCUYps0WNX6qrXYAbhiEhnYXI+ogyFP2+ExwnYZinv
DBXkMFnxUuBIVaO7J5Y3DFEa0VKmyDYt/27H89iQYF7cJbQJXrxCTaN7K9OS6nGO
+ya/OmYxSPVTKD/uVp3DCNzmfzFyA4KTX3pji/Fvq1zl03se3EnbBie6nEGZER/a
680CnamMB+P17gdX6UMcOVC9Pg/NrBI52P2bncQPvyJkyQi3EiTk9+qxxAr6QclM
w16AnpNZ6kRtUauL1HlXAeifPnxAnD23Yv3d3VYhatvs6hxv4zUoM11HwL652Qg+
6XQ0N2KygI4R9A89Ke2MfvhdutPBuhHCFVNgw8iy2cVq+tDSU2E8G/3HKV2vSYTl
PYjSSq4i/9z5O0pZ2nVN0Qm/3EZ+BNkb/ftAOFbVZFsJJYH1D4D2/BjoNFW5y+rf
p5C1nsHe4lizKPZchwv+G5MC7PDabVxeC+fAGE/ZkjuRsLXJjctXjxKdDBeOHbW1
SWMCPPVkbj6RPLYp0wLCHe+NGDDHG5NKlkiLdm3f1Rp3zFpkgJmpKz/5N0Iwxj9I
oW1k/w7Zo6yGfIC5QIHM/Zhxv2htP+P9iS5pN+LyhDQH8JqBwp1x+pSO44JysiE9
HC516VBpB57Mn7OjaGFpYe3OVC3XtTShoY+DWuOloFGCMCIzlM/5ZydMU38k+4D+
0uSS67J1LDzkRorgEQYmHfUHNycfVsTUVymmYUbUeg+mGEfuRDNUdiY/5fFt1EMy
2xeSc+lSxuU0/vWnlUwDfCvVxFefduKP64F1+gaiNQn3k5WeegUOMx+/rWthpz5K
T7U37mxPzTF0TvxYisr6aodZKgCGzHaKKfj04RI0WbyBJKhAYaGXwC3Cjxt3SLje
+ZYDGold3c54Abwz9QuE1HiIWEk8fneQjF4b4Tpdcyeo97PzfUEfcERxn6Hiv2JS
QAraKhLAwQEGIFhggA/EDvdo0WT4cqDQik3UgVmVYHnXlncn1UmVTOfrTVvVAQ8X
adngblIjiA9bkOLZzN7Fpx2wUI4wosb6kwhJ9EtVAKCLPjjy960XkGG9zB+mX1/S
zcpdZs3iJAsF5lNpivY33qnda7ZjKqUJ3EfJvFW/j1n1vy5Yv2yBSn/agfNcIYu9
loItfJqDUduWVEXTH2JzNqz1GNvWhA7ZkfOhxcW9/op4nieMPpVH1IJP+2QvmJal
NAMht5M2ykdk6MzMSUmc2X8dmNTut6aoo6m8GddddQyHZXxLtA1MIftA3DYZoMha
mPPIzphnm5xxGkydRgUPiKPdPBYj+3vZVbSvzuqv4faQZ9wvDBrG4BF+ZQJD5G3P
AOvtPwjQRQ1XmytNu1FK7Xp/tarvZYCrAH1gyrOeNZaMISVcpzHfUQCh4EQlGJtO
W5HANGw/XWDh/PJyKnpHQnwJ9g/5+bpm0wbTGXg/L0p0SwVGIQcWxDETb/Z0CKw7
UycsAqoI2y05OkmoHE7KWjFvxGoZRyDMkOyq2+W9bPUf5eoH8201WZzz2Kg0pMBQ
7I+06jmO29FshIzY9YKhTEdOF2ThBbtOxk37avSwtvoNuqWwh0XxZ+78wzW6OMg8
Hzw8to6RjE4cER9N+Q6g8whdeoOiV7iHFazLzGDBHHqwBkG8y5qbWr590ugABHrl
V6wwvQ4K7Vcg1joorh8XTUT4tSWheUzJoxWGf3qCBge8Ad47BzytuM2u14Rvzsx7
IgD1DWkuffrzJ8irXWZiHrQvrAk0yQkLRWgW7sILdX09M1J420CMiXBCrrR7YUSf
8a+lNX3FseYksh6rVvy3REKIigjqtu24oP1ICbSFiR8RYf/Jo9tzmfZ20B2hpk+g
jLY2Obu4gMSiGpyayVR2Pkq80qnzUxFIi/Oo4cIE49mM6aaKbN3GXGFeIs1MVoeu
a6voKyW8QXf67YZ6+n/MRcF8GP3NUQ99Wg/bPlQBuUXrYMzFwsdeeAXCGltfCiDa
Wvgya8tTgpoatgHYRhDxhJVyy5R2smH9CKdrtkNfRuZQXJFMHuq+YUw4HtKQocDX
thqF7CPFsInS7cN78pBgP4238iVt6Zu0jX01f/QY/s01NaGYFis+qZ1RekTj0xd1
gsCcnRd97JSTIYlY+Tf0efX7v3LChczL2128KGudPlsXcKH7uMLC0cYlew3HJIGp
5h8hzOc5Pnr6rFFO1V+k+/BBwuY+9Js15gPpWZzYomHIUpqKCaSQpcuBsMLLc5wR
oZ9vAVAHr1nP83i1+q30a4KlUQpYL5zXE5ZtdyUBkfjp19gunHWxmjX0jX67rPNJ
kD4bU+c2ZZjf/hEJChaVVQdeyk9evqQO4c2Wz0xoTrU7uE1TAqrTeqLhcTDuTRvM
5dukxHbOCY2broEZB0v/vvbQKqrGV1fxZe4Gj3GyodFnx9+hnvIlvKSKnDp8mZXF
2BClM45dEOQZz0oafcFyGyTFC2WXADChtCNx69LcY9FgLS9FmcQuuvs5D0o4ytzO
Jut7yy7knFBphjajrN/nsuFCBu+gl4bK7q+0AXSPT8wHKOYahDHKqzU4xrc/bL5T
1LoA1i5l/zsbXwo3ngGj6jIvy7ux2dL10btcaXOWpllGw93w5KujgNvuPYNG0sxe
yhHC9ypStNZ5ewVD/rO5PDTXtwk770QLl8yikSmbrnazNCmK7h7J8b6YSfUNIgou
g54/hZYCgKrURFEsRQA2ZXWXMUKrSLo69kcV6+caeddPFfCXIIsz9knHc9jFb8+h
Fn7Ba7J79yFa8g51m8pq7NQOmQpolJtGe4TBX0IEN3UthjwWIRLCRiLO6hhjjBON
qU9lRH3ewiCQ6/cHy5kQdjJ/EMwscmE4W2ux8lctpUwb6TTRvXlmfTdfQjGlieXJ
uzxdFErbscSfX2z7o64iMEvvEHccdw+KZEEkiU57r8YMRUmKRY06pAzI6YxIAXwN
Cs7zQ9p7gZAGodzKJoAQ3ypjFX9BJ226bG7LarhSpAM28sZf4+/XURMzOe7zZeUl
K6oGd91j/5c/L1xbxDHttmgXOvAHby1HRK5072ujY3IT8E2A51rA+Hg+ZatCyVkk
w4O2hCs7Cvo1zkZl/XX9Mcsr0pBy/y9NOhtM8B5O27qPJtfigbb1PLi0UieOb4Ce
ScOZT3el0QSxZCTzJow/dSgfl4Es5qjSdjzCE3MhruJwps50AAiGk9kU2xZCRKBw
ILMDbqz8qVvwV3wfPUKPBCaZsTjozDLi9Dx6dEWeRnEiUCvUyvwjo7kj4vXqGOs5
cdXED4pT1ZK+v5BwY96WLNkGHHw8hbUfWGx+mLj9u12ZoPdnGE4V/P/aRhJfTu+v
fHwQxaahFsSjOHBxk5UHJGFSIh7kZpBUNdTdgTgD+GRr11HpfpjU25ufAzKNBrWo
s8Ll1ghKS3FOeqFOVJuGLZHbEf0nXRO+cXAyVXpUfK4RKRz6l9d3hmNT/v5/OwJp
L4QMcDNOnDQpS8V5Ofc07KS9HzfR6mJeLwmcKCo5Xnallg1ahZenZaYvHwcM+nHh
l6ieSUI90g0OJ5G4ATHoJNxqjCmnWHAcM32d5z2pcOsWYImWcb0FR10pV46sHvbE
6XK5cMtO/v0xZpxZPbZIplrKfRWyGO1iIbfqO10OjOJbqHOc7aujfm/X7z9nqeGc
QpLGREEeqKT4Clk6BGc98GHXTEstGcmMXExbckESXaOnsm4jXk/vAkaHzrRUlP6q
NUeP6kEjn8eZ2QObVVav9vlOCV2zBiZIy0h5VUcF//hDJIwAFGtDRyle5f6U/Z/M
AC/iXHwuFVNgOriaLMs7Q0lSha0VlIEsVowPstCcvZWUAtN05EMNIYa98GV2GxLW
p7C6O5MGH2XHDovdDxbFO93LOX5YLVOePxJpGsqwMckV/PzyavdgAO1hH/H2YGZa
S5GYYLt7P8mJNa8wVSkfrp2xferjlOrPeKvyfBYJ/nFfAb+ykl1LY0yLfum/FG7y
8MT9pOc+KZjUxWRkWUuY3neEwQ/LY1yXuJs+NcAqdgKEVdVk0JyUrU6+12WFIye/
dYZsvlF+q5BFoeR1KPdH8oyi1zXqpvwsUHt9ORIuawCoFeDVMwFJJECmajCvNyZW
5LqgR9vRDEuOn11swmzythmaEAPlbxQRx7MoNZzK6wN2SVv+u3IskMcqdUdFbIlp
HKe/EsPI2ll0E0lNeMZ3zpwYeg3NOUuJrgpYUKzKeP+XdihuXD2U89zZDHhL85w9
TpVsOVBNPqyg6fpYg/KdP0Moe8ycTOonQdhvkGGCJElDUKMdkEcv1zQ5kbhIg4Wi
WCE3pxfnTqXAYm8GDJpBA5F2YbZ7LdEtW90dVgT9uxRIo53fvX53LITdXPt4AHIi
TsDk/ucKOiZC0OzKqrpndty8qw52kcVEUdI3o/Dm1/nv+f54dOdFB6O04YDx1Ph5
p9CE4odeHEpGbNDIoiQwlVGM79c5fSo3Yzm+u5TSw39ixBR6Twh4QDjTWUCHJVIC
1itg7QeCI6q4T/LOu+hvaeNCXdSRkZLjIt0kkYxQqksfkHzlVA82iO2u583iXMuI
gkdRqsAH7ch4TEYuuHAiYldUWTvNTouneQLyS+C6/aFGVzhmLGw/hHBZyeugxdDr
bVRHOk8nU8y7VjsTr01iPKWl3X7lf4ShMBm0YxSAb4F1G/PDDE4bkUUmJbeC65vZ
nsw/CclpU5FjH48T7ROB5UpAcLo7KPmPsJJxriGCQk4EHoS4BNv/voKHLwuK11yk
jRAISR691vem7/1KwmexrbvglAF05+jzDkalM5xRzk54l5ItcMoHZusNbd9qDQvW
8w6fYo8zDd4uNnftBJl3JbrV+tz7lyAC/4g9tH6waPtaFtRT5g7bMJjv1/jEhVTs
dX8FWTuhO4KrxRBTg+q2xIGiV6Ix6A5v/QD/LtWhpIOZwr946ujACbXyektEvXBC
vPylYT89mgnqa+z+K5CNgw3ZMlDi+OunVdDGAwC7zYoF+sG3wVRmeoMxhB3kQN3c
UbZgXH6ytAVWofa3v6eRqUBjYet2jGH9NozTe4rDhKdX0KLEPUho06dG4IhVh7gU
46CIFbrSZv4vzoVgEj346G7ktR9S6cJx9c7thwNmPHe3t0C2bbZvw0RHjE0H+QfT
qDtvn946IzgDTQh5avpLyeJvljhzXLb36kY3yCQzBfN/PoWLuBbbBKYQ8uQcfMto
IsBIkv0wCqc5TL5tKcubUPqtMMscu80fIa1AKPLA5eQ0EH0zBu6l8YrxUrGzpQUn
KvJMFoo56IflwFImL/V+Zc3YV338it3Zp6iPKJJ8LQKNw49dIC5sq1GAkp2sACr2
CBldMIroo1qMryPiwBNd3r13U/3UC3/LsCwI7NjGaELyBiMuDZUPzc05chYYuNTV
/bJMv0XahpJQkRVxuES8DBX4xVvem7MMVPO/sAt2SVkEQPOZSdHOMdOpxwVM5S3d
I56UjlXzVh6UPklC4gKcaZcTO2xB8dWZzhIxWcsO4vFRndGnDCRgmRlVIHLpqmvG
VTcAAnlGKK8/0wG2NKOLTAIXVqxEVUUIfPEa5hnWXYSky9dcfVEG4yNwBHNEgKy/
OXiavAEhCq4NMfZC25CkHzJz9ZwmhgH2xNPQfYTSwMknu1h5EjvQN6aQXOBHtELh
PWjXQsDyBWUw+uUP0yzdQAnni7Y4TagzeQJIVAdunUqjvBPgRsP3FLI77dXa/B3A
jmIJRCaUE75v1mfprqOlDOINE6ZRxKF/H1BzuC5sXa6sIia744iHfQdQu0xWpU2g
V/Vzrgfj4E8ithWJpctMPwajqLhf8DZgYx6p2K3Bbhw0jaKS16nBwspCCmLAWQDu
Ajy8X72CjJ6PNqN2oFiK9Eh0k8pQdTa2LO133sWK8gnq2nTQnWFP81nVJyrh2pin
0K276nVXJnD/BoKzKQwEoWwkt61p7W7qM+qplroISjexpxtI1i1GybMEN96HRnMC
vHbjU0oNQ1VtMDnew0qtXwrCr4h/rdxrPWY7ti3avhG/9JXvNVIBs0hp41kD3ivi
U1pbhrqh02RUxSeS10rLL6R/P+up3a7Xbn6yyZItsm40i6pnmhPGwBGMpUCf6KMa
8ADxCa0AFPK+E6xEOLSsXVe6tSCSN+88OsUWKoVY1qfO6WQhePZVYi4Ua/WLO3Ni
+wvSpVKjJA9mdYqSlpQ7X6AuMQKxyBOwZl5cD29Y3LYJX5YAoe+69fBXC69W3MSz
J1wArYhELiUYsjHvCM2r7NXdseRBalhhOmfHt3owSZ9khQygue9de5Zl+VPpbGze
A3by0bwKaFfdqa/DVtojy8rHgRs4qQae6WPlrNdFLi6iNKKu0AMem/MVTdN3BYZP
yZwAmKAU+5eGhFdxkEp5qtPa7Cu/OmjrFatisGjZWeckJ3Sisq/3xhUi74Axmj0S
Ec3qwBRYDHPthVGSI4b9Js4rzk6vWFuNcevo12CeoMPcJhZWCWdzwQ51fM9yBxFg
0eH7yVmMaDlbqBJocYTfk/qtUdojwiws51qiPF3ZvaztofnkfDkpeLETwED+1lN7
tPwe2ACLkSt+Ngp4FCA7m0a+UAwMSzzBmWN8xikK6fajLc+6ORnsY/kh9AXC7S08
rSDzvACDkQUTGzv/F48jJQo8/fIxyEiAh3WVszJ2iV1nEi7LCuqlCitMLWZZRZ2r
R6Bb+ayR/pwoBVY9qAOM8eON6SXCcSvP/w6xMoBUu038ZyLROUyRznHqrDXO3XNR
88dx8gBZhPUgEp0hOnlWGABZW4MP1Z8aIjCXxwJy900JKIGIN4naXlIVyjJpMcyC
Y0vqpI1nPMlRXS7hKkHccHYzKDllHYYEiQ4Adz/CN1gROPaqHxqLs/RVpu48GOpO
U26uPG8/XNyywQSAIg6F0wKEpuQ5qcqwrvIu9z+UPgF9hpCH7UgkBF+3vuRa2MB0
XiDXk60H11AOl2YIDjosfRaVWBzo8y8xZA9SKuUGPSdN6K8wNfAp4YL0KUHj2dST
EPO6awfCiHaR9c5/gx/ykzkl/CiPWbqyzdHRo5Lf2cujSISraqSstxlWtkkr/8co
SwXd7t4NNlr1ZYeuCmmqCGE7cgQ1u4N+Bw8D/JAUDn5bBJLGvCDhwMVe4ipwvsm3
sYKeEEyMFmY6TpTBAtn71XOjbcDY1YvHkaoDVMvH+YJRob9FEJ3MowkhiVBz8Tw/
XewFQC6irTY1OTpUTMJDsdyTnz0xZScotLb8JJtY43pGpXnZrpCkCEZipl2ixjFX
cBJhlJBwPCqxwLXrpHm0d4aw0HweEejj21rx4P7hOXK9ANi63w7AjAVZR453OdnH
B615CcBzFEWSEEfYs5Imd+Ivt+hujKJ6I/p9/r028NSaUiSzDvIgJWKeytQgbWoK
ap0Hoi6eSS82nYLmeH4ntNbjckGBQlacqnzvKFAf9uSIQmBcmWfDyg4eiPkZ63cV
4hQsDZMBxrnTE5hyp1j9+kdZHknqILqMc9dBUMi5eeZYK6MkQA0pc8Y46WVYDSyS
nKLsD+95cBHIZ8989wQBDK9OVdfyPrj+HqB+Tuw00oU25/8TNFQFWIa6CJcn0jF6
qc7OOf5TitV847MAnUvCU1WETBx1N/GjKdoTjqB82/0NOadgXEe79IRy5IVr/eWC
DIJeEFOqiL4BE3pfyMDsLvNfWU4WlaVHyW5GD7xQn1Z8iCBmExfbm/0s0LS/AsLT
Ev9Wd0gqJiuUgZ9YddUfhLwSbe+SHlHQqDQVLTcmDlY5aqvjKzZawJfHEFspveTa
xA+/uXLJ3V7yJa/LkMb+jC4SyGYMdPyPJxzY9FBaoMVrwbhg3dWnyT6QTG/aoJgD
S8GKRu4gC/Net83ftuNTHhwMmq6TnWnS+DNeRIwcvfvfzy0hhILil3UmOAAjvR/Z
LgZ6nee75jq/iItoQYJHCdUwGrEjfbiGK1xw2fchtAz+ExAygW8906CEwp1jRvZb
ti/HkxJDLBcx/YcotUurUHf6VsgAYMNSE2U/6oZtFD7rPcvWKp15bSIc7lRecB2z
tD6lqqYwoi+QhLeb6LL3xEaOY++D+goIp/e1krHbhqE8vQaxnVmlVu6N+1Ausuny
3i40bCb83CSZLF3KCjZX9hCRj/SOE6AgrvbubMe8eb3/o69+Py7dedi8KAfwLNmS
d5bgxzQ91bkcm+r02sV7YjaWN5SXsnht1FbSkCSeAXPR5shFrMKw7TefTlmnDD4C
UNXJxM2P90vkWYllpXU5INgbjYLf+VniX1cEkqJ8eGq19JEzzoPOvL55wh3BkNw+
C3OzDwYqk2H4Fp7/UabkPwLKZN7CcurwqRZ5GVxeYEITCoIHUIvyYOmAjV3Rqq5T
MayYnFcIz0GcCcDQpbTw7xE8vuStt0SPsiQBpPYUAjBflpzdKjA1r7XWvPIoCcRF
s59NdSL8YW0LwaVZ6E4EZsiGdds/sx+Co/YD6g4y7Lq1o09DzdGujv2OZDyJIQwg
JlsdSl4jm+AGWs86ap4kULnWJJTa1ASdNRZ3qqAoz2kpMe0+rWWXsdqjwJ+mWhMH
/DWGkiRJ6rtpruWV6ja+/TuqA1AXdM5UIqgMueqiTEWKAk3/a5U04fPzlknMPN9T
bZSpyhNadsBHhABZPDHefWlvHWW6ib4TGNSlVPMguB+laWJDSj+/HjWNzVMu1heA
HdyP2TUMgmjVQUYmH82kaSgb4zROizqk5+UB1FL+9vAVdivNugnNjjcsKlAL/eKA
6mtZZ2jATYGwaPnAR1kE7yakHaD67vvgN0nOtBiQPVVuoTxrCYWd65gEXetngih7
BDcazza3KQkQL9/yxZlRWKF/UUN6ll9sgEBm14cAUbMUUa4k2EkSriEZRVynMauK
lictN7/vK2x0jNfjFR+NHcPhKJNFPz76xS8xVlyc9Sse1vNhwfIV6k07Oe+akdh2
PKBjwW4rwRJ9iC6ysz7kBggz/9DEA/1sypx9I5y5TOoPS3dirtBDUeiCyIZtZfz8
BrvJcC/hDU9q0HVwKfFk26r8lOr1r9+CY8Arp8WfqBvVwqkmGEtGg9Qo6/7ac3Xh
swviTnGpVuhTgbVu6LwaqLN8GOR1FBPsgzSFz2ZwRxyFR6m2pSlehFmggRcURkdx
aHReYa1CAPVdvQkuiVZxwqI0VxQZcI1HYeTquU1235eOfo+AyvdBSAvo1BOhYDir
fzTiZqqCHJMc7WCpvixZ0LFmrA4b7TZps/bNMa4ckoEL2cner2ODZnlyCb+LSGec
0lCBD52XpEFecZcdoOvuaLiKbYxQpv7sdTAwynsxCPWOmrI0LTDVKIrAK1iThsd3
bDuq8/uod0kwDWkMTLNna+lPo0HKjjovsY4EYCfQf7c7N41xgeQttGmWu4HP1gHl
Acepz1KgxSD7NR6XnmO1K3URbMU+hQnIXW2UHnEMTkkzYxWIJQo6866rFU2OQtmR
VMiQB4jndA+RbOLmUkdZYKXnC346CYYBWiK6B9QGPItXaG/4moPG1l/vdJqgaT+X
tQveJAJshdVDjyx363PlLDEC20DN5d2mKMjwdU8iVmcSTwf3PWIvIvuusXOXTPH+
obz2q0/nEk+m0jZs/LRi+GtwiaHK6xgRGeXjwAfyNqeVcaziuiPyeClnlCTvkjPw
SmRuNPnKR+vGNxAN97oSPNdaIfrHf2eRyzLo2Nswx2Va9fktcJe2RavOA1qD3xHo
W78qrZPTF478caCZP1xLZmuv+tc23OHcOX6zS6Ih8sjYRR1/kDB85DEmh0i6zp5H
K6u64ely6cjUs5/yMxih6hrSDOadGr8Mz1gjmqgcjBU+HXQAJwQMuhSmqrzNR7rK
/+nCOhzm6b6ae4WzUbqDy2QrQyWIkj/D+0Fhya+dMw2dfuCuX4w92dogTwGUJLXR
3WuxUdbtqsxCsLGKFPuNog6Ai8WgPGgSMuWk85JilGSXv0z6vPK3/d0kQLOTwunM
9VyV++vnJwUPtXP97BDIWfbh3L5b8Juc0KRuHX9Oz3rWcwj1YeHuX55UofGsS7+R
dKJ4NxWFbwgdBm1/eTBDu6koH7+Ub/3URDbo/fDfjsYqvEzkUiI88IZC+J4Dut1C
Fa2/o22XhnJYxU8KDT76v27GYBZoD/GjRY2YuRSYjkJZ2RgPwLY37J0Oi0ysvN9i
K2wOMzhck5ARfXytiGZ7QsCoBGDcDpN8r9SWs6lMs9+Yl1Bd8NWccIHpt+kM8BX0
xvfG1Thbfy4MFOuoN0hGRsB2/a3FGtp0gMtK9mZbETXZsCzuz7ls497jGOz18IG7
xaNjM5dOYckp4z+0h7ofbAL9HZTJa5AsXNAnGOjkj6wuB2OpGz3Ajn0iikbScr14
2Ag6LJoRcjCCpPyau1Gh8y7VMHnEpZha2qBj+RwQDQZLU9+mhKAOMKP98ljw9HHP
q6jXOnNeODwGaWuyQMyNKHwZycQm4Xm2sHKG8cxiNmeBWs8Ilk0uZVceK081ViZC
4e4p7RLM/6XQru1qaapFNpUACnL5OBt8EQl28ffYCodj5IBI57pzdPjD6/Uy5H+k
7eZtE/HyZ5RiO3cW2spGxPTvglFiMjGkvWKVHczwwfiAOLI/nOHM7gMY3Q4TD17W
AWOP+IZcXMeKfJ04QmDnWGR0NlWeUNd6W31HzF45v4HaaHCvf0hT3qZf5+BHPNZk
6moyDuhNn1kxVBt7aM9XbLdIB485Lwiuh26gvw7cnWsjMbiPK+gLdkD7de5XXnGm
Z62AnWSvY3U+NajlMB630k0cFEognw3pOfrog7RTJo4FqgngSTom3KtwvGlR8moM
XWxGwaLTtjR2ZsMuOCGm68GjIF6ey2D7ojvmmnY9JTNJ93mLYhC/GzIYArBgNeoq
Wy40zNPc56NzsfEeqOeEgeAJX6ufS7KedJP8KKbb1DhhH1QcJTELCI3YdC2qMnnV
wAmdhp88PDkQHaFeaCPCKNXaDoeE1ff5SWUYxZma9D60rdVaViFOKMg74zailmGO
LKTGd5FSxee1hdo3gtz9UPhtUg+0Nw9tL2iNe3dIjwaBmHIhX0jU5l/VnxJgSFli
uiw7QGVH9ZKuUhHm6bYV0I8Feq0m40yJr0J6xSmssTzJIi2hzQux5jKqvyibjgYp
xPDTu83hxxsgxgGR/ZfWCFjW4VGGC0okj04UvL30N38EKJhzoFWFUzWAS311t+WJ
ia9EBs4mvKHUj0GWpsfN7K3Dblj1ULApfALhdS3SQ7hw8goLTrJsa/1jw0Le+Oif
k74h71zIu3EKeLhuqXZQbavmUx9GJC7Gk6RebqraRVFocLuYJgeC9SQPlf4w1kuQ
yIvmg9eqqETXxdWVnVhdMintLO/mGRsd/x21xlDF+mpcyHTI8oK7tsggWDzV1+IT
w9lWAcqNMUhYLNb3gije/6Z9DrmXC2CswCMWRTwOSAE9XKmvKNkPU28MPliqARJz
V6zGnMfg7DNUaWHV6d9vCb7W2z/MRkJdkHrvC1XeC2EQwBb9ydda1hGRVz0NuUeF
yi4iWQ9oJ4C8H30xRf3w4+5VEsp9rYqO5dzF90/ingXnNHdoqUz6E0aIJu/zLVJC
kxGWAxgVKGmnKcfbnkyFArawDI5jhMe1IHcVoMcw72zi87XpD/G826Mw22wK/FbL
hRK/GOBt43PLjs8U9iUwyk//eL9PEynbl9gPUvlzwFfbvzebSR0ZCR7OavWMJt51
rcpeAeEBorn3yJJKgPKgs86kTw6awEnuybi/Qd+PAuvB2ictQhtVMOkMWtwlOK4C
IvhJmcf0JAjA2EJneOBmWamEocagjzSzUKcbgRL7/3so/0+6zSfXy72j0sSSwN4Y
B9Si1I1/+dw32CU3Nz6nBMlvkhP428ePCLMe8rJZ07lrOQdgE8iWUAiHqfHbWpGe
DiQSMRWngcKDo9aF79BDK2YXQ8HzgJdmeGx9IPy6+lj91tFWJLAhT3CFTKQYPTr/
Xyqt4suGuLLiVcjx7XKnQUa7ZAel1bTpAYlKhmWx+Guva5yNj1IZ93AnjYkt46k0
18gzHIvk3U5b/J0Eq+/5y83InXrZPP4h46rijhRccoe5bgyUv2Odc/+tWDK4Btpb
DyX16VZbtXBSOb7nakWoljOGzs8LBlJ6hbPIBvys/FlUeC/IOVNp3/a7dCGc4yeG
uObbM99mHVAl5z6wfBmi6bEVMEIEpBQqIgdXLPhc/MgPsu8rQK9qnXrueYFHayKS
isufzXcmW1HRNXHKAdlAz3F8IHPOId6SP71CmgfPC27MIWjFu8bXaj2ILa2p8wgh
xJ2QHA7XaxvBPi6eOWf/pgph8PYcsSQw9F0byimw09YjSklypi6YoVSYzOdyQ/RI
8WZM8C7N7NSaR+eNSuhQ9wmkUwKUCvUSDxx3FdZ1r7CuEnndGAYdFyBdebN8KN/J
a78FQn2sz81Wv7nvtix0o6GXFPniiRe1LI5hXVLsoePiZKBWpoj82CGfVwNAUWIN
Ge0VejxPSZE2B00wQMwoebSIAP/vEUjUVxCdbVYOnS5BiFT743B5nPlnEAYLFyov
QyDKL36rS8gEUl5yDUd7vC91FJqVq6Xh7Pc1jSXhZyDb5zb7rg4kBi2rEW/1IksM
faIQ0d0+GJqCq0WM33qYOktNdo8SaWgesoZgcluUb0wXCyG21Y21Mz9z/lIfhlFl
d3hfosrk/PXgvcnwOkDX6S1wX0WcsA+JOVf2QnYDAwHiwguJEaRF/hNCE1M2QKfs
TDEt2QqgkxPdTpvrWCxEpARy+qyZnlnD2eVsub01r7Qed/fkzayurOlfFMih6I89
gZxW1/2N3UGLgQGQbKgcMKCLx67/MXro4SRUy/eU0VNnIvZ2N9VuwQXY7WGl2T83
6Nia2CvMkSiyquJF1EkaN+lhi8JkD25L8AI8RcMq8eo+HpDa66AhhgIS6MXqZHOv
jdxgG32OLmXarGbPGvi1aLhSqcQHbo/GKIzY/8Gnz9jrRLNLlAKeD7xrNs/rNkGY
Tix/a/nj+PS2e3EqBMDVuQ99grzvqY/spI5a6ske0H8U2zju2v1w3GezgSvHYgji
czqyuETebqKxZ4Bwt3OQrudd8fRBQDCBt2wwAGd4QNkuW2SDFQgfHAu534LghNdg
o5yrJ8YIu+nN3jjSbIBY9DVpz4xxpcmhYEL+MyXMJaGv7GJXOeAm7mcNu4vLjBm8
ZRRdA7OEgNYdcMdCeCT14Z3KDvdGJOt+MeNEpRrFTXeOE26wzqVb1zvN2inQwD/o
6MMn7vfYrLEyg26Ye7Ckk6SjOBeYyvpbpVqi/AAYgQ39ckAzvSeqL1+lghM3pEDI
aVfvP8evgg8DUUA05ZaQQsYaTsd8+c8wT8jvC5vg1W62sKUjWgJsI/j5pKxJDLEa
TfS9Kgmhbsp/0y+77RQZdiBF+JmcSQiO6Clt8qyoOUNhE1NQrEeQU9mMxqWlivbk
yLGCqsQIWITVWUH0lqApcXDguFZrSn7+X+noCYTHsVEpTa+xQyL+nXTZevi0efyc
jmqkr276fKdxhi46D1Sk9RHxFkvxSX80at3LZ2sRV9jBAHsTLSaSKUnfYVk2COak
ZrHvy/FHuydG7nJqabQqCryS7YsWQE4Bbcxrz/cGg6fmrDjjnO6K8UDqESZYWIbb
wiNFcW2EZTAo5X2JpUq0Rzpq/sSAqGk7V/djKsaagmieLbkflJj1qYZqVs98e7be
infr8rPKssVtNs8r0FA2fyh79LJGtuccStOLTrgubTq6EFwXRKAUoMDyH6EE2ieQ
2/w8aQx8p9MQjrg5OG/EaMQIebAvJKKJ2hndX/FrCm+qbIZeemjeuXFfa/63DgZl
u1lwZm+4Z6BLTGQ7ZMA1mZxzoUg7JLyK0tGcZcDGAThfG6o8VgdCDDYJ9HxFsW04
c1sMQi3jde/0B9caJ+QBqoWxOnKT7kJPBZeAWySVtq3DtD8/XBR5Iq/0IFzhLl2K
LIb7IiwNrYI1eAmNgtNf7Eg/YNCHEvaSfVTdC8gGg7HFRucQ3mPEz+BA/dCBTfuq
2nM1gKMzlRHh1eFeQEODiXJbj0OUDO6MEoiYwwwJYDaaEQCWvZgxhLV7a+dkDojz
juDGjfA7M4W9McXRrTbW4BSaM+wf+9T7MdnXxYTzNvYwzpKHBs73LT/1kQO9V3/O
pG5oXCKI8m3d0O0NFd5Sy27sHaAOl/OBVViN539Y5yWigDC6EClSzeGk7ibw9PiO
ikRz5E/jybeuujne+lsp0WYnaMhoM9jnLd4Bophn05Csw1AZf5l69PrMq64pI71a
1E/b6Q/bx9J2RYKg+A9nTR8eJMMTlDmMZnedJ/FtmmYjTPu+/XRxJlFhteYktR+k
QHAdU21DgaXFBhcayvgLVtLFQSPf2sKxTSVeiOHwgczIF33I/DfsDaWAaubKLxdU
qfKT/uhAm8lyPDAPcLjWkR5nkob0uSE1w9mmm1n+LlmSgdlO5yizbx3Joxa+lkcZ
RYkhmGk9ncBm1y6hOaqey5eMCjIGKgeMY7H5/58iwrnb9cOsx9FPH+oYiS2MULP4
JIfAg0QIhfN4hKNnZ2wXy4+N16xZ1kfgljtwY+PLeVSqtdAsAgBkJZ9E9mkNsqYE
jDZHXZ87Yb2Rw+G3ypUArJETwWe/OJvwpf6BhAM1QkfR0XsIDnrHMjhjK4kO1SOg
8FnDNNR7oR++55NZdYdytvCvjJDLdF/wqkcDnkegk+QnVdix9X/Q95W2e0rQcEzZ
RyKxQAmk9mCQXkNzwbmoI5Ieb29HdHrKo3cN1OLUasYUi3dVd6krRN8wUMgZhA3w
Lk0Uac4C1Md+Qx1pBIx1+5JV028jx8jk8LxrGWu4e/dXXbRWOdD6pmvLtSSr6GAM
8bjQWWbDgPWAx4iFDtZPQQEWPeiJnwrZxOr6J4E15S6kSIvw84luZ87Ow9hECHL5
HojIyvZ8matb92uHVzL3qcLIMjfeE/tw8ysBNxJucWhFYc9D31Gg5JW3CwmW3bt0
O6vr2wTNqz+a9WbKW63+93LmRm5dMtvKyK59X9IYBNxFZhVGvIAp6Yf064K6STRF
jj0ufvOQlyttC3Jsu4b3rUa6ZvrBQsotWHa7FkTLlQuYFinOFJ8y7z9Xnp/HV4Tl
pOBxqIYwKczvYJSqaEo5hckB6QaUzGS+jkgXEWJMssj92PSWmTSAwFWkMilLkKSY
v7U6pfJQjuh7G4/Do3+2rkOnrv279mTRkQrJ1BYbpIDlzLF91Rdz1XjX5zKz3YhT
r2RML7IRuQl0fGK2qhrMsnwt7fEe2rrG/4+/bbduHmM8B8H4v3+5XS/Ajc6jv5WA
CQcDx8hYfFA5cW84UwOCc96icZ3UdcO1NCzCcarRrfGyO1dY0EhCWwHeHGOP1FK/
DyOdWnEsShkpQYcjusv5p4jdhbMlY17jRN6Vyvo1B/Q5J1rpfKERQSNLggUgp2t/
uZukj4Ja+1fzFTd1ivin6SCiefISrQWu098YGjh6qQd9DVSEh81TLvvocAhowUt3
MhUM0ycxdiQdpMIhsiTCHmjPuWSkSH3CbxAZPAfmgq9bQZy3xdZdLB6k129p5P1a
p6AhhYkaj00iP9CWxAic+edjdtJJsKi+f1oEAz4OhM1YoZ0TNTXfbQ75DLM7KyG2
WpHsLgSSw/foXcGll7eFo6QhNQ4Z4n31IEHX4qXGrz8sgJZxo8a2c0EelILbSIby
JBzBh6SmAlD9Ih5Cd4zN9WbFx3CN9QoswkJ4qr0Zy6GZP9gqRmWHxYT6zF07zSmp
9W9UNH0+1F1Z4Ng5YVaaFuwtu5gzaOYsSO6vtx64EzDPnAMOtmgIgXRSHlGEeV4n
ImpGO1GgYOy6Zv+kYKxoaBBxIQcdVmeJpAh/CaP9W1kg3hWaCCEg4F+c3VdiC7ud
1AcVSDTKxNCM2AAxV74F4dOCz6cjOdLQv3i9Rk+exmZNzhLRG2Agyw3mNyTv7APx
B2RZ/9hiIBMs71Tx030j81NxBLCGRTexsHA2jzJsxQTWA5yvd3+TBMw83JPt3Wgv
GXAPYwy5atGX0UAoq69rgBguRlNXfRcR6jwvpP8nnCYN7n8wYolrtMqKcHJaj6ck
7DtxtSEde76fH6QKQ3pkevdA0xxAz/2dHGjR5GDse7hRMayFjYNbOSJ0KAmz6SxR
ReWbMup9+boQs5EvoImgSrNooUCeIqR+BYIQIO/2evrz5bgJqfJigtX1LW0XnQ1T
76lJVMw3J0C0K9lET/OdSBibT07mLOX3Xck4Uf+D1w/7XCiI7mUfcWP83kB6fkrL
h+fxhojt0UuT01bvJCxCK1GY/mMniMxZUHr8SaYAv3wiaYgTUXmTiFndSj/Vk2UU
w/1r9nSxIqd9k0Guzyi74YTFodPslKgG0X+SHEGHeOZViDALroY6AQ9lZoT8izey
jn5K9QBRpMalpltj94ojXqwdfdAjwXoDepwaynkVtvQi7NsL1+BXQ73NqQIjXnnJ
n/8esxJ9z4gmtGkV2tIcldRmIPvezk0Jqr3uYdoIHWJ3CRQGWI30xMRRhXFgBouL
hpI05zVsYZ++jFIPHkqQPduJBqiWlz4cg/t+oAfD5ChppSj9KiPh2L5akWFwFD5y
jMKdxCZbE6TdcpBeHap9f7Usgw5u/KLUfaxQOuXyx/uF6HSxzhVfijDFwGji96kO
IQyvk6dkyXtXCqotuF7anfgOUI4Kc4ZUQaqC+xH35A/BRapwgV2re+92VigsC78z
eclskArMoN+epvdTIMixYa7X5iVSa18yA3fOHoUC1idRHiq7e11D4h50X++0I+2x
PRVkghI+t//kPsIIUejXnuhLlodYwN9sogtji3xBaK8iXE3Om97f9y2x9JRt7qII
NM1qrT8tpxzLW1INZQjx/vi1IgwN1ftq1PG7u4361/8RtZb0rdfqaXrT4QKrnEGO
qkplEmrASUPr2jrqD8sUX8y1wJL3WP4V27TkQItWkHbyOpsOJa+ncCTcMO8fcrWv
tTBlTNdKyuB3NjOfBnjMvmNGDlAvZouz3cxmVgOwO2nG8BIbr6k/cl2a3clHzzJR
QKkiVgaZ7OT2XryNv22dqc7ri81iAzQZ8KzBeNoNqCgB5zaSVyxaITrJUFSvU48q
bK2MAZdqn4M7JR5mdoS8KFIgrz1qWQpUj3Cridl2yiVLEd8ZVnLuiwmIrWJQ+IkU
bGLm2gL/qHe3RtSOk9YuWcyQUqe1NjtlUhIcwctUKAQTf86q09rANAidJsAV6O89
OoSywfQ1aaoVTbP8Yr8uUSd+hc1fTWsuXjrHUoOByVxaXzkW7bHgpnr6JhSNSl+w
CP8bouSvZeGqEjJgAwRPr0Xu4yMDau5SXB2tb3EkY55jZ7JBOgtXwf09XGDRtqOP
VWJrKSlWeu36a7mcLEsKkD1qhUeRcA4tUAAxEUVdavRsdPRtgy6ciHrB0e7hPc6f
bCJk+dNGciRqC8l5neB0jRtqwfh6fpItaIKKKdk4b19IZvKzJLGoip7hatoBZS+L
+eqR/Yvmur/s7uxbkpPc6ZUhJgSD37LtajeG8K4u38aCWG/NAWmfgJWZlloxWSyc
jM4BQF33S/tU5YWExtxNIcC/tZifi8GrffXSwvprpbrZ7KGEQvLvhu0HQn/E0YiB
DCogFbzIJwkbWqjwXh8jVuKATHj1wkwcYQBR7fqUBncV+lGQwQ+3DlO4CqUlKHOz
14hpPWENqSeI517tPPrq1XbLtg8msao7T86WmUzJSuVJG54N7CX0lTYR6qHK36Yl
B8ow0Xw+boYTzJjlMbfePOte/psaae1LQ9oyDQxFGYVVIIRERVpOKgyAvsV7n1X7
wwx7opVi8Gp5sYiH8rAKBzuLeQTwrOvGOXNHlgLrnHG29WEbiQS8f0fkgpS16m74
wwV/dCsJI94Erksd+mr+oyw6YQD8pGikytfu1jxU8mniE7vT9Ph07ktfXZKZHawg
exDGZNuyNiszm+6EeDNexcUE0p4t19KfP/YlbYAmg89M3jJYOL3smI9cnUs15MVX
SKAKOKdeHsBczS0S7d2z6wr/EH8b55UphbwwdXjHsKiHwoRH1Bx3IiLqutcz3pMb
jvYeCAhsxawT9FtAEXfL41p40bQ6KxZCPzMrhNOviDiygQvGmp+voDtPgyNKMoxK
4ja9mxT8zG/RU3OJoFeTRzeR/8eGHKFo/or+c5zXp0+Vp1Nm+LDu4pLtsRybQd88
XOVgS1A2QZm8Ydw7BtOkCvfbdbffnEqytNrc74T+SZ86HWvZKSYES4Ty2oqDNp7p
upYefw6zj1GXAF7LSquDtHxKW5cH80KLEin8V5epSIPCWTXfiRmzJFJVrBlQ9tcL
be0RNJHoEy3qWB1Y1s+8myZBbscb5uLPUcz/p5DCWqmW/0GInerWMrnq4+9CyqCw
vD2RRo8iTE7Z00gxb6bHJdtXp6RIuIsJHt5e1dCl6tiIY+d24fJ63x9WsWYEx7cP
7CFefOxkO4NPLRAGLJj3T4Art2he/yT2HrNq6Cr1GpgBwjPMBNuVXbH3WP+NZiI/
F8qcBUDhAMyeHn0Un4M1dTf/MXhZil9y+J7VQMpcUx9KogaYxzSfmCn8XfJ8Bk/R
WA9Xsldki/Le0WBBd//+Ky2rnKRKriGZorPWd5b0ajmNBbm4iFl1BUXQ/cU4lAqE
MOsVakCyqUDzpqaEWVxYPWZb+ilHeYc1t2NUWl46GrcZZLSdVnaxX2X6toKHWRe4
fPM5MgtgMWMlnGTYTaEaQz0o58R20QxGNzTBnvqmZrEG34wU/6HOE2IHf7hgVjWQ
3f1bq2z/J1zNTvYvuoDmi8G03RmLOHUSAcgKStaxj3pczrleq9hAnq3gOJw5sUW9
HAWUreKRJDjbo/T//KSEy4jP5twI/Mf80KsiO0Ut8TNh9Qvz4r1EUdaT1wg6AIA7
QoBWfA6uNcExQAFau6focsM17R82Zd372t+N7omHmZRu8XOy6rG2aX6POq4cGLJV
jVDjTkW5C4nTGza0pL8cK/HVAnoEVj1gVFwmkcM6wsaupkgjPkaTSc/hQ7OXa7pa
e/eX3tPvNwMENcpwGyN539w557bV1zJ16xRYubwB5CUkwOk216nILWvFFkiiTAg2
sdgDV9JF//yM8ICKld6ykmO7jQA2QHMiAlkmgGl6Q5ulPgz3e5P8LFoUI/PTJhPR
UoT/prb0DhkRio6ItN5UranhMPKE6dvclnYaXn5gIyExSAlnALmygiSfP8tF6mLJ
rSV9g04H2PW9AzP55JOK3+ItJeepuSsuP/OQcKjZ4Fc8DnAsqPvQxrAcYXuGt9Y9
b5CkQTQcgd9KwrtWIzVpZT/uLXAx0VziIOON7zwCJ4p804oWePI47FTnwDITLdhZ
kL98uF9nFNZ8teuY8amewh7si9ygq8ajTee3jCRgR66XKu772t6G/cLaQ5mQg8Qy
x1W+yUmvPTVOPkOWmeKphczfDc/IJ4xwy3ExQ5sjzAlQ1j5NrqoEdguX+1UCNlIu
P0yGPnxggKvW9rGBQ43Q8nLTzKQgnC0bJDouKfXHXKI3eVVqXyhPltlGgdkC9Fo0
ihsCgQoulEJEE8p26CpxT8sT0KGdJNLot3WaPNbdA0bVagZ4k8aSGznKzxudiLls
IJgJ0n4oajuPMv3fdBMG+/CNQAWJ4zzxaZES69ofBVcDZg/kckLnCXVYHU/PXFX7
H2fozpLj2BKvpwIL4QDHBxqB2Hv+u41mSsT5oXAcCwgDWDFZ0HvSsJcAldUxMQwO
MCcK+CFdHsxC4y/sFHvY0ZsF7AynQgGIHU3a2ZYpVv4gg54zAhClV5f1AG8oEykh
eLMllpNQ65HYL8Dw4RPMpqkGwYKZrrD9aNVsnBojiKkehCOO4joqsopdVPT4wQQA
yC2NyAo2dpfGWRP5sBLwgUnar7SdFoJmFQ1nQLZwXZ4cdQ07SgO2Fi1IK0zCnqqi
kP26A5tlggSxRwMzVMyKjpmSk76DhHhvp9MZBwLMf9n8jdvTd54qU6goQVMCjbQr
3d+mWRcKF5Amkm5Ugg4mojmEyJ9bfS85xaMLd+cr1WW74cphB8ZbJe4RoRoxuP3D
ah5u0MW2UVxExBGpTohJBU1JV5Zt/8uAuxXV4FhRQ5qHAQqxlSZlnTytzQbW4Z89
PWL8z2vB7DkJf/FuGBZ7DnKaZtV1czWpEqi1WrW1O/VF6AHIwFLXn+ktxuBnXgBt
5ItEGWL40IkL1Q/qWrZ3LJsa+Ep6ZOVHjFgS6+xYFpdUbaqf0seg+2RPBoRLmrTR
xjPiUM5StvAZOLMDAbi9V+eofmeZRaFeJkN/y54Q+Ygji7qegqOZQkYKsd+ZZ7gl
IQHSIj17vud9/+dNr/7MudC9aP3xbbqVkuKGLgMQFQtrRIEgW/MnzciP50OoHpvZ
+yP8vDTeByPrJFamW7QkyPUwslOuU+qmkDO2YEjJOxEi12YyYmLysaYiu8X1Q9Ji
xa42nZwK3NO6PZqtNuMufVGD0UUiCcbCxf+squzBNyTwhcE7iVGbpbQkSXBv43Jz
TKrLDdnCuq2GL2snrY4GRKMmRHM71jdIBVrqqgVgUGTEdo/gvHmmFbeWHO6pxS24
uVuD6kbg0rGLOUJnt0oVoOj32pscOYA2UmIExnePi0dt6eNhUKJhwPLDxnr3c6OH
HJPIFgXRS9ydqhvIDz5QS6RtUy0c5PgvAfMqnKmzntDi7UC7Yie2OfbEiBMA5rQQ
nsaoqlVSGrWQUlz1aGqmmJLH4WiaB1duj9/ZByhGB4P6ZoSoLiA7oYQ0BerceJq0
kYdvIHO2ogYSndD4HbaqJv+mYOxxaTA8YZCtWs0Dtb7GvDkbPZio/NVqSff736VM
2njz31yZnC2BsHEizLe/CuImfIanoMYxMCTb9L1XssnM08a1RzS4VEXqu8ms0lka
4aphYzVifAagiEoIcTK9ZALS1scWfwC7iDL3xnZRc3qnIIyZlnT2NbdG78B5GYwc
eUiLkc8JWgSLGfwD72qULCCo0JkCJrCBVanDOdqcXSBkHagyTDtoVMB9Xe2XvhtW
Y+6orznjnUatLBUAKgg/KLIES+1wKP5qVOOCU6aSJHdU10kUNCU9YhghxtHKNyLD
syxZQowD/0bT0fzlasN58vsBH6/DbCpdZ6VsKFWtWMNxzTrPGf12yyzInVaGNAEh
u9qvZm/Biz3W46NIxjLUfd2zOusojspa4SawsnTBy4sizAFeockvQhnEQmnKPH3b
DYRkNBF/XT1xfehDXl8qffWpk4Dc7CS0AYlofH0IN0jPBwvYg1U0EM1UfxFi1N5M
xgnr7vEYtwMpo/PplYFzIxjYmJyykR5Zlpru0lxyppLHdFL6js2ZbIdZXK5KwOqc
rADEYtFvGauMiZFjEi5gQ0GQXlncIoQ7g/quGoh0u3NrGaSlKDY1YG0Hnz3VQs59
PMET07KNsOIOdk9DxxPpFtGvgYQdy62Qv56fRqE3cD/tFMYU+fzpwkdWusg7kFPd
0NaeOg0osEU9GsquAtM9S+SphJgdeloA8775yr1g6dZC+PtVtjerq+HKQyIEA+gp
o8K3EE7q7Zb/aUYh9W2oqJOHPGxHPddyfYqkxmVfdwsZVu5y2mzD73QjS+kj40PZ
G8xvgomYNRw/v909Nt/w1Drv1xM4FOVro5ouL7jCBN40bpO8M/8epOh3etz9dRpC
5H1iaL6zno8asxEVuLbUcFgrSuquUvDZMhZ/pbXTV/W8li/AZccE9HWbQFxOvxKl
NIQpzUiI823HNYM9380jqCnjGih/TBfzDXvagXqWe6MQ5MqYTCLlnKXwOhIXhJl4
UCJUfFRGLTLskU+U9nrG6A==
`protect END_PROTECTED
