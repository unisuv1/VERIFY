`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ff+1vPfrdeXYUjMxBFS1T2t12JfPpPrPSmmxaDPJ2Fiwyuld7NZ8PCaLYUvgEh9Y
x1pw6XJLVjw0Gf5mLwL2uAOsQmSB78GxX/iZ8xRIRUoweE+99gJ2oEyIQLqVo/Ts
GvAupEVHPFraSqZwF3R9Z3X7/+WVja1seO3q67dnzXGU1Z2QaIMnpgkBrUJaWVPJ
xOSpCJ+Y3cAAgIhdl3DlI13/R70H+enHN0mqntg57qjMVuPT4JHTrt9nBH0fP5rS
ic3tBA+2K4nxfeNK+an51DyU3FfqnfIsU/iQZIFN1Y4dxUEVwV5taON1NshcGzWO
J0AI7/bnLZKECvBwTSDwGJ+0QjeBGrWBqn5j96WtjB7SQsNwfQ5bt9De1o7BLDuQ
vn6FAvbDbepH/afcYgRv1eQV0C2mu5nrMyLXO7Pr7fLDxoiRhMVBjuA1wqimLwuH
5Vi+NHBvC+UmKFV4f7Blhf0UsZEQhkPbJeqh9iTfr2SUDnExHHoTuaPB7PwB3HWf
TjMx97b3mzDXT+4fYRc8JLfEqabNXMicMYqHfWiZ509D9La75snoxUhTA834dOtQ
XXazZdJ9v7Xx8e6Opmyp9mW25cczkkfGvWx8VWyE0DsmkwZtmf9vUW6pbG6YDxPr
A4nlhel+txMuRDwO6ngCBSK7zJuMeYeGQqK45JDplU7IUk8zAbBfVbhVq2lfAtqX
liyadMzXohkPWd+4j34xKRtT3vatBek+6dHxwvJ38dgiFfvI+efgOuzMGIq0kjIB
8pqoaMG3GI3n1EXNpvVYIW1w+z5HpfBOpNBBjD2lHPzMYKqUDm85aI5AF57BbtNF
c9mqfprIBLKabS1TK7x9vfllbYmWmz0ij7WR89GSc8s3FkpZXDxyjIoamaI2ekI/
WIzqhusrQ4WApg6r+OCSar2Fpnb3d79tEAD91gzcYNJ6ApdbQBV7NLQ3BTwojED0
PSo7es+gX+UumUA/iMGIOAlYr1pm/fEcJc9IJgNrKlxvKHEZb+DuZCdMFPRiG7OJ
yYX0PGZCdY/WL4VvOkusDbfw1LRovrBy5gohD/9XP1LNG7hZ8sC86FKd+f9kgaD5
R33gCLgHZnHjAnu5NrdlewghbsUlhHb5CweDoQHAjI235yAZxI/VbMyo2/QlzPIK
wdJUbxmMOXNL4tbEluJCJimr8QL6iadI2gpduGsXY5bDFWB6XYT+BfHP3C/BHWjg
85zo84UWyUj46tJNfsQ6n1BUCYRhvYDQvibfxmqNeHaJprnox3ayo/F6zYfw49cW
LFIJnDo/9mkVc4pUG01G7ZzW8e2THxUDykqFfe5/Ai+TKO2C7cB2ZZ7DQRJxEWbT
xnbYtlPnchcJB4rWpE6klmaqzup6g/dVP0AtaF9SC4y6pOK4laqSjDkpYHPCsrFK
MWHK0+u9A5GbVc2DvLgvGBgeGniCJtNdDlm/gFb3QfyIDupfVj65JdLsNrCiGujT
NOoUxu7g3XVs9b0wyjSPNdTt7vg9hZvGKiatRvlsQk1EK4nXWPg0gp3F/jrITy/9
oXBuoolPTOuj+XL5bcQGA6HnNrY08bHOqOYodd3t2UY=
`protect END_PROTECTED
