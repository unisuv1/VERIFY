`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
p4XqJd/BK02fQMfTWr8BLofq5NRdi7pGxHBXT2GD7SpO1XbMfMhqvOvqhshmbKMF
SYPVPJOFkskYgJeLJq+K9jOHn4G5Ug5NyHroOJcTILw3D393wukM9SUHZaZNB/SE
pjvuqKnONglaw4fBuohS7iXxbDlXoVpQeCgplAAeHuel2pYgK2c61FQ96JRV5hg6
kJnTFBhpzsMUKiMnscirpw==
`protect END_PROTECTED
