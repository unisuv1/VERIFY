`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
UZcK0cD6jQrfqFFUM7lu9/luz1x2DXtJExR2EN7TPQbg/Oq/asbOXtf1eaYlQGHm
5KO6RG/VvwtVIhW2TbZNKiSErjQbnLgeEE7AJpoIb4GyPsUnLeTy7cu2aOjkSEHO
pjjmRqbz6zMKg16vYkIcdZW4pYTr9peCK+SDRPSme0AvBBNdIFxhIsTDd3lAOc4D
q+H3xspVMGm9rjGm1Gtq9cN2ezWM4bShN2OHWxw+9iAePjlyKKtwDE7CLiXDn047
wUMW/Vyj39Dk56uJW5XBvuGZrw5LlNVA7SBuoH6l0Z/xIELH5gsM7Eh5RM4sHXpU
Tjo0QtpSB/nt6nPL77nmIqsUUdTPX7K9Qxz7frUqVtnQdf/vVI0MI2t9gW26wUMn
VlvRdIkgZ89+Ie4JNXI09pyrFtXV/X9hVIoCP98pJqY=
`protect END_PROTECTED
