`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
94bcFZXBpsc6nA5uhOSQsd618//59DzisTE2EnilQBIZV/b9/obYnhZNN7QPAgAx
aqXVSon2sekhJwDz0lnWZRBIKicKQ26EJ0LNBoDQojbdRvyIe7RZN9Ec9kc7Z9Ow
oIJi3Hdyh3c0qlS1zdBf3JChYJY7uyD675TP3+ba3IRdeeMWoAcVq/WzYaVu7NLj
PRyx1p8ajtt/6FHaOLjw2e8QYQoVrgJxy/nTP/Z2cYr9wYlt81fjkVylWBzFJpvS
7S6IA77ZWzuoajmDs507wtl9Lqq6plxeqsfmUNrpOAlWRxidBBEJo54AQiGpSMBG
7hUy+Fak4dnqTbz765aP7rffF6cUtR65hTQux7a5UR2qRVCLuKXSY0QHhw+77hxk
D+8su2VKYwU3lqsvIatH0PUVHZxa4tQrUZ4pI11i7OaL3VF3qrS+vwn9eGZPxo+P
9Y3yOXlykl/PflN/mYKHbIqgEjr5ZcehBSOX6lUxNCCcST5MaDHPcGb2kvBss+fX
DA5tRIRvH1OSJYMRWXK8/AQ4lsMWxJy1vLQExK0IAhTHf+gOz3ZjEr6biQiNIQny
oDC+LCX22RYTQyEVOupntztzgeb9hiKOXeLq6TWLutOC4cbn7M/bb+/XIQi4Go4W
X6VteoYDkeityfQecr6NzsAuJtXm/+YxHPwrokrDverRdKNP2nCgxpp9H3k3wZhJ
l1fh93YsChUfQ30YmrIk+eGAbGY+zBa/mkJ8Tnj4jqwbCJ9G4r9R0RpiseD5OC9k
HtTcoiB6si2k4zRAywXi51kQKMKEeGxyACNxvLMID/MgP3Wfi+mVem3AQlzbzeHK
9uDmemful2B1TZgPWGnnTJi3r5VhN32a7aZEqIunIhD6CsaHdxuIeh2iB2O2xzog
xvK/JTyGjaF+BH9Z39opu7J4VHPLeOWhxHJOuBXc8A1F+/DBwaf/eTRADxIldPwU
rYyo71r5iY0foD+oJtagekbHzPZqAsXhx0zf6K6bdLJA47LHvM+tPyPMhaU04SIA
d4FNlU85YvTt2HrXbNxy0UBiE7X+eZTrw5n4J14gzMf1bWVG0jZFB5aa/7dCbbyQ
Tr1ET5q+laMZRvEkH2fdRsk/mbD3lRxH7geii6FbTyLnuQcI04xHxbxSfhjggLyW
7f5bP5/imMqSL+e4/x7pCUFRAWGva6VVrlNXeVEcF3HajHGgPeFboTovTzvZgMZ4
6pyuq+LTyeSLT9ycpoS9jmJcCvg0QESB6rXSqyckROO+QO3OZ/1eT5+acVmjmSRK
xaPO/tKnukyUL+7tvwKgH2G+yT5X5krxv60EITEBUH86m9AkIA2xvSHwmLtrI7ye
r335gM/FVrV2aY1uumJzHSQs7R6DjiKb328jN25l9fArp2fn8x42KMg5QLkL0Frr
0EqfU3cIHho5WTI2s89dojQDpVKm3GyHhB2Wq0p38R/yPA/U01QAE0/O6ZEB+Xa4
s3a0dzMzVlxb/FscZ3to9IEojGAIIJs1/2WDZ2SPZ3+Ey13VCb34dCEPfdCydnJO
M3rZGz/75mRgj87Jh7OJND6LdGGLGcqh9x+i5iDaRcJJcx5qUmv72uMgTNMmOBzI
dJLjd31Wt7hV4546hZ7qsVk4yOJ/pqBqQjGRgbghif3/1Bza/tmqNRTegRLggSs6
Ld5LsqPKFIKj0XTvJlrdj3rc05d0Gutegw9nU+Ue/GFGlrYQpyN1ZffIRxWYJWzf
7FE834n5CwwVofEdTk/7NyfNf2LVAp+I7ew0OPa7nB1QHBiJ0S0A3ks42vg26pkv
Y2fdgpWjG5d+UX/kQKMV6K+e2GlhA/42prcq1VKwPqUgxjSVv8yZIj317W3ZHbdH
TZFVwJTvn6H+AdXKke6lRjpzkSX5ooDQ3g057UxU7ajtPmnVvXs59jLvq23/l3+V
mwWGrIPGnNou1I2V2PeISXV6d6R4XLYELluMyu8BVzPpBv1YfKC7Mkpy4FTMdIDp
jkNv7vzZZhjwntR3F3deu97c0e0rSKcbvG8EUi+CUx2upZi3SbIbfrKQqHKfsk6v
EncNACbvqpeFVzRF1MU+oDFn4KMc0jW7hOcZo6s03uDC67rkZSH1m1utL+rCnrmA
hc35mp4xPXGWZj5nJVb3ioGbAdNzQQMval4DywtlnttWkmPznDXgoc/NcgFJ4hUa
DWZPNhQCZrieDy2TkOu/RrK8GPASl/SjU85AUpqSMh1y+Ue4J54odKhbqnoB04eA
2me1oPlrdlNpdr7hUrsoR3/2pmo7x+u9qSm741Xr2ai5ABXBHahm1jadCYRDLsbF
Io0w+PWP/CHrJ2tDSxo2Gt7DFORpzVFQ66c4d++YPQZ9oxNMoRLDkqlCtVhDgq90
6n/un3PG1D9yhElXjODjLjskvX9agM706huz/QhUiU2962YovbV90xaLw9EhyeYD
B2lTSGT0J6TSOicRDTXngYJhWCtiTmr6otb6KMA1sa5G+OFbppxRjO37C9sxT6RV
Et4DlvLJLE3U7hpRq0M91+lznTrAB2Ic8JDR4rO9b8UsNfavg//ZQ1TRv6b3y/1u
EaDWYmoplNAJxO/PgqDeU0FGgyfTWEocr8zkSiO5LWjrsajojUZDPhvN+5PQhJVu
yeaqrBVgzyxuqMrQAHKpub2ueANUZPNE/cGWz5WeXcMg+hoZzJ66xTkc3DIfJJf8
oSzn9vuhHRL2x30tN97q/JpPiyg//slfyv67kVQPzYMQn5yUH3XBM/xS/OdcGKvT
RqxaXPE5KTzQnqevfI59M6IBuhmgMCqNlfmmRCfWsnNqiXJ8OcDYjHITXow2n2PW
Ctg1MHLKFuIGRV3uC3Iz5iw1pBjd/TrNEn350kPewwknzetlTA8ejHRIGgya1kGL
80xSz9syUeTFudQNM+OeMM4f5Q+TJ/dBahevCcB92mXWaBP0euc5ED+Q9bct+fI9
gYVTeiUxjMlJ2gmEazz+u3gs07fa/MkzsUlTlvIdyMhkwh7GJ3YtuDqjdXSlYnCY
Z0nZr8+oVbB2lfK7rHb+ypP+uGzvyX5pJDUDGre1qMmNbKo7n8GibHKKgWOKNieV
IyyCw9J4VgxCTO3NCd+6nL113vCGcB/fY96tWIzO/TNVFNZYlzMReVrGqkswXqGF
KtYQXmsnRTWtffru03Jc1efYloLyEvW5Pn0St6VWJYe0d1YVhOWDBPP1Sqlmjl94
BDBT8pIy6c61z1K6nyW5MzPDHoEIysdHofXdbfbRJYeQiHZaL9YjhyhOove6ualD
+JEaSaBgvdhjnt5iNdYcjqReOK8LjPxA9fA2bRcZLIAhN1KLvDlRQAZe2Xhw+5Qz
ETPc/ELZ7DJTO84ieNlyBPiPzEXpzowcGhdhMx7qeIPktOCHFcXE1YijnGPCZAiC
2YsPo5o7Xi+KRpMV4gTQ6kB+HzJj41p/ASSbC7fQl9LFxjqcuHrbAENvWGBlz41D
eURUHiA91c7FDmn8ICOohfhufjVlTIRRm6WIpWk18uARFARsh5++3UlZyQgYdXLB
p/lqY4z1Hgrk5ws3JKIJdFKLgGHMWIJTXVd5P8siakF5t7f8EzpfULGLKlErsBw/
g1n8KVp8cQN0HZm6J2YdWqW9tXcZ0HzL/n45H1CKCEEBl8mEfxnrt5JfQyCi1l4O
43k17f1HMDZEYJ+ytGHU6uToiMOdxFzmLFM5xItXlDJ3a4Z93levEITJxU5mdCL6
/WNjXcrp9FVibhJVVdBxmdnscSPgQA3LRohvVI8bWk00HGVJmQiX9k5f7sCmiSFJ
+POZUZPln63281ULkilAKjRGmNGCXZB7/hcq6cPGmLhWWvVeCYOE0NlqbDJDo+N1
8wf8HdrVioRrsrHECrj3+wLFPf27mrQeb91/pfvI8ySpba16mrffZIPfKriKdR+4
5lSw31+bg7R/yz/AwACy5KEk9K11+tZwao2fiVFkW0wbBqjeRzuPWKrER5uHVsTF
W2HmqIPMSoj+4qbhw/IySVJmMaTgqI4/dAoPtXGaURgUyfJIOPFa6qN14COxDFF9
r6BphRs4Kf952nnp+GF2+Cd8tGRlVxAhxgQLIj77bf0Lb6FKeMnADpMlkAUpMMAN
Yn2lc5vLwdAIKxB0p1Pl1EaCjIIX9Bzr1PmVsl6uAFd5GjHtzNJmSBIiSdlgJeG7
AQhdP1uUu2Wp05H1dEP2iYdRu2gl5SGkiAjwiTwJ89OcaUnFuJw0CCurFX9SAnGP
7iKgcaQdjtfmRPjR4QBTuyXo36X0o5Gz3lRx+MkzFBGnFwW3FkbZgNGtHd7Ua513
KSfbDjU9NGOxPpjGs0trN349mWtbGu3PpZEHwYgpiXnaCPqWiqcc6xbmY3BVp/9u
e3oPl+t0JT6PFs0CzIGEV04Kx8KeZmIaDpCfcXTSGNUzGpG1x2VosZxfEmUP9qmS
OYPYETDPyU/xS9/gLZfyUD61LOgckBzz0/vktLwRpQltrQQJV3ITA+vivhebk7BX
goPJjwXlWoeQVJY6bUkToJB7q1MREuWwtXyceBXs6R2mTqRTJk6LUbvZkGJ57H5j
2BqkGHN2aRq5gWKV0dVBULTg62VuzWtrIROpzQmlF2sjho7uxzqebGQowwoxr9tK
XC0ueM0U0GgETC7PP9NA2SSBoxpov7pSKcURO/RgMn7Roryd0x0LJ+dul/ECZZoF
EWk9GAzGMubVyMxYxEeQ4RqHjlUIHETjY6xeJpMZaVL4Nnttxj2f9wnhzetq76zi
ipL0QGezsu52kRqI08Zhlm5pJVfEgS2kbkcbtxSD4WEy40u4J7sg5yKN1F9qrIGb
EADzx8wBBJZCY2sT0Lg3S8tsnGYEJo+p8kr1UksmtfY5PdpDwF+C8HlDkYNNnnkm
FJ9NZtO9uKe5BXyn1qXiYjwAQVi3kml8Si/TwLEgaf0SwkRceRT3UYxiktoHa+aU
CC6sIY8xPdkjH3LmHUXlOBaZsBXeQBWVR5TheMYEasXW6cLWHk88MQFnjn/g5TZc
ekMxUDEqGLz8k5+5o5qSQv9JmcintpjnZlC7LRqftJD3pcwiYLjpbx0a34zZfF/K
0A3Rzj+PptrZPQWEBOo4KW4TekokRd61TuPCq+dwFkMcD5acav+AZHNVa7pw2yZ/
xbko70Wqw+bYzK/d3oXwRgtPouUTuuC+BYECD4ATT1gqMQSUf9j5Mye1XBgTieof
QQ/Y5LfPBMWFeb8Ytnn0+miTqoGUJby8MYZvG1uDw6JcwiWaPqidhWxBqie6dYPI
EL/7Tnj1UxjtTZxBDSw8JWS597eJ5J2pztoZmtt59YKrtORqBNz9jA1hm7j36VJn
`protect END_PROTECTED
