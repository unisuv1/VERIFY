`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
KaHIRRYouml4Dfj+RnQeaimdWsIE1hRvppck8O7SDuRfnAZTsy/rJ0UC17dIlsck
N1QJW1GE/QEXwT2zHNUu8hAWtZXpc90Ncs8VCaQOF7ab1opHuXto7VBAHzeXAg/8
RfjL0x/fi5AmPevqH3Qv+vwpOOjDCX6VcOOryM8bXANm+cyDIOMSSE6U1jTYEM3d
XdxSn6WnmmsEwqyx7LLaqtJCT65XPIpDbWAdcg7upgwNlKHX69yKGg4wYTQVPbWQ
Oycrl26Y/AMB2ujgmkFzoW0iz3Z+om6IL2eMUGtlnn7QKKPNO0WMOtwVghLaC5fo
bOREJax9xXiDzWEHRebsfPpCtBa1Tj0WBlWfVrTP35zVXXS3EiclNSebJoYNmd51
jlRL5kSURHp/exaOhtpFnnbC7/4ROHkWK9WRR0vCkkUKDOxNDUpQKxhHx/KqHrNd
+Ln82Lgw4JPfM1wwpAbqPsqcbyKrNp88dwNFUZz9v1yvw9TiE6ykgFL/N7v0cEfv
jFgnAyDxzEtWDj098CWL+Z/tGEeo9MPY/fcMtnC81yF6AQLARkJt0C79vFRCNGAN
Rm+FuqQECzL/ocJMaNp+uUwsN9Krw0GvWFYnaWdosTtz3dIanJn7gChyrIv164g9
Oiws0bap/BiaPXekRL5kMEm3+53yWQLrSBcnPgFaUyhGWAkcHCTej7fZ7epPpHbC
1wj1NmUHGs1Wr3/Tg6bIMe7Y1SYAIguk1MwnYTycuVSKMf5tou4qDODwAivPUrZa
Ke8M/j8GasUjpX0lUBIQLN+Js1+iv1e/zetwTstlZZu8nBc85JA32lR2NMFTLxce
SrwFvsCOYMTxa4shtMBFcKh4ZhGa08NfGRtl2qw+0OLVTxxIkBh0229fEaYn5Ww+
KtBHsBsMptB+CJijKhoDB3/e22Kl7q/Y6gFB2jvyb52GLFKx4v/jAsZT0uGgDPLX
BO9/HBc0k9AQyDm5LVRX5z15bNMD+3X0ndVhy4NRZYa+ckon2HWgBM0yM0QAjnH7
MEZ6bAnoNupxEbqNu58Q/uGC4gBgnVpYrBPFmcQcVsX/PsrG900Uf3I561ss3iJm
sxXhumgZeKqk7hlriuvdedmNI/HMX36B8gFsX2/d9duCMVI7CZRPMGzQRJFw+cdm
K6+t9fGEHQj5WsI4zUeQ7uGswS/MdWFQJqHdcGMUD++6xHGXmYCSZe0tPLz873JQ
jVoeSL6Zeu7Hv0wyj9egqbjnIq/oXrCWvcuV9WAYE+2H7iWWxkhAcdHmTUL3g9fb
vKiA2r8XtIboar84iive/JTatSyTpfRVE0iPVUBFcnjDT1Ht6XfOT2zCKDdxeJCc
RTM0KX1VoMRkzSTQ+/1GHLD1VGpcyCztxc/6i6n9qHx/YF5Sy6tseLGyXH30mrWv
eylxzMTxPQVZGSeLT8YNaxsJOFhMJlVQrm2v/B4+UrV+CaqeE/xigM7A+rObYqQd
bAGGJQv4Zz22boPeMJ6COIRcqbKNmDwyoXU8BTwhDN4hou3RXON+uqU5bOzc0RmL
vhJEfNt7VzsV5oAXgaP+Inyww6gZHMKHfMXnU4Cs2xxBaRJGfjweqcqq7bAqXi9i
3rNMJb+R93J0LwDzcllz0JNNirQX+jJvbio3spr60vdKkB8rkDBAWxIwppgGr1lV
HxMOWAzSVgTIw/FJpDgVRT+/BVx0vcpnBWrU/zTcJSKRubq3lhVQ0EfxLKZO8jMu
lviXq0iTDTccN4is7tQ0WG7Ub3j1WD8ZZzjv+N8DZsFRYG36TI4BOU6Se99GQviZ
X6aevuIwBRHd/Vxu+727C0pBPnhKsI2rSeg6wrPaaNfFoJdo0KvIe/ia5gs5czmM
BrJf3oyBrkfmiNnby8TbpU+ZSTq9CE/dSoPcAPeFg3EGXVe5VUKIglX5l/dwbmVo
8Wkh2Pex7RXJBzkKVE2+9isqO9u9HaiFXjcfm2R7gffDDj48aC02F+HuceWXlnEH
6PwWzfOV8CKwZd6vxsZhoWNsQs00R+SQjzXPa1oDqKVbLwjzWUgCAkxaP54cGl0p
BVxaqg8UTnxqVAZZyeTZxlhfSDR/zlpaKGCb9IYgYC8+B8cey+ggQ1DUK8VqcYFG
ZuDJ12GUvz9lLF98RKyw5PkZ8ZODos41KB//ITfkN/dP7yO/SpUlEFLftDo51LiV
lB7XuPq+qTUGvHiTHh7aHndvJb52kwzXaTOYTWqMKkCth5AY6XFNkZWqD07yHyYL
/9j5dj102AnYXg4wwnR25LfjH50F3ACTBAqU42ZevlgHz36nHsZHJsK1cXZdq0S4
vme79enluDYNQAE79Z6cXlyh0Vsf3I3K1NSrcBeG6PtyjL+K9UvXDfABIoM53rzX
1/KDqMOsIr9ME812cSM3I/WdEdLCiCUzj3xC/Yu0nSS1ZD8IsephP5JoX2fqk1l/
B6kZqSvNe0xHdW8pOQ7nC9QJ6ZyIrK+5AaOZ+8kPaFj7z9tAPoL/0BhEZDr06x+u
npltO15bOIOvhOk3SSYoCRZuJkdxnIAswsY8oVH+NJQNz9cY4CzQeNjUHcBT5qJk
v94wQaUIEx4ZvZJQADmQytCsD3+OFrWtbf6gTeS9r+lTvlKbENHI9+q+ZxFBZDpW
8xnyIKmwLIAiqkYz8kjfJ47bNSR2MnTMNWwtwqiLk8uSaorQ5FEEAA1ir4K9xdvq
GGtc359jVc6FoziTYOIjN+3FIL7IXD8EqqltG/iSWdPklcShcQoGhNPZK3YLb/Uq
YC0hfn+2hxaKhohRfMyqutdjcUUCn/82zHJ/iUvx2g33H2cflNwogXG6WUrKo/VA
p4yqtmX77lg8IlHxjbsRovkfGB7frl6FZs8E4C7rmZ8IRQzeQhT2xZlEWrgwQIOh
y2cP3J1hCEaZ6ZDZsaIniwDfh3lbPp7RgTSP5/B2NOP+eZbHUyntyzq7WpLm3D5m
55xCg+xBhUsE5mElfoCunhobd6t/6EgCxsxzW14loAAx4g9zYR1yfm39RWr/BuV/
DhZiY38dioi6qH2XzcObjJslR28HSGyIf7no1mAlBrn9UT+FD4o4LSfWU33TGYTV
Pr1/249w+Bs+byJPg9zaXpMHoAr711tE4q6pxYR1YiUDoW+C6I3pc4sti1d31/4n
r4E3hojO9K44dcxMdnojF7BcFhIA/of6TEi88/9zVG0ctaWXZh1tNObLPYUPaaar
asmeTE71JM//DXGqc7qIP3F+Hah3Mxn+ER2Ggbp/9MHwl/dJUCUfglFiba8JtV/7
DGNdyXBXl/td85Nv3ylmnp2oNq8rXQB76vXq8rr7jzzSPvvhlHrZXpDTdhKRvEkz
ZqQuBdHaCo/9io3g/6zNsiitJmQ9qhcfJIs5gtjf9m8sizzX+B60QtBKTFunktaC
lRb+Zk/oG/TEqYT5+nxsFoDY9DNYfg/mPByowFj+4qaVfKQ5EM6+WNq9Yd7stTpn
QxSHw6fswnbJ7f0NvErmDZ/6RaQmyphdL0OwsxXVPZwtG8WMmV8PR3cyZ9PJrD11
GmSDKyjnZlhIPcOCcoWr4PQYPdYevnkOzN+WIl85xvVbYr9WVbT4kGDM/T/0glVS
vgVOYiAbllu1xy19GnPVQE7J27u28SbSLobkKwWe6ClPG0DT/0i4Pe/TsPzdy5VL
0jASgk9x8CvjL6/sDho9M9KDIGAjIbQw2/xN8s7bbKIkpV5RsyzqZWnq/1oPSeqh
gdc3qyMiSFkEmkvmWC1eyldf+YjnE+DDy2TTXH7AyHctHcNPl+kTWfQVJ3UB12MV
YrG2/38L/GVR2JO5eBILM2CgjQz6JeprNTUVh0sNiRMiTzB14OWk3lTjAZXhfHqB
x4XjCfGs9F+LO6g4aH/sDmgjQBcknPAeTK3IdIX36QYJd4nR3USsb87tvMg/i9ch
k+w4bzduoKLrKolzZWgulnxy/9+qH1nUO9uQpXD0S4yN5626tED9DdEF3sqANJ+r
/FmrWq+/CFrkT0AWzrhuQnl68zdy8Un4AJdBoJDomuNpZZ6Q3zrcOKFo6zvCCms9
UkPys7QlIKLIqS4suFpy+El8AhFY+r7sEFY7nWrT7CJP9M9qgereRDeR3Vns5CL4
YD947V4VVNKWd+L6wS8uJGDitPxNUbXXDb+FZ02qrHfhvd/gbAMXWtcvuM7ijM6z
3DUNtqv/bCgKVBFry0sBiCDFETGBfjQzJczPve5vzbAFySxSmYME3/njw+wteC06
1bmGJK3//Ql9RYnvGNxIJDNX+U0AwtuPxYeBs9AwC39/2lUVNwqIH6BozDeOrXBb
gNdYjlURmXAhUNsvwUwYc91EKSbxoPSCdYJWE3SbfX2YTSVkERCknJG/m23qVPwq
f1B1xLPpOGcFFQbFaVBcG89pY8Wjus7SF/yL+5kGk4gmv4zfYYcIGOeudV3vu3Q5
Cw1bXLk9XsZrCOtvrbUVWgRfkXHdOP0XSKVYg5D5cV/d860wxfcZ3UGRhHThFWis
tI3Fx0LZRyC4j+ebpJPj6G1gtXFpulSiwKiH+rQtLPUJH4kb7utMy1auVw4NZuW2
daa41L2ehgTo56sdUAZP2n4MUK2g8oYtF62In2X0qziRziokTcHNl436VAsMYmmX
dRqrbduEgolr4kxTKdm9YUwhP02o0wmmCsqMwSRQ6iAXCdsk2cP/XkPVyPnc+MLk
UGkhzgsnwo8+f2hJEJxC7mOTIWp/9Gxp/tVGl1tHskIziPzcH08aaULokq6X4Gp7
8NdRiv/DuR+PSNc1a0adD4NZjkUmWYwR58/C5fIOTnBUx3d37fXAeMg5hE8sSgmy
aA+4sLvwbxanSyQpm94SNXfAIoTB9OcrC6WzgEi4BOqs601Nntku5m5/egrMPNVh
t/AN0EdzTyciPljl6Hi+3iaTwZjP62NcmN78WMmmFxXLWrLZLT6qsLSc9kveaWjG
mp9dBFMpX/2sCgQvDmxXdqCxdjMEmdwSLF3MnrD0SajEuX/vsq6rztlSASUOIp0a
nfu/IrCyL0pOIY5cri0xzpIP3CYqhPBU5iRQy5emMo8RQcbKn3x9LR1p+Jyl5KRj
FSQ58e0vXqETGcxmtbYsRxuTEVd8ynLulIAkoAJz+viPETmesfbwcDZ/lEAicwUo
cqkaLn5FtWFvO2zXS/ue8tnD6c+e7+8t3gEpKLxNt0LBCW3q/WhVEMPtgqdryycF
NWwxe8dWWg2+q3fPNjstkR53rT24D0MWFB1H7UKNFNSaT3PNllLWkfnSMzW37Ldq
AuUDFVSye887sIH0fJLpcfoLm4aXxK1mkQ2sBteSSKHXtYLkqdIqqPId4birjCD+
Hw9enGDaOLDLbqv3oRZYA7iXB7uiOJ/KHWNDnLHqFvNnoGO4g2RJncFbjypAs1Gk
8jss0IESNWJtqr+//ItnhhD2BRPZaFBDIE/57YF0S17t128pXkYntkOQ8vrNJ6M/
LWvCaQr/aBUwAD+cKskLwJYUAryYCQ0PgHAEcswgpuhbog1V+acimK+TJ+lVv9VF
UeeWVxxYCXfN2kJFW9crLwYgZZJU4RFziT1Ct8JDNh74pTvBncHQ7DBLYQq4Zd+a
2uAoGzVnj1d2KbxQdHQQq+WXRu1qr9eSvnSZMSYRbLH66h0usQyWu+YSB4sTVVmM
XN4GPg9dUFo7dA9C8cwXS4sg+TnxHiqfUy3x1aYdpdNDvedXxxLv1cRJ48dXctF+
DDJWKnP2wBAbiHOkBPuy9OcudVVG8MJdZiw5toNWuAeStM9Xo0a+vuQ9Vr/P3VDP
9s/vAmU2o6NvSc4se66TUkoU9POLmS8saPgFt7UBBr5I2zeV6C7DLD1h0qi6SOxz
EprIQNjAQI6xSTYm+zMcWF7g9wsRsfFoA3A4IUfBvjJt937Dp/YscseRg7zWkZKs
RtGpad0rD6tWH8mlxj03fffViDh9TDd52Y6NlQjpkVUpDbw8ll+jDv8o6qbMf7sG
wc2YU3IIGVm56z2VkLyFxsa7yNEMMMzew7BQbueHVZbHws00Y7t9KnUpSIcvi+2a
qgue2zr0o0zjzPEVO6ZiCHYqCCiOx1m1YExYwTDPG03Sx9uxl7vvrLFc/IytpYKG
0JN+zvB6SR9Taqph+RSY2J3Y2ixzKv1K1ecghSD6yxdQKLqs0kRymsuvoqBAtbgh
c5+wWm0JmE4mukzfgS8aBWhpLgAuMG4xHgIJmOrcuePOsJw4ZHl3e/+mcfhHvlmP
9iwevnwmyjLKbWUgs65Rgwo3JmpXKfKRUbkkqI4ucRJYjapuWvsGaqZ0Semf3Mbf
y3nrc++LOl4+IUnsfR73horf2r9h8hVBiN2/Kgtnrqynu3NUKWvpC7u6u0ox5Zcr
cCpQV2IqJ0jjqxKnt1SZFPdr03EzGRqzJenLTswQ9r3jCRCr7ZBNWYB+m5IqbAxn
+HuGH0+JuGFEostdz757BrjhcQ23E8OVvIXXSTFdYBB9y1XvtI7KHyejBdzLEv8b
bQwd+swVP+ZTNfu6p7qVAnR4yCcfgT1aYKzZfQtQQamK5HngesYdNhgmMGFmQjVn
hQKNb/3Zn4jJt881zM/gLQqcfuASz921W0A1tCQP/QJiiqdPPVqTaovDwgwADl6A
2z324n4QpsQYjboZ3po2uVXAmZHvx37AseSwkIbsztQHkaUpasIMXaQiJ6MuKXTi
U1fRPrFsA0plMlzFTL6W844lSIpKVpYP7z7U1P0OD+xu9UEyDtub6x9Gtwse/vAK
qqcpJzd+gNU47TgjueUmIUzxYQCsVqGvIYarSosqOyNVIh5DNkZrBRcT6heFtpkx
Qzo/r7YWRN+oTE7AnHzc32PoJEBDBa4JpMNMNNpXCbzsjmdPL0UrmsPQBegF+22r
YjLybScvdmkiY+nLz2/717k/oAEyGndzpiR4zDZdYCg7rDOAyIbYdBv+SjVw0zXt
f1y22tj0hCnJ7EHo3owddnw54xrtmCNLAJWEyKMkqv+RdsgmqztBYrl82Bd8NmPK
uwLCB8cnFbVh1+gyxlcJtmNRj1dIbQ16bL179eetI0W8roDwwiSX2J537xPO6JGF
qbcl2R7WQCY8qXvrfcvXr5GM3SHYP2F4gtsHxe7oFm7ot+2Zcnkfos3TVSgnN+hG
VCFj7pzMrcJoxSNfg+Qx7ohDfP6XFBrWlgSdINr5WaOGXLqQaXHUNX0vTwlfCRfT
hVKlTDKGMWDN0F2yCWOL9fDXiuzX02bqzqMRwHtm0FwcHy2JYXRKGFXIvPNumL3T
azUWZj61FtZzImygiEYO3iplzBKR6Yprc4NWRZdP1/dG+UMdFTgUWES59/ZxlyTn
tzNLFY1BGG9Rz0VSnQRPo2hplt6evfhFMMqyKrVNxZvgwmBbSQYGvyWzmVtFrJoX
IB/xkHykcrKGyBgPMFf5mY+gZQNs3R1/78BBgBfNugpGbcfeQg2L9IgWbWC9JNgd
BSAIc0TZVnmd9Yt69IaqhP82c9NC6EKMn6TReuara0TgTy49+4Y1YQc4t1hAi8+Z
uplDnwZMm1vy0cn3iCoudoRivaNzJ3JSFqAYUYYkFTlSjbJfPO+pE95YaiKCnD3D
KgEEY7t1iPdn1p28AmrFu4LVM/xOa2qHvwM6qRQxjk+KL3fBwmsSU6VYSws8t0x/
0Twik7htF5fC7LmxDo9zbf9MlryWFWJ60yw+JvQgqJR3QnnAiIfFXD8vVIA6rIAC
Elz8TG/9fTnCMQFQowVeNqDAmYYeGW5c75w8bl1v/9yiQIQIagkx+6eBalsXlQn+
PZMPD7dt9q+x9MKvdZaEf359MXZD/ZnwO88Q+WLGz2bajIUwddafi3FMr8RUvACe
fIVjsk8PSDlEwpHY2YPNe8VrEvwJ0sBKsFgKU1nAAzgNFchwhllEfNmUCu7NbWgL
v7sdFbDb/CDx2Lex4Dr7Xn7ieoeW7bM202SJ30f4ebPWmpgbTxUjijV7ujo7zKuV
vBjglRKnytXpunbMsnWgsxzIl367sI5PFAUO6GE0I6Ts2gcNH7XPSfaraQ07LfVd
GLHZnF3cyvDSs2En+lC576pzad6LKPhCBWXLSM6ULZwRBeU+xCEf6r0pHjmZaJf6
nUZ03oPIvMo80au3L/Ygcz/ZFvQbIN7RQuH6Fvi32kXrIDS+VnYXulnuAOCJ4ksl
G/UNCFtlt8eNwuEparK5WRukzMsZGEvBs1F9tYHDuYh30hCgT3yLz22NKnWbxZGr
piVbxy5p7lnrI82UbMKyKp2oLdmYmVIRze8vmPIvqt59Vk58/zjuD+8C0SuZ0udS
srNN5FlCMbRewOmwJfjL8E0sS3V5YeRoX/wAp1BzN4Xq32QYEYoFXE8apRKc0627
ya/cJ9MgVBZhX4eLjYsNjnLI+ui9KYR1fw4jV1DuH0SVvRa3yCFtAMeTrdsuU94o
t3UnqWysBubc+RA76Bq8KJ0g0KiqJNZJ1C36+LKkh+9xUpCSqWYXY0tCUBxHleGs
ykjO5foJHJe8VTUIIJ778SmamokSZwlvSZk44d0k3yXvXsk6gG9PU9bvbfc53K7Q
N38p4LnFyw2XI8hr9aSX1uYmtcBAdS4Z3YUm3IH6Yy4QoEAgYF8BtJ6wYBwkOYbI
22f0KvWoGTP0W3uIyRuiU5ndocOy2Hdr91AX6ykitRKCrCY0G6n8GOqns71M1ZiP
hCrri2DibGRtPew9Z73u9ze7jRnJqy6JnK9LSMKlBueJmJt/BOQhF5PhKjeCHYBe
YIfJJ4A49p/1DBfTAe4BpO7Jb6Vtn/7HuJrsoVTv+8URHK5IIZch5SzE7vBSWQ52
/Yv6ix2gx88uwQFUcwC2PaKV+notpc7VECqV9bKpHog3XDJSLuTm//2gImdGcjrr
GX3vXnXKEo07lkYwwH2GwRIdyAlTtZF/D+GEvFiCkkm+EZF4cabFv+zmdP0VWdzg
1kwLDuG+JY0mXvLH+RqL5zh1HFo+onWxNnwS/PeAg35LZBiu5Dzme/CUsqHP9K6E
c+hKtNGkTup00N/FNT/LR5yYzoW6H2DoBRQ4+QabCIkPe7DSa5uEMv2a1SLVgSpM
SGhOoeD7+WWTY3q0m15sriLqM+g+IGLjgmHXeCk3d66lkJ+0UiilB/bQBjR/XQJo
m2HdrD9pYsRTG/SBeHT67crmltZLZ88tEAJNT++cQ61Sya7IEqvFRje1sTW4mXGr
8GGWxgo7pnL43R1BftdX+bhLH+EEWaSlj0vDo/iewHTh/8f3DhoH12NKx8oiPbVf
ClKxEOgFG4cxAv02PTt1MwP++K2zPnsf2Pr+ZI/SRo28Em+V4jRLSh11HRRUQ0wa
2wPEgHr6ZJNb4nf7MEMi4JnvGT+e0uJlQOpjpQOg2wWyoyXpFCyWubP7sLrO8UCF
+yrL/3s4PtnVKO2OJH8DcyYvoAg6PmXX0mxRBfQ95vdcL2Axux+Eb6LOW2hESoPu
n3zUAsrP7e9ohyYhLd5jHOvHlAQ8HPleZRjlfrrTY9vpmkOFL1WjDDFEgXQU/LHO
ycIUJlN/NcnFm/3G+pKHGn28sg4Ob8UDi6ttsKBDBML7W6JMY7H2lA6F4OB2lzV0
aRtRQ7+0H+OdOQEmCBlKZYQr3bli9Ok7TlH7yZtYirg/tOjB09TR9xCrYsro8F34
mrsuQGOCrkne6/Y54k7r8dhc55HgdNih/ZJx7mmg7OrlmkqHxER2bU6M1W09Wwm5
EwY+B2PQ0voohEtK3mS7OikLEROEThYFwkIEvx5nmmx/EmsA+JPIbGTiDGJXP7Ja
e5FDTiArI7Dav9lVy13nLtLR9FhlbghSXAzhZFd0viBTfFGDHmZwETA6WnxyNT6x
94LK/8tZiMnP7pj9JDHXLKZf2mpnvmtf3IX6Yo7usU+Vb34RDH1Qp5n4T8c+4JfB
F869n+N+wRMy80DsUzhCA4AV6UEVRt/w3mEOCLVMqVouErDh+WzyPl9CqIa4uWv9
WURLD848kqZFr/lp1oYwuLiI10D9gp91vAXwNzFviI6TXwmOMWhbEGn0U080UY40
LaYh6opuRbsy2kA8vq60u09d6O5aqOCAKvgj4jG1p2r5qL9kvJBCXU/46pmfgxRV
iS+Lnv9fXUzYk3hDZ+lxuHQi7I03b8VGszP5fQmzB4qjkcxFgUJq4TJk1ukXBh1B
UK5RuB1TgNFdmJAtQEWKvNCQi0QlzoPyqE2eXuZIkcDxID1sBAAi35v5iyQZQeXr
CfJmM5Us8N3xqPt0jAUORc58cQf0WjmOSAjRJntpP5p3pmhUCbHStj7TK9raccUA
3Bbnz0qDc3/7Tpbgq1iirYWiup7ikJi7F9EK+M6+kgma3cKlEcADy1kbQeg2hLvi
QMpGhGVr1rBYc1yOsBpSgmAHQqC8RiFfPQyZH+NenluPTrLCVg8MoTCGyjBn1qc9
LHLIWg+GmA0Z2YevIwHQ9IsSKyT/ZudUJUFUSI3g9PkPqKB4b0n6xIXAIemYfSTl
CxnyWsQ/a7gte2f3H99sLUaNSSVP69KBuHvmybN63GkQmdoDNTtFXbEMPS9Ujv1O
BlS56kx12LR6xBNuvQYbpT0EpN3riMxbgRtjLKcrGHmhjadny3mCaNy4L0K3tvDa
tOf1JFwGa94cjbcxzYLY1lqFK8sAIPW00/JlqVXEARRjYkY7RUDqnxO96SY0x3/J
JWCOvOT4KGJQkPolvW6jzuUcd5jGCJ/8KXz3W9fwvx93QRxuJhzngXA105XSB+G7
TvmRWS/lgHUv/EYFK+lVuoYMguocjH/SzfxIqUyqL5yfh1Q5zZKq+NigOLF7B8eS
bj2aDWJ66ekC84NBuZTgdY82Z1UHEJAFyMe+G2sNQsC0L3aLZ03lB0gXbk2A0crB
S0RNDqxo1C5wjXdtkqRRy66JRi0YAG3yPdbjylm4SDslbedx+xVZAB/3Zr1EI3Q4
zJqBecDJoAlyTv7QWBLRlW/42FwTlFgxoor8Gt0Zgg+BBjQrlBJlCg+t3DXiG02+
lI8f7pcsQOprYq4dJilaK7zccS5Jc7uBOpKarABJ0recXwZxXIs6agHFkYBmteOk
N8EKw1TsRlkNj0K2GDRoh3WZ3/iFW2gmbk2apA/Y2TI/uBRLgoYsJAc8bPBjVX7N
k10bJbGz7+ctpdffEhxtEFOFMwFjID4mvZjWS5biR9sLNoVEV9mUEUGxPrubQrpo
33ebZvkKpvrR/i3/PtRPlpeKeki8v3HQnhjdjkqJuC9RUjOCbHeno1qdkaM9YVGY
LFmsfnc2velJnAaOKl3Otff2He82Dbv9UhpxMC3DTDm1AGh627EWZMtRB5IsOKMH
BXMxywHwhd+pDrGhHlazGwCszg/G3nFGsrOcdT3f4/iG8GpzrjyNk1mZQBVRcwj5
iMmfJDHVpyWPgb0iZKF3H/In4w+0Xdk8VUJuLAeHBR7sp2Rs1Hsq4eIQYrNj7Nnv
6mqGTdznzJJxSAo9mYsqgrKXXBt5QG1KtQl7O5XpVKA7qHnGIyKzQC2RylOPHA31
AWhqfWZ72cVdV3MlK+9da8C4RZVDUn46sTX68sZ4jWCj9lgUNeCvc7cLCPSxFBpX
5o8mRIAtdFsr6jOY+HStzkwgDP+pA+Khv0l9KpWZu5+28Qb/kXaJvRCt1DJ7l1mz
4z9opz1X41ZJeOkf9NiPS64/829rT5B/LdbI7CzQm7N0Khir/4S1j/WZ540Vog6D
9/Az0rGDv4wgevMDQAFw2CLFTAcv/UoTIlH7PFhIecCMPMgIwsgO9MPS51zhKv1S
G5Ga9OaE6viVGPIy47OjJmfW1fvjJSpywMNVISD5jTXdgN98LOny1oNIjsHwW5v/
J7L/fW6dpmIC2qYbIZhZ+UJfK6qwZCNy7tqrR5SYSDxxBk0wLtsagtc5KqRtg637
c9YFuiVHFIUDiD3sT/qR2QBp2TniJAz5haaK+L0azYJMiQpQfyR3WjTWVdvXdoK0
6byChoua8soEG57RVho51pHFQ7Jqa3m0jjRiaMX+W3lhySdTWDNp1a/e3kwg3DyI
qhBoATjDWbX0NAok2PUMOX9QstaINrFwUrva4279M3R/sS8qPeo4UpALICR2XLtA
mSzfLOAyAHumbLw25bwiU+/a45L9AdacZ5zcNAtR2l4S24Jr3wYIXQcYf7l0N0ME
cDtOn43ViF3DE2AzwPmJrA6R6HO9PfWScVJ7X0XkMxkm5otgWdB65ZvunVsuvyIp
lFaJNYxTyU3AjI7b2i+xHqdzRW8459rmKUOFEk3oP6x3U+I7RQtnBp1KTF1ZZyrd
d6fvAb6byUyyIP1nzeGUPK9Axev/TwZ9+TMr6P4ssXZ8jaq3OAuguaa3l3UYdIkN
v5epKU7aghxtcTJaNdgNDGilLpjulBYOZ+fc5kfUPWwK4OuNPJcxazmXRfbO1Fin
4HSXPAURKTDs4wp+R8lOaLzH0cDUr7HzbhjWQEJCxQw9+Y1i2A6DrNkfkiHWgi+p
Pr+MwD1tjst9ZpsrTz5abt6DhaE2Z/dSuoiWZr2PP1DCAUA7zAzDij2M56yzY6g6
5JdjXBVjxAUO/a5hOiTRg2lEs+blcOCYbho0q4pVcaXZ6Wj/ofdelnTmEuunNwTZ
HcA4lIECX0TF7/kh5sbe8DkHtaKpY1HFYlfu49Ow0d7RD7uaVfS2/oKWIdasFIzL
OMbAtW6SWBnZJMVOpThA3CKcB7kIOnTxDGB3IhKAiFjeloBYRU2Wgcr1wtw3oGqm
gzamZ1Aw2IBcFrUFGFNTKFO3y4I7rjClPQadS0VKjhWr+Q2lqPPnkXXW8j6JITps
lMvKIOxQCnKPdTYL2TSb1aWRfFMMlsA6tIHfoS9iXSxpPrFPfB3oPh4fTceEhdvd
7i8gDQTlrD2fDadYYLz2VAIY8F9iQn7+YIvQBBM4gKdhXPfwNydh34s4x9/wX6jd
m4+53Jaq+6PblBy3Ug46gzrcDZUMpnefq6gBeE7hUFyOORWay33dOwgimhozjVYU
1VwakRN0meuV7+iu10245sKTJUyJwOBO1FsyuEaY2fjHOAgV1m10kTXElbZ36zn4
thCqCcCQOIZJG4VzOoxtQFXSF2IZ8t27RDl7MrKJ0ab3cNd/A5RtlzYxVB/9of+n
YDUKwDjGvHvpmDOIk0w/tPzGIbBlZGGcMGhFwEExULuDG94/ZkwryT6iEeO4E01r
vIpeT82vuK/py+yPziqljihzmBLP4Sr18ROUk4sChXFGI7+K/U1po8j45n5Ucg+V
OfMCdwjXqWD6f7wR0cQ2Z1vKBFfTtEv0hWSmLvJm2PSm+OwLQfGBA8LObO36PX29
2vZEyWTCmGUm1etpjoQxMeG7YXo/XRT3frmbYWkytxXPrJRGR5GF52k2qW+agJIj
1YBlsd50Jec76htoNAyzH2ZmXcPgHEgGFU8STVVPu6Np/z8JbE3NOiCjgATFwXW3
x/27LCuehjgmRYbDPCOAg3xDXxNmjghHHyWmMnRYvftYSkC9RQGj7f+DxLpSx+vK
KHliLI4m3Difu2+9XLWReQdhoeuJ7n0paD4k2ShNUs9U4Cch9LeD2BQ50480z6r2
VSKWq7tssX9w+XADNKweIYc8X78EshvGZGM/ycpaQ8JRUhudbHmKaGCLvTLCYxZ3
YQ3Dy7W+ZSNVrMXuJZgzaw+LsBK1hfdOit/etJGaYq4qjPQxo/yMkGLu0jASAF4z
0hwJdOTkchNqnazDsZmwDCfbiwNvs4CwEVpQxZF31Q9+a/azeMWMY9x5QLr8Igdg
hrHWFcuo6kK4GuayjIPyk5z8se1K89xICMogJeJCqkgjpms3GD/bZVvsLjqwTpnK
SqXQVKRwqgCvrIWJdjQdn1rPQTWmF/v8RjYQlzG4aLn+yitNNxzr6GefdxImrCFQ
QEfmACa+YSSMbSOIBU5h8qQ8dsnd8F8iHPKR8sWePYve4fee+9ex7XSexzHWGH8o
an5DwlMt0wuwP7DoT+q2re6yVCQcJHni8XVtCE+StFPFaa+Xa5PH0+01aa5S58pI
NQqySoNhIFplXeSZeaaqCRswuevaj5Gqn0f+lAFqDkYoTJTAp24DGAWzZgacKdy/
CKmlF9xUWinI/CRfBg6yKGzoVPwO62Zf6Jv4PXM1h/oWi/QrJ0iQGBCT0vcvV55W
btHD74y1tXYpk/bVVEbdzSj16MtHKfkSkBeCD3V3MeamVPXz0yVL6WWELl+aPh5W
E8dyurbDgLttKEPqCzUtoI+SJb3kCWPB94uPc0DMWI0+aWCN+a4vwlQSCfF1plT4
EO76voF5HkiScJq2CjVQFXhS2lOeuXlDI+vaiUBxO3/z34udVzbLLtmgymlBU8Fo
R6RloAD3qqZ+xebImYnsptuNmHxXYgsaMiGfI//STHz/Jm8pWk3YoFrAfi1vjxqT
hHqLBCMZgW/5rWraIlkuZ5/B40Acr6OWZ5WeAuZ/0WVAJgYa/Ix6klwXkfVxWNTQ
5pR6Zk9iFrVXaqCUY78oGJuIj52XKkXqcKlrUCgkjQToQG4sIrKd+8VH7BOTt9Je
tiTuU0jPa8VLMXMb3q9yzsa5wUPTk7oBYLIw6kVU26GLZaepjEUbCxrVnXlreytv
4tTUbkSx4k9vnpYZ4hy2GI+7q3z8e0hrb6eKy1m9dmNe57hCzMpqvEvxcJxRE6ZQ
BbQZycGl3N3+WhcwklpNUe+bt/YpEG9R3j7TaGQwnpSsIsZYWhfgolEMm+orTV27
ADDGaMHEcGtq0qOqxAdzDQcmBJ+04UUssQ1G1BN24KFxZjlGwjYogdQMMfw/braY
bFYM55tmhXmwPcUIuKdr0uCSFKRA5sBo1KvkJ30MVG0QplyEVZxgW7mqe1cJsarA
09CRsoksJTO1MtdcaIAm6w8Gun7RxJR6AGtI0Hvhl+aNPIeADvSWbdOpaz6wyxOi
gjOFbN1DVJOyq1fUow9vyOeGtcpX6rO506w36F+ElzMgbWjIr4sy6ByTztW7Lw5X
aIyO6XwmWu57pyYePKdan35KNhRe8uAOhX7KrlP0YLxCuJYMGx34Zt992m+lAgmJ
GKWxy3f5p0SWr8IOSNquxaXVxOqHrN5K75UqRMvNifxUrUvQGIftBpkAJeDFwCLw
+OKq3BU9g86Pgw44ed4TQQGfvDlz5wmfmC4cU7KtVgGY4MKT+rl4nLSav3t4l/NM
vYzUQYvcEbNZSOMTYh0qf7JhtQhLeJfcoOjGTqCSBpJS15o1HlzTIA8G7CzGMIKz
B04R2RWyWKXyu3nmon3tTFgHXmwzedNINKNwSgz5rxrcTQWDpRCd93cgzA0S2Tlr
SjGOREVTZc18O8EUwBdMQLxDQPRz73auDS5Rmah6T+WA03Brpn9cz/VpuWMCvXo0
UNLjuQ+EDMibdXN/lKJiuKQMq4sW6HKZFVaWNO3tZE+CrSCHQ9aErto5pdlF/uJo
8qrWMT5yvgHdlb0IclkCPv4LOA8SAL8B671EhrsuGBz6R5yPCuhIilTTtfr7dYRh
zz64YoFKpjq4t4TC55zqZCniTY35cBy/1w1RBV1/FYFgYyW+talUbZ5Vajg4BYsS
fTR9raPGRfZZB2b7TuFySX1ZO01Sf2ktWD7y8YGGoJb/vTdk1JIhuKzgIHqkcxIq
+IRV11haccG6g8FfcVgeRohppukon5Nncta/E3yNkJQcUQlvKQER9nLDxeAk4B8j
hDQYabHi4342QdaLs9ZYaXXEl8XmPpyUjD+oXjhQoQwS4gULTWa4gfvha/OjlGoY
kFC95GlJ3tKHIDym8akAK7sSXpvEeuf0OsREn+QF5lWyZcCMFfVKN6QjtMBm/EyC
YTxR0PBgl+e/R91VWgqtzOn2L/8jZn+DESKY7si9JWZ3kWcUIU5S+8up0pCj6Z+T
cT8k5pqZ6RkZMWgfSBtqZvsNwfo3lu8ncKlleA4HGc8uK57Pg4s3YKpOFix/LyRi
jNNhM5mLG/EKsjd8o4R2aRqxRu/E2LwrPU1G7LUQwTpEfMFimVMhrQLfk5TjMMM+
c/xoSF85DVAob3wE2/bTYmFqT7IspQ1dOFF/NAqMuXUEkdHSlgR9tpNcl5pIOqW5
1GZe9v7DgcunDwSovgoPuV/dABY287tUZR4f/34g3LUuUdqIkUE2ZQrpFu0Z2NiY
pkDv/6x3nc720q5rYeH/2jXj6gwrT0EW0xaVqd2CpqdO5AV1SyxKG07zJ4kp1+ye
fUTcHULRtShGHSjwk8e5YdWcmM8XUDBlbHxQWnxmZBubwHotxSA4VZ21Px+5sgYn
VsfUVhJZjVn70e/NP8XFT/ex+lPUsXJalUX7dV5XRhhicWREEL4TRedV9mBKUiaM
6uvs76FylwPBq0ZKcexnjtkHfhGUQTs6LzVlgIgIkxb/OKh6uTw1ys1eE4fAhZ9P
ynVl5wI+E7+bn6PAW2+fbSYbmKHcpJJNvKLA72ZL738TTE59D9UtCNMnpEh+KI9v
RiXg1S9NYGs4dVUAljhqMQ9bGnE36q7g60dph7d2QfLQJ6W7sAHOtKxiBoxfhLmv
ouN+EVHOfbX6XPVx6ilZVyykZbi24eH8osi1JTd+EEa6hhNPaM6SFqvM21X0XPa+
1k5pvTdvHZPXZ+PtrZos7AD3qrtwqVkL1TB05fEnyWfKazfWZ3Hp0Km/6G8GHRGz
m5KUzq1TzQ+eU60nk0SVHf4NDbcbmZ5LfOG3Myrsz1GvKMfANI1tcbkNhgMcVkTw
zsY+lOBQxd/J5A/x+9y2uPH4o9PDotTVyBFX/45zkqgxrBVz2PaSUe1XceM8zzbA
uVFUqpxdZJ2erDnBZiQeyPgJHxLL0WsHX8labhtVyXPkbIYunWwVpNfToElutW9m
yGHxVCfRL9vK5H5mHS80TAyQ69ly2PlJMnhEeIkmwPdlQDEw/bNUhLAOFNGD+dNn
e3/uhvrVZKe8cajPajlkUOHoRdDKFfoWwfhRN/uA1uwrE8Q4Yeu499gfsRE/DxCb
g+vXSZJ743cGjtqVeSvyTQc/p8NpWzt3ImoSx5iNxwx6AeUH400GmhTRqrUqjLJ/
zOtpiU5cLc5wX25XevjMkc3ODA2k98/3gvsmlVzd36ofyg2qgAIKLj03rEkbFKO8
drwE2txPmB5nbDGpLrrSRX/OS3bb5qB6PYD8ai2cWTA8D4+bIULq06qD7lzzEtHO
0wJqP0YclUsGxLQQpor/HgJxpjgWVFnYTVYw2uGLvl/5Mjafb0hcHUIuSMR+J/+f
QYqL9uzQB5HTRMm84zwcPQik2/5jjfbTpj4UBvE+GstVE8C2sW0SNnQa36stxBja
WKUrLDX1kvMVAGwBUISCmbnciiEWV5tbu7/SLUWiW986wDK+1PqoAhrSBzLl+kNm
0+1SpekXcmBOw6VESjvi6dY1bLhon3eE1Wr7V3/sqwqeZr2aJY7HWgeuRL9SvLgR
C0s84juhPZ3krhLw1+sukrvLXVVF0MXo0DbNkcSy/0RLmSvjyryprio5WTADdYzE
TakuMaYhEfsx1A96btUFOgfySP6VZkZGso4Y24aYCRQDBiFtrasDDdVQReyn9jR0
t+f+DUzIuGWicwvZs7Mji6Jve34tyIrbTx4AOmVhpmmLNezMkYCrOsmpQpEpwebo
QTzUcI93XupZWXqh38pa64pR2r71s7jR2oB9Y5dNyb2bNFPKIYfIKWVTDag4x7W/
8RC2MQppdav2BgnHsBPLErKkzFl7FeKjUmoAr1Wk4g+A4tl73GsslAU1mijxuL/w
aMcU8DyUJnpGxLon+zFNFYQZYgLrZQScrk5QW5otxsZOHqa1G2S8qZjd3PHLDzcw
R9ochJJWlCpEFFA5PIrVHGRTV2CWmCQ8zZvCXfrWYQ0SsNYqG2yA7rBFjICc2D+O
/HtZVnN6IiVdlmVr+2/Zi326Fo2kQNRe6KIt+OJlECAK39P6dt0qqy3L649mA61F
NdjOUrSQEAVaZXJq4vhWfDt67Sxcfm0T4L+HKNF67BWjyckS8GTxOq4q6vCuG2E3
hh8x+PWOxkaT0EquMRXtU6QbpD2UEASQhYCcm6EUpz/CyOuS/Ysc9sLWOmgIfIKa
ez2/iwFt9GC6ksVcFyI50wzXA3PsRTd9cj1lkwMQRkvivZ+JZxYYhrZUi3mYLOVF
MXuDCYv6n8hqDcmbP0Ms7ssNJzh3WBlEHy/Kqv61xKW8OeG7y/Ilg8y2D5lvR4Ov
HZqh/NMV+9fjb8Q3HABfi92gRqC83qK/4xTJ+s+pZRHAL3RurcfZqmps1wpoytSE
9itgStRV2INiSxFiNb4+eLg35TA/eskyen9XcWznEvydZ8kszTfdAvOvsET1owIM
ujKCaMwnY1DftsrC0KfwUa8XhtywT7T044z/l++xEJV98foZoGrOOnPuZhStNIMb
TW4v1Up3dTgbP5Z1m3xl5WMxApbFZqHvBKyMqosDxk0WZmIh2mFFzNHu8dTokV3X
fwTqWP0iVQeYK1XX/QHYoVc/GFcfj6A50xyTcanp3BEbVUE2dv/93NOv/2JtLQP2
TXiL6VLm9wYqxiuawCEbaPZSMlczMctfMhXfX4NLXV7C95DMUP76clZIVYmSfg0F
EmSJyZd4cIbkj+PcZi44gNa/vWTZrwnStg9b+AAVKD/ACBgcxr4T4mdWhuoQTT6p
DHkqvNbNUDkD4grzyutSN9pzKMtAsudxEvbWa069RC3fAnl0DTQnQ3ta7Tu2knda
vrTJSM9BTHyjnxcsINOc3qafxbuiWNnM/yDB1AGUT6rYrBy+7+WJBL/aXOXRNsvZ
YB5/rwjboXtpG/Fe7RdRT1xfae9Yt78ijx3xgvvcAz6s6xv4/zq6bRQTAJh4dP7D
NSkha0/xeQX0aj5GDNazv9OJmTBOowPQKF4377UyJxhDcPoVn9hZKb5em/FQ2Ziz
xp5fSq496ANMsOwtIzhEX3RUx2Gk5QXatr+PtqjvMPFM4ebQnFUDgRLSjNbYQ3KB
fvef2XhXx0FR3SqM6nXVFCJO1Qgx9KlIGpUvoCxQOPrXbiyfxGHIBSvEFNOSSxtf
ydelMMV+nx/DSmHcRwZu03nX6kDVNW1ekeaD22g8+zMYL8hdMy347WhXIovJIZ0F
dzhUDzICGFt/u+j7HbNpbDIBV0XpOC1DGE4gjMJE9I+bFEQzs70dFtmXqJWcxa07
R/N47JvqexIANuwqfNjzvEKqEjOnkgyEZ0AHFNZSexHjuaeQoT3G8QUE8H47I6h8
JRPnbRKT5TitcJQKx6+BlbMqTWUOJTsOW0sc7qEn8NuyLP/5muQWoGpyNP63tchP
15KubjWYX2GPgzlSG1DXaqT4ZacJnlP/sAUiUQuqkAFGTzOtzGOumpwLDzQq85DI
xyJitBoBOE+m9a1lAGKz4X8YNExRc+qRFYv6JeC1DjAEZhguh51sVq8L2zyoXWGO
RDvJrpfU+LzBd0eWVy7Qpq3Y48JyGM/9R471Gcyf/ANvzZ3ansMCSV8mGwEYeMHh
fp5VJygVNKyH9r+mEhoCPIbt3TdHz+uU16XAO8UbrBv8a8x/L0WWTg0jywV66rYF
QKiJCmmgQL26gw4TIfy/W4tTiYUR4kq16ksFWREPPzllBU5IzYii+4cKOkn97ORN
BnKmUSRp9uWQ08Nb1Y1wxZNj9FR5kCqw3RucJZmD+b9RZgR+cIx6pbTRAid3LCSW
DlpQwW07G1eRDvBuRJLd01W4npcOBYUyh7X2Ra4frlLQXqIjRJjv2tw1YgdvKjq5
zxJVzfucSuwDRVT30VXNzjB3gO0zvV60JuA4ZKzQl9bVmgiP1HaNCxkJRIeHu2Ho
PujF9chyf28FX6bnipYrSK9rPAtq6hayMG4DHWe7dkwftV0570dQYo0tuYlxSaQ/
/D8tTXO0WKMlOrcEWVXIRwXL7dED/4vywcPCnxq67nclnFYLb761pkQLTCYI9hdd
Ax92uNUqvHsuEnjUz5CfaZsobPPS8zTv4eecl5mpwFWgBrd+ce8LurQadnf4gO2Z
AFtqQ7cneVh6XdFOAL3C6UJ18CKVNAO6nBxVaooKtBgpkiXD3DPWkHC+2GxxhUzz
8xaeTYGR+2UE1niBcnofDHqTRYDNK/sIcQNY2GkC6THyuBW70gzSgHnxXHHt5hxL
LR38BGS21vmRmfOIbSTfbEyf2uc5PMjaFiVEv4CbKt1cuqwWkBqkjE6fyW/L3HBp
HZ/1jS8MQr20XBDO3ReGMHQ9B1QPP3QjQndEIJhK+Xf0YIgyA413X+okVh1N7Snt
k6tdUl7itBRShjNYriDNVqiUfp5vYAnt+/5Ww/weLS5I1oI2axZ+pNOiL5nw6j+l
bnXyEUWs3HGfr3M8ozTfqUpj+mch0+WHAf2GshyBCC75/v9ZLFQN7a2DuzwtbCeA
BX3Zdi6JfKGo7lQfPz5cBHzWEkShVI3M9VpUTc4QxYxuK3TCorlwndaMUge55D6I
kqcMyFrFTDTuJFd3bPgUhoc3aILFqktPZRQaPjdmnS4L+O3OHcBFcqF/VXwhgcO8
kVY4OQ8LCr1tgqQVZDjb+8xzcQka0aELvxQ78+1o+gfAVOhtzJ4D9q3Ucj19lrOb
glgrysp4ADU8MoZfBfAj1TCOv1BSyfdufoJT3aBbfa8BthOUIGEYrYsu3v80E0rl
pIqh0D9n8Rie2g8wbzDZWIFnA2bgnhB9EDkG8ix6iLwdhnhSMbWJRDnbEVM7XBEW
nzlxFFVCdow5KI1tA5jLDtl/l8TkV6AHAxTZK955qtdTfF7Qzuq3Kn/cyCT60/Gb
pVnAHx5TWcNLgBgFXx2wrIJ2x54j0fxTelx3+ZjnIQYEKesJ3vhbo0ojP3xvu/rK
M0eA4XSSjD7i9BTrMe7Vbu/68KjtkbezyPePPUqVsQ20cvGvI8SeBbWsirY21GK3
pq+GlhacgXqen4UDq2UciiC3lk6iQ5lmlNN4GixVX1L9Rtz51ZQgx52/4VmjA8qX
9x+4eZANlBWcorKDgKUGokuoA5karH/D9QBMxSRl7AobeG6H/GWBFHmhqywS4Lvk
GVLVHyV59/HTH8eZNvND7xanSKXnqCDQxzIDMBczWK8nXKg1Aw1UPPANYT8zd1wz
rY6vAWfnv1rOg4LMch79uN9iwEzcTBJGiKpg3IXSAZUBi7VGxSxnOSSSm6zDBePo
0/uP5vCFdBAp+ZelnKqWVXW4FRm2MF5exDpb3fQ9CR7Pqgk27LJV0GTQvYjWD1hl
3lPkDAguBKQx6XClHqlrUc/Q4F1mTU5BypMdULzIrn1KD+MNavBXG56I83kM3i5C
JqP9tkdV0gJ2qThUPtzxUb9tsv+bME7jExnkR9QM+w2MS8tx8uYwXDN24FnnnjiS
x5AwVzkg14mPciMEYZaa7+/5bph19e+r60fO+4Sd9nv6UCkQ1ilIO8jBSWxwYQo5
RCXwm5kfurvXW/SP+5D0P9YhlZmQ/D6B4wzjWTdIH0pGsy4QNkk6ghrqrvT3vP1Z
IsquL8+WfjM4C9EPhTBPBF3MLiLl6ABdVchXsiYo9rVvSg/xQmUVwI0I4/4UN3QB
5GhU+eRqZzvImcuReLwO2Q6yDeK3WYfqWZw2IKCvlsPsyvCadcRE0vlTiSHzF35i
XnpLXLoNurDDn62pUQgr4zE07GaNlch2efx4ywcnOTg3inVLaRLLLfS5atx7MDB+
gwvcIxm1MiDllrt/wmpU/a8fXkqAGmYV0yZuiI5sBP06Z+lKN/V6GvjQNSHSlAs/
R3fsAC8PiPN/A6Sr+Yj9YlTnfBZb5KjR84XWWgNmmqRnLYKT6WOQ2+prTFjv7FyR
xthdJhoJ7ZeZZcq1CTiQh9dfOT+kCHqNYM5JZKLoVwk5+eOrnOWSkAnb4boNQSy4
I0/n0EWfrIEgujA2kT0c3CZOt5iUI+wasS9yAioRMsUvsr/bmyvLEycAFxaz+5Ee
TIimsQ+WoMPBt0o9NX6ejix36e6C1i56p1VssLZmbfU5D+UyZ5sU3HvASxWWqPRa
kgA2bVtPo7EXp7oMNMTMPyGhkaVRS/vQLMiIV4kbE5E4YzuEhRvPgaiVH3Uu5nLm
j1nh2WZo3Aa+r+qVFZmX6g9P5HEGpKS0OxNZ2EOt4PvuYczN6ujL+HBk4fy6Fz3b
gheVQhbpmu7gkW+pBJe/XzZKLqYkyqS0zn9+mYkWxpYFz5htJwJfljQBAiT/Fv4n
iLjN/2eJNWz79+uTvXZu0T91hkoJJ/yF+Wt8lYCd7pQ/bZ1GIr2NiIwbJaQuqSqt
3tpz7MkuFD92e3vPZiJrqSljHtkdvuwdZ+qA1RjdAo76lAflFKprG8tuhaLuREk+
em0KBU7rRbyH6M0AkX6EbnNoG69Jfzs8kr4PBU6aUFyHEq7fzaOI3udIb5crIesm
QCbg+faiitAEx/hBJ3I3153c8MlT24mJpFUB3ZaTzK6+ZISh57TqV+EWRqkAAfpC
kA3f42SWm6vHs6H+l8EANFLyIJDUAoTYQE67XZaZqsLxUEFu1HThS58b+bpTbfFH
007W88mEc/NBpk+QRkgdFyE9pUEaMpSoZU7gLVJEX278jGh+tZjYp5XFb1MonEAR
v+/9/Tv8apmqQ7Xh73y8DCik2iE9EwUqj4vzqW7f1P1sQvKiYoxI6oEzSR9Y8c33
oW3L7xx/RuP7OCCA+epQdPZS4MFUzTSzEjv7TD9k/Go/k3gIG1/3sPDxHnYyzH5o
6Pp8uQ/2COy3YHqc/BLovUGbAauX6PL4XdluvPtiJ+fGwR+yz/nEvLQuOcO9Gead
sYZO1BmKL+SKz2ZyQXlXuXDy1GIifyt3wLU4Xlpy7PTRfgVAletBD6XIStIK2/1r
pD4CJ7OvNt6hxuFtaDsqTF/clDsdWIy2TsW91oPP5QMB8jnoKH0DyUV+HGL+lmqP
pRkyS6zDck2aH+4Kj9L3Ir6Ky26WXdQhIFON0EYUBshxrCjXBt/sudKzRwIGedNS
2j+ymrlBc6tDpaCimWzO2AFDOARPZL7szqkNTi9M4UgI23+BGqCHGSuN/SOSnCDG
+KzCVoYeUQ+mAU7zdREqtWWjvXIoAeiu+ZQ+qAbACqXjyHKA3N822Me1iqnswXls
Zm2Gcpu1LPlQSYWSbzKEFZTSfbNDqfD7swDH8a3wGKU1UQ4y8tixZZMIgLm71+r+
YVGqtYNOmEKiA2/BVVL3o4+UHQoWH2VRibaqFYyBfPSQffYorBsOuZmiX6hXpVrh
FDTry4dHRxF8eujSh8sjAAlVhHejJmREgOKljiY5iFMsSOXF8m7CJklbAh1JYHgh
XECmbacTu8yqCKHfaVfb/DrsIrHv591utBLgpFEkDz1TgErl2Ar4EPua28vgRsQt
rtwErjA3r0MEJ2ytxwrEltrC2X9KTOqv+kOc74PJ3ilmzRS7AQZnVo9d9AgP3mvH
p00yQFhC8TBoGNCDEk3csmhS1JVHN8F9jakSLk350UTzH3cGbMC7sS3OUM9Sl4Bx
2MjmY8dmTTfrGjiTDp2RV4yhbRb7SsR638bE5REv5L/p4pkOFDAO7aXquqlWy50k
NeDnkb2j/n5B+Liu3zsKKOyO+o7KbAXNj+53JIhsjX6Luh28+ozWRiDKopMMM/0J
RSa9T6DUAT8kvR6bwV1FH4k3gA+o1IIYE+ipMoRi30DO11QJYS2K7IuZalXVnRzM
bOVDOzsVYzkvU7irlOf4sAKdEUJbpoy6BV6Nedg8KllRWla+8eI/USbVoVD8iggc
Umn+XyQHP61pgGSTmN6NpaqTFoZYvPB1aUOTSoikwB+Lmr/bwQ8o4qIkt/LfX1YR
Ym4+A+KmSzhRQ/67nfNO+p6bQcsGwuuPFpZvgDmnekw5MdBnadiptjaCxXS1PZYu
R1y1yTxvFoy6ni+0tY5kxXA0Fbf3kexm53df8WZjaNn+8LNP70XifZMTsUQN8SIu
sNJaGIbJA2o0orrR0KhQCQIVJxGifuq6AJlN0iTPhNviFBH4chzV9ADURwEquPrt
lKinlFzEZ1k2ji86ZZi86BlSF/1OjhzsCSe/CtzwTZq31TKJdfJs97MhklTW/IAg
NUpeWL23vmKYo7i/WL9+Tgbqde9c2HgQsotvbdZWOyQ1Kek0ZtNUqq+z97uzOu1Q
sPQBPhGXrrRIhPlMCQVBVqJ26Zmjk9IfSVVv2QSj7TuVHjuOxtcal0vm+x+5O9a8
FAsXthbwzqDiFb3WMmHaS5Dch0MfNPhxx43n4v1aMZLCp/insCBhzcS4Gy5sCSEH
CmShPaO1yoWYk9vpr4yp8Of0sYyrk+B+QfoF4xc7FAdMp7UZi1PS9vbgWMZ4fqCw
qo0MrEubnHd1cwja7tCqOzZmFoEmm2DV5wVRyAzmqWDH9m+5/RDwCvB4Chy6jkBL
PXfMbNB3WKTceTUjCLue3UEeJdHNX03jbVc79r8OGe5/1tivK+nHq08+yPMQM5a1
yAAeacQNn9mSzAmEaPsnRtaVDjWFiAwnPtxX2YEUiYO1bYNOEM/RhevfuWi025E1
8zX7+34YpeDd4wXKwUcawubDus3OSROu/ivgDK5LPnjxItOsk6PmaHUVcLtqbEVs
8PS9gUwPAF1uJm+cWw+Vnx8lgoHI1niDJ2Q5VNQz6Nfy01GF0IepwLV9Q9+O87Yb
H2BStl5nJR/mws+zriT03kWjQSUkVsXeQi81CiukMfpMdClKq4/HQFmiIOSL6JYK
FE/KBBTE2rrx7/apPQyFHkhKoWr9MPJhBxrs6hiSjDag8gkxH8LQMI1sP7UeWpUW
o6HQePGJcIEZycLm/rZyy7IAM/7/VaWZTxKctB9JRN1pCb3GrccQS3+padTLRzDK
X6wkVjasdKMss0r4S9oA7ha1lc5hj/SGtko9SWR8CEixVNQDm8PGxOt+f990BqML
L/30uTA8o+vVXVqOOv3IrAZMNkYwvPXj8b3Ct35zQhK8PxugKZNYWfwZwsVKgGZy
e9NqdRXvsS+wZiIvgKYA/9n5gXBFP843pirrwcN/FPF4cH5dj6CBwyYEHt+4jn/O
KJhw2PUH7ITMrXPfru2/jU/h83z3JZxcF5yYiuEmBlfxX7JKE3T3Hgops45hQ3O4
Em2KG6X59y+Va/BMim/jiTSdc2nlTxWTIbb+EYqk48R2YuNQFaHcd2V5oHm//FzE
DcdvoVtUjH4ecEU2ASeC2WYKxKQXHRS7b+mMuP8AG7cKxB0PofPtSLDhIOG99gzL
NNL1dK4IPhffUznkiyQUUK4MIe+jo59BaR02DcWgYFcosj/uNBI0WwSMHcl55BV8
WihEkQx5+3q0UBf+utgFjw5gJc2bxqX+3BfCB6ZHu48MS1FdOEqtfF1WB5IUuZpy
Za8Jy9aTRLLhSrRKAvmFIOMqOLpjjI5tTuvTPNwN7MkzqjhE31ZkW2QC4+J9m+Ps
SOLVoSSFtVkrrW9DfIR/vnQFNwnLPdyvM898u0dsaGVw9h5jr1lq963mo9qwHt4n
R9685VEWVy+obiqAPUIcmzjXKzewwE6p866KmlmGEM7fwiTZvG3hur7adqEY0Psr
avLyM+oYnBscDFLXUB8H7ZEKFT4e/TgTmiCPi8xVBvLqktwdcIv7sraC708jcM3N
og2yEI/sqGk86tNd7LlqFGuz6KK78DWCEzK1d4/08OZiRZ+blQvTf/IqHwaMp586
kVDysVtBYJ5ytxZa6s9voGgMS0hvcs7/tgElO4+VXKkRsNq1spfcwHSA0BAr8kQa
B3W8MSJVut76ipuQvogih3ojhSBM3YcST93Oq5VE2Lp2VAsUcPnd1e/UmzUFEdSJ
BI5SUpdTvwwqLBR6ZAgE5mJGbrRa1q4q2+WIM6UtaVR/dbHvmX8pYRJh27tsEhRT
MYnRAaDaaBa7dgfnEouQS+w6Zdi1LgLQ/b/P9TrLeaOghcxfCTiTuXZR9ipOpa9r
a5kCTcvT01VQaMRvyOHRPhdsJyAHgLiJgWsCVccEbL45CXuNMivTN5aDNBu1lK/K
FRJjiX+pkbPiItIFi2IJBeEDLpmZbYfyxh/vvQ4CFHNDG0lRBmB7NsiTaLOXIHVx
F4Z56lUWuT1H9LqFLFWTfUUzSFIZgTsnXM941CddGA3DAGRTZk9q2EF8M7o8gY3R
SpRFgnP5gWtF1RdqFxqD3x/5vkH0V11VTu1t37/dKk6kCdF7wwZa53WQ7ZjNdpcm
CW6JjJDKMT7XQXeZIpschIiEgAbmmgx655bNwhuHZVCuldb20VqqOVH+8KQ3wdfP
dH6yP5rQuQ8yOOYhoAxXw7AkzFxTiRDnvzDKpmUmchGIE9yPFszTbvJZebKQ88nx
J0F60E6byK8RNZ0GuWSaK1dYmnr1TWYPS/Kk7dtYQMZb34JHQDY/uDwtGTksOK9q
5bbLGaZUAFQJ1CS+JCY1IzWh1SCWFdCOU53ppclsEbDG61mSs6UBzxvToGIjK+JN
E8kI6RPegFZhrUz+Yj5XefcwPlIbBz9TAx37tFH5PRFjwcG+KMWCK1sfOR1xO8JD
WCpU+q91oekVJ1V31ijn8xROvT09SZHoIR/gORPTWBm8ijhsR+c6ACZFvtVxtlVx
hS9qojj33/QbzgCrG+39aY1RPIoPOMAlECOTiKFVkdsqQJyNAwsc+z+oRQtDsZ5x
qI6TpSRJOZT9ept7bkvSmR8nb8kPYzHhg3AASEu6FVirvvcQcHtrWjOdGHIJqEcK
152o8c1JtUgMk34nSS1NooSlRC5TZh8kTurcjJEqa8w1XNIXK24banAl82fa22iy
B64wGL4YVkm3bxA1RMjmBO+vLZRPKWR4DWgXWeYqYwMCL/aG6734yGrSAXFPO/0x
Ig+WZxOKuGc6FYoN7tHrsb2ul+MWFwA3P0JpPhSVy9RZ2G8pEUNvQ/uj3XuQmoNI
PkbHa0otZes3hv8Qi2BEwF6KUIpDT8hhTCnfsitvvRrpyH4x1/3gltsJlOgElXtH
gyv51FVU7BmPUgLOXH3L330re3c/BQOgXA9cl68nq6Dj6HIRyZs9R9J6yIXxYo7p
6bwbTMEcOHuUy6p37uSZWipuMvDMHq5IUmMlVAQ3liDVZgA/0sSlSyJ7BdThrebK
NvB/QtX2ASDGG8m7FKik+iaDdSdz3IRtok1Z1ysuNE3FI0hOJ0fqrBtKQrAgMeJl
BtLt0gNXusqBtbUpjGHfUq0933OJy3KsEa614oos5jD0Llhm1BUSBRChW6/Ceota
B45Ivh5GVjJbuHrnOcvDTYXcBlfdEcHEdWSJFPa0Fmc91E9XECb8oK0LK8XPGE5J
jEENNd4hYX186JPNy8R4f1rRWx2rdLSQNvpQ1RaqlyQmHnnmeUPr8Zw/ZcQAK/Xh
X6TgGqL3POB/63Z+KC/6zhkxlvenJ45+xMiWAallQns36G2lRJqxN2b6SGQ4bZ2R
Hd+eWpo37jD+hHu0ZiDOHTgpnZJ3Uml3xr4A7DmdOV0r2Y4GG4wCOpENBpV+jzLo
n+UvAuxNdIiueL/wk3sHnlaBXpar06vB4m49NwgIuGsPOOaXIsunWX9hIdEWP0yF
ctHvwDdZ3pVBSmpi4XIVlLe0guOlJb4A4XaQYoSNgyUoOrnExqWFfOq7S7lcfxAV
S6ezEsJH61LenaewhoC3SnOPLhGiY+9Cl0UPK7YdN3HqnL8jqa5ZU4bAIm/69gtc
Vsgg9/djKge+u4abmYlKh+3EjcnWAsZARm0gXLa6Ny08ZsAC5pznkrr6mxyewYiE
18Fm6SljuoBtsUwPE7IeHVcd9Si08AhwYjtgCRnh7bsS/vdacMUcKCv/JbiwdTgx
cIrKC9qfBjelekEGfs82LNVJ40kRFgRI+H5xLQhNZiOCn5vDU8XvVOUeJwShE24R
Uv1uueN91BN36Zj8oXJCqEWRUhBXK+Ai2IghHNwDaGQKOhZ3X/FuWtmKv0MmU7YY
Jk3Y3e+b6lUnQWl8c50m2z5A3vYLsHAjDkdUt5Fd08h2yCCIYickZlhg9X8k/Iee
J5jE8zRNvzrABGcgvCLKrNEQyUH3FIVb23OZ1rHmpSt8DN1vg27uI4y//b0Lwu/+
yn6oIzwKAfXK9NEh9FVaLK1RGrj1R9BVp64bCA8JXHEfvrDi7oyNPLiMHMcsq8zi
A/GWgqGQl0jvhbrzj5I7fH/B21q7nN3fjAffLnuigDQU2XinL3lAfu+IKQx6EIDx
in9eZB1JkLY6w52Oy/X8z98XDv9kIbLB1PIXmevb2+re45eAVE7aUveE1Gr5MZgv
ebkyGOhK+Q/h1SXdwRAmKFeAYhgdXbxFo4zis4WJi4zEO//qjb85tB0Hv8YK36eX
AIciM0P9ktSwhgXbbakmZ9gV0wBpPYm8N47Sbk47QrwtLhZqk58HLJvTTQWNWw5K
2pLGk0FmV/t234MAMJCiK0bWwWvF2smCR9tBpYKiJD1/56lLta8GY1qzdgBK+Y3B
F+ys0ldeeuvp/y3nYLHMUgsmxiV/d6lhY7d02cXvxN44djCROjge935mFLjYGVsA
JDUyVvjETA1i2AItiPpMlcibkiiHEmW4BNPdzmdukEIFyDX/gLmNWOiiVc0nIvj8
491GhGV1iSyj0b+jN0+FvkB3hJQJQskBA5At4AmrmU+onsFbgVIqdgKd24sMYuL9
QKBzYms4ULEXTHT8tsFQpn/95ctz0smINrPBtCTN9UUw4R7K7ZwW2eyUWv3So3xY
h38yS7HRo2Y7BHXqq97lNgQ05JMCut8VStf6nQZvybMOJ3FYMh8vn4zfv4jHx4bu
9ikoHBArAnE/MrvIRtD0bj4kEFi4HMgyEpABUfexjYgsgfcxyGKADmV7R730iwS3
7wncH882TJRzOVXmP+x9cGDcpclu888ykp6BBz92S1nlw1jEIoCmT3viT24yhNuF
Sl5luHnxc9+G5YbmIGIvc9C+Bew07YBxxAoWfkK+tEtRMP6KtAXLM29Xte2XYgbT
jbDF8w5aD6jKjOYxVYnQ/IRAsnC5nlrgolEaU9vjwanV3BF/AlbuJ5ziJYQSS1FL
OKP73ax6X/VzMUuz1rC7t5q3V5ByR/5pDKsf7aJteZ9dhWYegNQyWaYfBIwEUmN3
bcQf9a8F/FbddO+jOTrJ/7RfKkjtpRjPxrHaulawjRr1RXjC7H4bUSwFXOUxxtZx
PhUEd/sldLV9QymEu642VIWCzr6rp/AVuDMgNzIN6dCZJQilYOV4D0lWfGp0az85
uc+41FlMzMhCpMSIKHs0FojUQYh2QeR+hJQ+sbvKWlVP0YAcpRtu31ct68T5n8Bs
yBfelGcNi2wmgRCiOKV2sX3j2XiGPy5IrirtEg0CS6qnobab+JbYEFaJIp09yeSR
c/KAraAhyrjvtNc+JKxRe0oFLM9BAv/aq1UpePmF1HJgNuTyJt3uwuMgJZipUocz
sAlCpqWO9QIn5xzw8aWGvRVpNiQ7LyFEVamyLom4e3UbrSIjKsW4Y9OQWD9ilYoT
LnW7cQyrghsVQfI2WHmal7G6POQHpSY+V4HOP1MERHNgHCO5MoAzsD71YwT0pHT7
auuXmkgW/JIZ9x6JPo/MOdM8jMmQ8qoll41h43WElGSdOIEMEjhjzUN9E9ohHJio
VSZF9Ut/pcxLL7wL3KNTbA5vJa4bu3m1XE0vz2zZC6AE3Ln9HLmGgdXsViwS7qlJ
GT876visGv/Dxfog2YUmPQA4lti+jhh376JW1MEM81fASpV3f8Lnz+6YWij9Wf+B
Mq71i0Nrkj5gcvNzZ5mvkFz1xI7Ke58Vjl1giaz3UiV/YKcIZMTCvaHj7hErs8IH
YNrSNWPxFFzPnCiMrOEd0gw0bJsaMLe0fNATPG1baR4OYj6rLPbJSHMR0rT9Zk6U
RSAkSQaK1kAtvGxcVfE+4R6FulowN18cOEUC7WKaQzYk+KmHAI/YEZfLXeNxghQC
65PNDVyX1WRmA6ghT8wVJ9QOuuYQ1XGT/eiQt0FDJlctCe5ce1+jPAjzS8/NAEep
+YC13TEg0nBVSfAJg0weANFi6o+d7jbTJqZrzB110LVU8ZwimVa/Kcwzv+J4lyji
3NmwtU/3uotcJuNJxpBP/uvBx3Y+GKZyQbq92L/XfCeUtlaZuW5IPITB9OT5J0ph
h0xr6OrHRI/KMpKYsxsLi+b1Tv90Ji4fvUr6c7V7OrN1m8mFtGWKU4bm7mXQaeN+
4cAQc3eG662Henb44YontQkUeOHGV5R3hacMnD/pT92xO0qL536TvHwUBfwPoSZd
K7aLsPRtQab021T58CISwXaKY1YL2/v5HEHRiNw++nGL0S/8QodFlqKYE5DCMAS8
/dOqCAihuXShC9AidMs1gizlOKKQxWle8UBDhtmYvBbu7K/n/V2NBOquwU/DMRNT
ThYGJsXurMcOdkqo8z27jfboRU9cyyqF8o1nBWxRQ9K+EaEz8j1z+YcE1WnJ7NAc
pnz1XijWSlCK9XyxMnvil/049mKA7o0lZJJOtc4oRhbksUNdLJs4fjivSUF3LvfP
TKz6VWzQyPpAfaTizv24ANmzHTKBuoAIdWIniDnKFSro0OkClquUhGudZC61Aiky
XuBvFDK8i6Xnyy+eM/kRGG9gZvYvjcIXQSF0TlHwP6tDsE7ilZ/HexBnZUMOyjwX
c3AqZA4P9+ybTySz7UjaiWiGdnrin7VpiG4j6YHxlVAWGScPE9HhSZTyFSyXCTxj
/eTZTIlqcj0y47gm2d6JlTN96S9MLsZAuIJyMymobVeqRylI5RMEz4z5F2c9ZcpN
DVzIENkikDBSGhaECnwMmuED1dApogpMRzbmOAH2G/bBBxKDPxT8S2wx5oMKvH48
WdEI4yWd+N2Es80aJ+f5hzIDJlLQvOFF+d1alzWt7dQCx79nvq4JC12YZjVmUxL1
GZFTQuXfF35TDAkRO6ccuytO+g4s5VP49BM1/OC7uBNWh78Hk9RpSKKCU/cFHZ+L
xOZ9+gg9oXqr5mrjlZ7RI++d6XCrTFSmW/uuRiBTIcdnIvszRE51WZTcukaH1FHW
CYpP8Dd8WdyfFy39kPUFC0vNqRoCmWCE291MTLiK8aCcD3Kv8nP1j+8fls0N3fwf
Rzp+QCX99hZ0VYIFBZHg5iTHoMmcApS1/INshkU69jvGq3CdSIGmSmwTMCQawb96
MHg3GlmF+NHsWAU4Pu6TmuFeMIfag3zj7+qQO5xjdLWHEzbOP7egqapfAn8ZEWCX
RXBZd9lixgrik7myoZDL5pl1sIDlZLYWUSzd7na7yyWQ5Hr/NNZCNCs9HmsLnbp6
sbZIdppSrpmiYh+xY2JlVnqeKWYHwB9de1syrigsfavHx02tqgE60OxGnBSfRoff
NIdpxo9AUlz5UO+UTLHv7lospr9a7wkXSTNaS4DrLNdT42uefrRFTOz9t5pO49S0
AUg1FPRvxOf0F9c/4XkirHYsRIyhZXDoRTHAq7Y7rd0D0EoBJECGVkGwdDRHnGWf
ddLg8N7n5AQMktaFhuqgH2yV+87bm32BeBhIlrh7WlcV01mA0VmMLtJLeiYlRw9U
/X0vLFloCL5KXB1ntR1jbreRY3RGoT7I2MZe89igo7ysQf5NX/tQ5QK6rU/O5fAn
AnD/Q9xTvmIjBV7h7BD8R9o7N0Lxwdbe/kIOEcypqOITqebup7zGSKBW3X0dNcfW
FWrLmkFPkV52/U7BwkxvNNjRYt2L5ye77uCEZ3RRi+SnLay+1ZdmHSlI6IL6PHTh
j2/VxdteYCxGubtQEmcnTYqPtvnykAq/SKWXNgLYpASPOkkgm4tMQul2fOzfEbOM
Rq5LqSOKbOUf0O70C3WkoxyOnKvkKfM1azTxEavUAvDk16CnxtgRY/kTjnO02eTA
kEmW0PCFDsxwlTrUMCAFt7Efjyr2XQQUfLpjPr8CyGRH3JM7dYecRI2QHwR6hbVM
cMSsIXjzPyAlQ+wWgV7yTseHUpj6mMMPv79GvTG0PP0uxo9DnPbC03At6Zbo88gy
TXqOVq/F+NRWQoazhYvXRrDFwG2i2V1TasgK8RRstaPUJiIwOwyMkoxDtxwSZ/GE
Bd9dRHQhlWz0Gev3mrr1NMpWtoZ9dJxOhHfrXSTz1IOUOBXEExUpRc3WryI/0efD
jeo1DmoLqAwp6zRX4C9lQ0sH0p1wCAmLnc3lUBq58ZcjM2tqh99VSq0+zsBCsf6f
mMs2+pbXPZjJBe2VH4hM6YH9tAnylU9Ut+jijYHk6/PkSrrGsqX13W07QAL/PQH2
Yo1O8t6D/K/lRjsmpqmpj1uV9sRXi/SPrLg0x3OMPYYDAIFa68saTYUZmHpIQTXF
hl4Yb3EdzsyuyeOiLZ0nJv1WbcXp1NulTzNK8BQ+ChEhLo0CDLf4B30LUfGIJFGz
dkYMPJ4hqEGIjvcEVDKxD4fSoeIAwsrE7930EqLt5YBaxelkZpVGLpkh6mMQdbWZ
QaPhNDKsTvNt/9JPUVpdcu+7bh0peGwY0s+BWpHaVaAz7Iys3e1cqH/E1ljWWZUq
vKbO2mhBoVFYrzBRyO3ChjAXMsu8BRTUZnmJmQYzzDT4DB7G81tg6jMDhjdhfQ+g
rR5YFAQC3kOFgmPjvqfgfIPyMdRdjoN+D8POco/SsVDrcfoQfo8qYlOyLbD9dbA9
hKTO0uW06z2hJv1b4yWMKwLB0HHY1CZBy4lz4INlkWGre5cvdl1ha+1+UAf71+2T
tttE8f/S1HMAx8sqerG7I9ya7BqevR9Ysb1hKpfbznvnyUl+GH2Gu8dA/UejTiKn
GUdvs2hn+eSADDhbaVegySIXycfZLLuJqH/d51xLaHMpbzMl2G/7AHJzLvmMQDMW
XU7er8KPygCGerwTCjGF4hfqQJNzFD28GKWWyf40mhxDZkLvp4CLQwaFeHWhGUbl
iq21/BeHq9apcPyYEAGmFv3mIcpTp0xaWo735dxv36M6JSgBDMy3TQ1KxeucV/+N
nl0ZG55FCk+PDcH4Oz0nZCPtDlcBK3bn36mKSSUIn0hHBWZOtNizxuHGp2+yPxMt
hLEKqLwH2CGpaqDqJRLdoHUIUQI5T6nBdZwaBBCGiZG8Jkvzpktx48WEMwGYJjke
0F8do0SV6L98ErdpuoyiyojSkvIKAZHGYEj4vnJRHjIM9ufVeQt8n1Qw0NVo+1St
dnCMj7xXn0JVpOJw2aCXpNpBYx4lAz0c/ZcWa8rNmkX4kejFrFuui2GsYeC/B8u2
TCAPcoQA2rfhTtcqfsngclN5mVMSwtroHU3G8aswmdONOGwOYWH7dubF/3SDwG8T
lv0Jyg9UMhyxpWbVJT8FSABaa4oiUnIQQ8m0OHE5EwTE1X9WNPgR8u5iP8mBIxP2
qXSHa45xL+4gJmOFVdB9vZRIvZVwDTtYhdeKeofWmjvdMBacAQPLrIcD5ZG6xAnZ
H5x/bLsG4VVyaOJbUwY2OL9DT2ue5KkZauVJkgygwAoJIt86cl248CQQKYCo0103
tLCRDOOTzpAuNuYb62IcQS5yCIyiKoAN4JmM4GUTlMZGt3XB7L7f1q727mTvW5Ot
1VtSES9cZiI1++YZO48GBdHaecn0/JabhaK+tI58iQnWScQ6LPLv7nO98o1Go+Tf
g5n5w+fGBsBJ2yEUijtveTC1kkWNM7aee22caHyC/LSzhAwkNOcsNkgJVv7SBARk
eOIX/eSXzIC95VWiZpCl81dAHKRWQqDksnrL+1SpGGMXHWqgG/+KbgLS1NG7MPgA
aMWQ+yxJHqdI/rdNOM9CfDWD+2AnMRHOXPIzz1e3r3a2p8KQcObtZP6jTUBn/QAR
MUzGKbB+hU9K2GOOWGHRDkv2yyznZATHzTVw21+J01wNTgYKN4giA2Uy5WeDhSmg
uF/TZmuFlTVIR98mk55IhDg/Cki18Y8DW3GpfDucTHpqt0ovf4f8L2qhFO1nxwSn
XN6D1DIl1qJqUssr0MDjmllA736ReJh7uoEcXBqg7Fv6eBZXDSUCiceC2oq2Wbl4
ZvFj3cxPedT0ara0rtEb5SBZXCcVm9L3z6L7rOHP9hDCvADJEvQgUDu+AGYMT4QI
eDIRWCC8kbSf00TdAZzY/d3+PrMs90eirl2UabarTM6SinC/ufvgenhMBb+zBwJe
O11Aa4BmZWopHG8W5fVJfrSS+3k9iMCbCNqSqYwTJV4aDgWFtL0VoAFvJjKYzPYg
oCPwBaMWqoIKNsNOKTn3C6XcNm/45QZnv6QwUZOh75ef/k94idWeO7R/oCPpeZws
wUhpF1IUj6lmSNhhBWabojiKapf0d/P2aIYkrzQnJW9o16IBwNG794ButjCuziSk
l5z1lS/6WrfQb7PNx465le0jwJ05c5ao0Z+xn20LfEoKM2M46cbRdAoFheeOTtz9
EqPIPWcOaPAtLuBTrFh2XSfcGSlA6ysNPu/plHn4xy+j4t+mmiUlAiyaUA8YiVVF
LMiED7+Up/JHKGhWshNKHT8hwp7d6SIpSSeZSNpvZtdDeDzOQ8x8iDts7xUJcmPN
7e2tldlfnD6QEEUPnfS1GMdZ96gVdE/i8iflryAp9rk4XvQFQF9ohw3bSwhW+AKd
7Len+01odZL6E1pfqxjFqKTsMKOMx/ZYlQ88W7DFiBpsJ2locDGz4NjToufi1Cug
KnEZZLETGFBBQX/PL/FR6tA2dh9TyWbfMchMVkyA6ZImRhLdGE1u1Hse32QNtbkx
zQ6v23RMrUNgNIDQqor30M03jStODvh6+ZKqqVyLkyEuLwH40rrXG+OMBpQgzfqk
WjwGZWYzY72OnPSBuaUDt+FzOVw+JAZJPqCyPS3IEB1ZsBuJ6/aSEbqg2Eent3rm
reP+vfbl8LhzRlHma9ELNOiIkDwWO1YEYMSPoipVuskT4V6G5ZqyqCHsZwchm8gK
1yPpPP15mtJFs5mnb4Qv4KdqLYNnjywoB6dUF34tYUn16n1cVKywYstEZwKnE1xd
v284dDCa/1hXOA4hjJqvAnfa6AsqsYbJiXKgJvwKBI0K/XT8hGgHGPGqd6AFahbj
OYDBB40wC6F7YCnxa4aHTYMFIhbzkR55Fg3iR2noYWkQxgBn/SJvuuy2thJL5Xa0
Ydh3VjkLzMkdNUKoJfVIwO65/Omu5DM5jUNEU1d5sD+Xp7w3ahMedDalLEjVHhax
9LTZ3BEdESlEusTkFJs89bJW3oosa8UyZLgFHU+KbVk+5j4dXDdGD5kbgqXPTrO8
DtMUs574NJYjm+uSCr9ziGhFpF9sZ22Eukp4glRHausNHBeKzx1nln1YvwA33M31
96auFMFTFNYS2aKmjg2aHC6PgFbztuPc1eXH25rAFiEunP+B9jsacP8KStmNDwyi
auflNBiP421zVQ9IzcFjn2mCrHtA/KNDnbuCwDVRcfxe+AhtFHlMnnWaF3xFMxt2
7lpqMwxB0W5r5pMGkx5z5C8BzAXQ0EIt+l44LGVAliiOgAwqKRkO8H7JxqfkzTH8
mSjSy9kGj1GW0zJyMOezjMCynPIu9dKDUuCXT2i63NVKfmZ6SjHdtQZ69PvLKrTe
6KpEo5nvSVRvIj10Q3QyXcqRr8a09rM081gmHFUv0RH1PQGbrM9gwqLGXnVYm/dI
s2oVnonhpRJ+l/BzFZptFryiBUs6x12uxYW6U4I1S9H9cpcGIa9sFT88zFtLnzw7
WPXcl5zao5NQfElNcw1zHDGYky0/FhwlJwhq3E24oqjyGtCMKkxr3smLtnPjU3YF
VP3k+osoT7zvqLE9KkXBUWFTSyJSYxuIPu3ZGRRkrm1TJTeJBFHeuHaS90BA0VtD
0sQSDRWsT2mHYkcM6lNdA3MLxccA68y2pUlh9IX/6jTT1tU3I52F15GQLh+Flh6q
axj2zGkShlqhlJMnApRnDSsPbUs8DYuwBskzfg2HtKjgkuin0m5MmeZ/lF0lYthP
1TDc2OOETCdtTugNa0w3UB/NcU7o/3jfRyIlV65V06vxEmcuKauKSTeGnMcYanp9
J20vanPvAhG/5ImaKwfGKyp6LJ/BiH3Ek2vw2ysCsBI251R0erKOO0rltmqwkv+t
8dS44eK843/0SasvKq1eHdyy8lMJnJpks3PfNiTDUdwSLOz2OKwtssTYxetsQIfw
1X/L25XFcNoHE9j6Zh8PRrxfkaJaCTrzRm0bsn5uioQEuIPtov9wYdA22M8EA2i6
7y/qce3Udz77CGqHTRIVhANKFzfFqNCo394FG3D9+cfbmnLGGseNXo1fx2DsEStf
iy1NGfuBmzjtoTehuV2Tr8GC0FFGUzCfG/P2EaMZvXqQOhdg2DSNjwePCryaq/Ke
Nc7shQVFCGYLzYoprYaIalqKbFCMf1toAhWaLQE9tRuhfLiGLlyxcDiPoufARQgf
bU6tYkyw+QmqwmysZy1MfP6F7U+xCxMGhcorjjRq6FS3DGv4nyPi2NmYvmzovrPE
AZWjGJuubZLTdhcE5iy+C1UgxdJWcVeSbzSsGkBNB5um4jJp+qFSTyRGr4LCJ5vN
MIfb5aIZY08MEi1xno93c63DKwcQ1oncL9Rk3kmla6gMuhEo/BZyKjuL722/6Ocy
k4cibF+H19jPInotF3XWcZ7Wca3HJcD2kjRcZacxnCIrzUovopgKuzZ+IZGPXCHW
USpuV71mel5VwfH+PYopup4BSjaMYWwlDftiqttUTGLzYQ+oTGAfXwYyLFZZt/Gt
cGNMtGRm5FLDP7dv5khvGo00JL8vMoejnuKjtlVxZfBZVq8n/qw32vsEGnhPSzCs
VGdlQiKNf78fsGcGMi3+p1i8uuLg+0ERBNevLeSooJ3UjErs4oDPpk2/mkLdzNZr
KkBcCL2pZTD/+w8MKKua30m9ZoYmWJAZkwqH+dcq0RoIXKaE9ZsEkHpYuevQUb6k
7Vk5F5n/76Eu+pV26TwC7OIf4bG/D1bRrvgQW5dxwopqdH3r7YLaJMCcEGeLxgAF
UqmNn5ydzH9nC8K61oIu/q9BR8Zf0mW02nv2ieFTmt8PFgt6cF0Tl0MxjT8Ts1Dd
mwdYRD0VHKYMlWExIvBC1ixktifiE/a/RM6RDGfnZFBfnid/SU6H360c+/z1wWPH
OWs0ILbVfCuoeJimAp16a+JUHFaoYgMhi/Kog+xhQf/XUfC+XUgy4yTyta+esjKk
Edi4XyplIaI1KzmTvRZ6h9ttJdDM6N4hdkqoSa2+plQD++mgvzju5p7fsg8Fu510
kLVNOpDoHE9YEpVSyDSKlMIG5orh6F+cXarIoME8HpE3Fx6tAZ6qrKBBDqYMuunc
XTifFGe+0qC7yWk8z/CTeFeWkw52eFQfNmZvod9lVaDorN8gd2Qx9jeKfAI2jY+7
9dvOB0nYEfahgoct5uhEWBUgfe98oAFpIsKjiiznbV9ULTFUhSctmznTx9G3J8UD
wM7OvYMI4wKxYAvDJxGzLQ4TYkWxP50yjx5reKf0Z6lepeDrvKP1tinReCpw1iPS
fB+zmFCXMLthnfvmMKfg1A91PoHNDgcjEK30onEF3kXc8e4HGw68eeAl9oZTQ0KO
LrbfmExN5M3UvnB+N4yhEoTowgL15qhMzg6yeYhXvsU3mZJgkYNgBcj+OMa//XTe
hLBfpkV7IRVVKpxlZjJiGdzXvooNK9bDFRx9FYPN0lR2q6/+Zt3GQOLUW71dMrUe
KAJdiTZKCZHNk7j7FD0WZcf4Rs7vBNiSCxk0xW/TGMnZhda/vLkWy+rNFdW9m4Ae
wL7btZndmY47h1+NIJh/6W5sCJ/nlb22Mfsp4QQzM0LXTKDSf58L4pOUtFChWVc4
tTyzzfUXJtXim+J6KtbaJxzsI2I69dRythx+JsGzmw71/f5FZHQVjlVNX4DcUtY4
R9DhxnwRJkypBj0XdGrcNesF3sWJPjrVd1EQrsylS0x6QkygYeEgn+NI2rlBnwRi
+EdaT4r4sWeffP7gIh26cgKkRhZ5BBSH8EzxMhfjFuZRNi/srz1ZeDKYI/jmscSZ
BQS6VXjV6EurNxE039mVqvblkR9F9c8AWqCL+o/TgRjYAiYhPXFMZQjlTcvA0RO1
Gd055YQSVpB8DKevV1nYnYf1fXl8EQ9zfLxebiahgg2jnXTGEj9R29MNsKoiPbBd
fVS95w9vG6PnAfgrnvOXGjMPAnNw2iQJw3DACzQmrW63pKSfV7KL7EV92MXqc1aG
glpcnGcYa5d0pr5N11Tbw2XHGYgBUt9PXhuuB13MDRSDv2hMiURKL0Ys+lFTlL+/
XjE+po3xvkH89wLH4x0PeK8U8E5vFBH/UUyinfL/qq3nmuLOIPQCSIQgG/3OZhRi
34Ip0hqx4/7W49LCyxWBSsAYbDMMqbctUMSZ+Lb/PmQmgsnkxHIcuayr4DRMX7Fk
5k7+GDXrnPRMZ9rJ1s6GhtNMKLTGHk5jzD4c+b/4qIetoDQg65P0g+nhnUP7BL7d
03/KBBexyidLOaaoHFJNV3TgirWrl1k+cP4w1hWxv+tK+0qen3lJAyYVt5AngqZv
2tUQVaBIZKgqmDNsAqpoHhlhTyJuVfKDVY4ixVPLD0zxO/mpDguiHyNaWCLtsvCv
oODsImM8B+/U010u6BEWdGueuJedzLnZMlhVRaUN5Ag7VNK1TtuF40CsQUX0YzFh
ZKj9qeL3nhNgq5yv3ssZ3rL3L5Hza9kWxqGPAZTd4my/3/bteom56YdydJSw8gs6
rAxbJnD2yhu7C0jsVb4sd/8Hv54HH5TgzmBcwV/KpNKLkvHN9f/gRMKslWbhRciG
XRGOuK5JgYpDRMjDwUOB9hlLppoqqyr0eFjofAKEDMsdVVzXkd2zFzgOwK+BBKbd
1HwnChEaobmXluLoxpv6D/2VpcUTTk2CWLE8GwE4lQ9R3s/ezHdBgWXxkzM6fBIP
/zFhcYxyR970QJ4hWdwJ/oPwSsu9QLjjYADFxFmpzaD8/9Aq15MWhF7zdhSPThYa
X6YZjegnfw/kYpQLNs1MQhCEO3CDrY6TwpnAXfEnZJ/XS4Nzp+Qekp/4DY3OJiyl
idRVTx7btcMuqriv+mn8jJ2Do45wQWK9yYdL6j62u8pFMx15I3sU0aG/rTOv1YCi
BLcMIqTr+/nBHtawSIewnAzi2rii1c12AZJZ/aPneEm8+Jb/vUic3t1P/3PweKlP
lpp6ejms4CrMnGsNP15Xa37Uy5TsUPZPB2k3tpzakrBg4GiiAJpqmCuGiSvVUv06
yvFTNS3qhf/gWoJWVhKMsT9YpMCGafCZim/HsMTln529z480zg2pz5906/s97g+C
mg4lgo776QpeCu7Dke2c4gZPqWt/EGdq6i5R/tF6pidBkDyQ584Q8hSZJwe+F6iC
TW2DTvwJ9zGMcefb+hILfFiI31ioj7O6LNnTp1GcovcxkWQVi73Q00pVhkciCDnA
HnCFew66JZmkdx9SBeKL+y8rZLKP5ICmCnrg8hxkjO94FI8u+1nNdNBdCtiJ48ua
avpaZ2EtKRz36TGPbOpTLi2oHn0qM8KblR0uMN33tx1KUTqsc6GLVZ1yNuTA9Wsq
SrlVkEtudiIDwwjQoalBKZISm8i9S4QJP/HIQiwbS4+St4iVpx5EpVy21oIJoWW3
ijmFv73p/q0IMGgbCvwTs/xg/Dpaef7WYoO3k7AcZIF6mHHwnKsyMglK3KsCvsXj
kmmwRkwTH12++PcktwCYW84vlUKwxFaAD/2oZIaB4HMV05A+87ApmfZFx4sHYqhl
C4Fro9R/waLeOG32/zj6TGNd7u0Sb0FJ4wgSTwHTwolDOLI4RD0eYDKKk2MVTnjI
vheysTqTYfxcIyXmFkRW3fFGCTDhft0vEs3i7b58PIn8dg7lVcINYBtMAxaehr1a
ReWQliMrNOG4RjPB3kv7ssnCYSFVM0NWF8MLSs6vYeyVaLVL084D7modAJwVVU2w
DFYn6wqR/GCdXl6ejiMSoWrUNh1XgHduN+971lO/xJy3ofCN8y6BPngX625Hmhak
vp2f/1897Gj7xNBYbg1Xk7+KhX4UDLMpeJQ0FEL44T+YBeR8fOg1JmuOVPmDgstG
4arVZrX1AYVtXMyt8qbg0XyOYJP8yKjwxQVNUG9NHWvFRQchAjr23IHFcH+2tDPq
mcD7IC7vyrqy8Wxjb78wvJz53TA/NCLKHaVhXuspoV/Enedrpi057FyiwxWD/+b9
Bace+ucSmqhraXQbs2izUaMx86sh2fY+VDR1jQEXFAdiq/QN7qdD/hOT71XfLbJJ
2OK3oPlqDw19y9/brCikr6qjoU4Hf491PKimrqThHenPWlUuFfWsz5ulr78XJZoB
bK1MMbIoPXoFlYXHvUGOwEdpwm/f7iglK0/+cmxXT5LcpGa+7ZQEqrBMRJO342kd
34VY0vqzlX7Ccn9A7FroJpvZ1+kMG0x7WAjWer/bUYnaQupILbR9V5dPaVKvKPuj
0iyS3v/FrjGW/SCDoJ9ym27dBEl4B94599t6lSEu7UOIcshMg8R2BlskCntWB5gb
Lg1Bo/e0Sk8/JOLOcDTAgs96L8ZYlQJSyESFvTH/+xdxpYmGXkwvN7vq3/+aMD19
FW+F7mnuFe8K3AtIeUcEEhTaDzGsX2ij4o2o8lm2nbYXbP8SwDmNcXHl6eElGxKo
zlRD3dglwVIREMk9LNkxwTE/w9+PTFvMmjU2QpXDGtMWPBJH0vkRRW8cnr8k8Cz6
oU2dI3Imu2SMV1kvDieXP/wzflgMIYo1J9DFRqYxqhggZcogtBrSXDYkvJKZvVBy
PHfsnSU6XycjD8g/JoWUNfyFklGNrurXXUIw+KldRjfALcGXkdexiCuwXLNOTi4/
yFB9qt4f53lJs809BJ3Xlr80Wk4MY7nQhhVWanCyZumRbw+2ocFBrqEMhTSKPVDy
4BAn2QllgBThNHzJEW2fQCzUEitp6OSoRwv8qXQKNXRrgkvy+JPO18+Rm4RxBREW
b791UcZ0IeV7H8gz/qoO7Y90EAvyPdmI6fbG+87T59dSPwmCSGLqbPJ02Tq0pjLj
W4u/kJS09oHa87G/AtwDwmqpKhsOqz6Xzyd+ulWkgrsPi+B9fgEfY3DKeXCG4q4j
JTTm5sl8l3wIPH0gU1NTfv8vZ2QXeccKm6/nAv8q0wxWr6stS2H8WhLa56ShyYiN
a20BR9uYC7khfDGMu/R356auj/USiLqedzbCAX5jpJNQnQQncvXPTn+nc4hiFE+n
7CJcSGZkJfFjQoBr7rOKxQ/vz5d+Ex5Qit6wWuGUrxz1w0oCLkM37Eo2v6F4l0ya
ceedWCVjyaqPp2Rd0oxq/xu3qGwa3hy/Gad66+FYHG77noNReFl9PmMsNTT/K2v6
fafcW2WKMOAKJlhoBennKScFDfYC5bXzNrvOKblLwWLuDLUGYMx8/gdhSjs9+U5D
n0Ih5p/G99syO3+nOCmwhAY/gZuET0DTW06xEKW7frNTqJ9MrfG3C8UI0AWCH9Hu
eQ8Pm83t4O9JK3js+3/YashS82mDiA4nuXL38Cr66ZuOJy6PXDrxxXcoo7HtAqe5
bJXmILAdTjzsshZFQJrP7k0KE+i5K3cT2M2ffsBUNwmod9dUO9GfjnGCWmcRbSlZ
HiL0DpUmGtvzFFbzVCKltbs1YsyP2Er5Oh3fv4KCbJ/Z6xZnVABKaNqcl03MfbR7
27MVjWcZ1LAEqLfK9tw1rqR5jnMpm0lRa5jCIFgzWBcUF65p1v16sx/oXrUGbY4q
+xpOxZ81NORTRWastwYP+5IxIhVLlAU7GETqC/ieiz1gur6eMpOaNA6FYEiIHlMC
UOvCw9F+ZpAtoa2G2+nJJkF8aLOcMgwkuTtz2iBMqLSqVmJmX+aiRK76CwPdr3BD
R+T/jnOXPzCT/ohQEPoH3NK8tEoz2mwpmA3YiyKvoK3sxTaRPKsxMTzIriDxdhdv
MOV/rwyVjPrk7OiSigidp8H6x6tJgZh8JFl922cmWtTLniVQIDMstwatbhPABfyv
zb0Gw6dl7hPuxDJLFcvuAXrrIals4XhcHhJt7PYImueNPigOANB0WW1Wzzke2K+S
1UU0ftOdBD8zTdDr0ugcVS+HrKKbhjvz5PXalXRyzJvVKO6p72vaTfJaLRzc7iqt
2oxe+tiAjcQnJYoKuMjQHtk427HQV098v7OIbjwkZ1L8RACP0nJsYRQAzLG9bCB3
67WZaCRmea4aj8LYwYbgZPulLXLhZId6c0scfrbY48hVkrTt+CY5P5HtZNlJnEqb
7JmNv5cv8b4DEWql53oiIH/8CohQcv+hdhxDgVvz1vFqogq0nFruMjXbp+fqs8W3
QlocGxPqZY3LeqA2UEItoXyPxaAAM6209nI3V09nEIiihc9QVgg7qQCuU0VY42EX
q5/8t9XiUrX5u70S1fjs6ACvQPcXgp8CdH5qABiUasqU4M1bXq3OU9UNCjuVMRGM
4Eo7yLmjTWzIitlMJL42eqDQat0oaUkq6rl6pvWWeTW4r7ybcviedt9IgoQ/H4rx
Y4KLz9o5oZ1V7hGv+4JYRlnTATaSisZHRTEHbsctrdeuq1eR7NelLWunrKLc6coX
FOTI5oLtqnTUpb4pnWkSQEeG/9ArJPZ4XK5S72PzSLC/FmRJKuE2pgB0l9pFElzv
qpsg/hvikJ3FUJH1dzJgU22WFilDk6qQzsRhXXCw3/o7W9c/cEVAro0ALrYaNo0W
ZzHMDmIOs6dFEKhEElE5Nf+DZj7O46d3TQVZUcpOpp53+niV+wO7lxVxFVNad0RA
KuQ0GAoPr67qnSUUQj3Uh1id24Ccw+PTSMg5vER9unqUdbzPI5HJC28lGY1lUyHP
Dxu8+1BYM0555VoCqQTtVHFl2+mNnZOr4uetduLv8sTqQf+UpO5Nqvi/DLnBhaWk
hRNsnoTTSH87npLE641Qegodb3OS0CXW0k8NKYxkeooo3yZgPqM83DgtE4h1WIE5
lzgA2LqyD0LiOL+UE+5q+lTgXfJZ1fF/Eh3DuXyXTIyvFahMfRjymu5E/IELWP2v
XQYYn9qJ+k4lwuU5NKkTN9UNVgESOgCopWmyUzEIVFvm+HY7j8NQhQv7zZn1EBMi
KndljPuZgeq4wrNvchHQQdrjQFtI+W79O2Z/EzkCjY0Rv+VePyq6CzZ02J2DMDw+
KTdsKj8wLicTTqb55uPuTc2ex1CNGjR4KWxQ+vNZwl3n3Ap8/OtSgXCi4oOI8dr4
8gqCsWAeI2sjfUmKzfS6b1k+eNVeqpGXjKr/S58sSeX1yJi0sIXlWUnJrQDCpQY9
vjM9QMxTX+wPppv856WVGlU2j2B3efToY2bEvUYQsHw7MNUdxZGz9EgV7tcQhK05
tqRTWU50+twP55P+MAj9oGXY3LkWfWXgKWLFHJWk3IY+7fZArZX2IsCkB2W3iJJz
eGmJJFW0Cp63WgNR6RBflIPGnLpaFba4gkf526RWzO6nv3szE8pUfjjhU5ksml+g
Snm8t45CLU6IsE0km20zrZ908RNrrIixN+teJANCtQ+Fo32AVeY6oTEsVMp4U1kQ
/yRa/Lk5bUtQBcDyIwioSMuVyk+NUEYqSDDceCCl1RlN9YvfUJU9fM8Ls0JT0qSW
epFN0g86SZ7hqS/H3EFEvBh+66NAA5lahCtl8DbfhtJ2eK8/Fd/HKH7FlK2nB2q7
9J1K33q3q9YdXrNOvwEodYL6LA9Em9qfpZ6Ia02DMZW6TUG9+GwDPrS68yhi9LAT
o9oInXLwl4UeOGLluxhz8jBOK6/pDWlDn0etNSbHi+55zohwSZ6ctxumQCK7imjT
SuTyXY2WMFSBMNIGHVtfpmV0GG5T+hESLELN5hF5MKH/ZeFmNfjS9LoZHMJCZjDT
tInhk+48Qw9O2GDam8S0fkw1DqAa02BLRi+ZJH0CxMPzlDkg7zzLq3iDcZEI74ka
jhLCQMnBobtUdGnvNjoLakBeRxxwC4HjmWfdN6hhqpiA6ekNKBH+sow1buPf8NZK
JjkLcazHFMD0+6aL9yqvy3FF69/gAaFTDQBGvak/NwzdBVOEDn3x27SLtZw+XWbY
wHDF4rC96HQvHborgkDR7F+vzqSzxX+fgP1htJ+XNq3rFguzWJJyXuVCvbxbMpIf
cHSHaOXTSZOiZSQvA7FpGVyNx/5znO8nr73cYFtOoLMMO95rt6tkb1SX3c4U6NCA
EupwMF4EncPY9Rc4vGNoeV30Z9R59U9k+cnu1Fp7K/Wlz1K0uDNNNhlxUbTJ8hPg
U/SuUswOKwodOSkScttGkUvfPuNoQMmLQWuu+tzRP/ofnrFd6UdAKLg0h+gRLeP0
h+Ouv10U90V6AuTaCC6/JIj0gWKQyFH73qqa77yHXvkkKarQOuJREbKLOtdPl5KN
Jae2Dz3NMMC9nv+K1Cjj0uWy+D/HCowKsdX/VW6PwF8OS2Q2OUFyQsvOE9RISR8t
G6yOSmfsJLt0B77BodjjhJ7jhLPsZRFdF3+0JNPsgbZLCg0hSH9XwDBVqioFWz0S
ZsX905SOrFqmRF/izE8CtWAa0T+Rj/E+IRTjbQJbuMwldw9tD8tZ+aqqR9vcbyc3
aKJgrUt8e180AssEF0Lfcn7ciFaRo30Grb+9ATXWn/A1/Lfqy0ybBFOTvaR+DrFh
jHzK71b+jCrbkwxOc22XJCHv9dVbiKnvNBkeoWzuCFNomSYbMIPxTvVw4zvswRWf
/KXT70utYeepOnb3ot2vCi3RiQVTs+wExyMDWV62eSa/RUfKL91tzXIFJW8RF95F
D6ViUF79m3SEbgG23AGgIdbNtpUmkq4Xfpwems/0j4wozZdphjNFSOtikl9YgIUm
NoyX0oP8XlN9JPZeXZAkysCwprHtsN+1b839fSWDyDdxZtgjO9Og6H6z9svMzZIq
0URdTxPO5aQq2PNEjp8dZtaF9bGLbIPJtrHBwBefNrb8kgcLJ8KWPTiN1DIp4bO3
29o+17LmAigx9bLIsufwiI4rKC5y0oJS//oyfMEW0kDsnm0U7+fACseoXdJeOL1b
BbpyGjmQE2/t0E6g5KAoecwpQnk7Nrvgp5eY+z8xbOdTXZ2gVIa34bSWzq9gFf4A
m58dhv6csekIcCGF0DyRs/lEFTMWpTiuIvsZDWoPP/owbkvloW14YeFlQF+/JMtO
L9sBIkFXr7UXYcuu4RpmDi8gS+XwyR4yKPaZ1ZmQrsuxhtv+NuWL2p0XCAE1DH/Z
dEXr5pSiUWpC7n5D2MfSY9ZOTn6dRegSQFxZfzZeEnbjRipV1pcHeHsUAayq8wwp
WNkiTXxVRMuC/7jxJjfSL8tP/HImjmO1WuxCpRmYQeXaPuG4tOl+CiC967foj/6z
eDiKmxzYSec2OMtT4rJd1zDu9CKfxgylr09zU+TyKdoPraUNTNwTcq4Iq+4Ni1lw
iOM88ADs9iexns6EfAJxcMGud9GIiT/TTUv6JCclddDQ0jzjJmoi7dglnufHCI7i
rk64UIpRL4+nau6lIFzECMlSJZjioPs2NpVKUNth7MyjFwTRXsG05QdeF/ZvZp4N
1vM5LJXCEdSQvYRratyMcY7W3ZgVMyYokeu8dDx4jtjlPfXAib1iIYAq01rnZX/t
Wb428R4LepzlGj5rM6U2dV18x8gg9pPyfUK5Rorqjc5Obpun1GrTESkbvrUE/rIp
74oGc319HHhm/Z3AAYunhljlKACo2axoHBPb27zLnypbOhUdy0zAci6qyMYbuO9f
e0VktVHZj0XiRl6g8acgRFdb3yJYoC+pYBC+6KZTBq/43C0tN1iNA55qhFd47/Xz
CWHFy7LoSF7eJzHpBUR4+gC8CE+0ERZxdMYxCYhz3p+2uGjxt6qKZ4tvgmsQjZM/
RANOtEMmHhxr7HXftcLZZHogF+XxOPN3SssVhRD7KpZUlStFKFk99c8JzxUj7Vvv
ImulnMG+nWHGLFLHEsN5lneNssHD2Un6SsBd6XwqIPtu/iZwaB3E0bR+RuxfW55U
8Kw2t6UfY4qFXYKNRsUCj19uu0AjAxGB7VjA0scNktPMmauULx3YsZ+siP5QH18O
O+OByiBWaw2IArGDKZ0dNWum2M1dr856c0Wz5oIdv8MMFVUAVk0p2977WKCWaMQA
qRG2ikZnm0OlVEJnePQ78hYo12YUzTt8OucnoucadE2Rp92GftlXIqKzy+2it6Pv
o3ybcAuPa87rsXHhlgI2iIrLGxjoCo+wdJYl4InhDIt+cozP2OH7jNSnS/PJtzwX
8VADRR3n0BD0ccO5XPkf1ZIiWYVeCVhW3yt2F4GttKM04JMOKgcwrXn6T8pzvhYB
7hWp5y5R8xap8uFGE2feZ2bEUsbqR+eWbl3wIBSAyqyG8AHRsBj+X7HmI98m2q0n
L2DA3+luZiamffUInEbufEfKey8aZVOsm2GGmpGZo53wUy1tRSSYEiZb4XtOphjy
iTOjGkIOb4bXd/7LUeHnOdfVFprh0EdQ/iGpV4EXjfz279I7t2CIXAvqgbxY//S1
WZTXloVkmQAamcc74evq+x1Y7z1vBBUqrwS204KRy057/ZVqarmnlpQYTPjler0q
Fn3xBpk6QBX07X8jmLN/S3MpISLocWCdx2kDnMbrQzgCWSr+lAHxHioU8YlVUzdg
uTL54TkRj7DTVHktDsea9NxfiLfAGN91oLOED5/o0M7Db3p6bEEXBLvC8MdsJbA1
eDWYo2AzTFYxL4lpMmPWkJ6Lmuy6xDEAPr2KgLA/lVFa0+wNbt2nRxiukZjvJP7n
4mmCqcbpgoWz7St4KfQDpkHmosTjJd0MFhQ0/+ZlDA0Oiun+Bs27SuWeZ6RAcSlX
ghu652EkRUq7ZT6+Hb1bNu8P69qS34nglqU02EZq9NuSk+q2nbF+K0sVb4AZ/UGY
bQWoAYlIL+qcSxmhZVkYqp+iJdR4HfEMiu/02+Kd3oQwV4HvF9uPqFSkq9XcMQ5S
rkqsg7D5vJyf+lgN8tkPKynbQQL9K9pljez9gixhGCf2MTuAptDB0YK9ePlDaL+s
V1Tq9I/Kl3jlw1phPqpqCXnDBuAALOQsJztkqu5ZhoLOOKiQieMDZEkyzlpMUCo5
1o/j6VCiO8nEG9cAO8YeEZ+yywLzxBabuc1fJS4bNj8ACQ0ydAj7nLz96IL9FXfJ
bIdgkCkxjRgwVXY0erAOeTbFIhaoP0SdCOTaCNdIogywD5hTR3omlGtFN6kXe1T/
2QqgDik6XVY+iSII3Ot7IW1xgYWKouiZ60332ln02c+B/mFkZFokFNtviLoG2nPh
2F/uJYfNJkV/X1UobDaItjND0u9F3hvrulKb8wzYvcmgW0FaZcmz/ILY9SzIkfP2
5X8AlnDorvpjfKKJyhNC+I5QnFlVe0+TILH7WYAfMei5S69WWqnE4LJfw0nv2KRo
7GVO34mtNyWw2/ll6pd+1kXWpAMeCkl6vQ68ZlrQEJs9/kgbgMeemyBX4NiNZ6d9
K70niZCxzfnP7QRNVz9f7CNDwQXFTKSTfq+slPGRGlamgk56c3wdkc4+zXUEDKYH
5DdaTmWYIEX1wPf2OAYQL9gSkxJ+NpPuLaf4WZT6ITOI+llY9VduAriOs9prJJsJ
tg4lU4485djXf++B8d7MY/kwPJA3dC7WSf7VmwHZMooSK+CSQAj+8OhS0lqL/16z
Zgs0rwnr6if/plMMZLcpMsLjHnzTkCQkRP2CbLZ2fy7h3qFCHKoOEXp86kZuYEMH
APpEjyPV31+qhTyIDhMwVDqNzS9RwCD1WBe7pOmLXSmzNTNE/7RXwEUHpGYDDc/M
5cytgHTWLStUNews0r96/bgVM24OA30itmdVVy2NwhcPNGxHzG4Hv7qaHbQuxNuh
6aZAJv64hKaIB1KommYu0153EtvrfSPye92lMAxMizIWIZuSHQRo8BppzBGXWknT
RSPxOBbXWotaL4W8zaVpL9NFvjCXsCjcTGIuYh26zJUjW8Vmvn21sLYridcG3+Vo
g8H+3tS0Auh4xGdk+YN3xc+q9FN0bZOg+QmONIDfin/LCF0DNYcoKldcRACpJ94e
0VcjM0DiMZBVBX+zlFrpJm8YJ45RjBgTRiFVaHsj7MA9e8IJFhWKuPA6pZibg1jd
BlVsq7YHWN+LLiXl6sqLV1IStzZ0i68UTKt8t5ksGouNL6huVagmxDAqDmeyXFlE
PgyefkJTw7AilHSpucLHrGiwpToNy8s5ZVttndT5Sbvt+F082z64JxT4VTS6IROF
lOG7A2ZF0hsg60QaYdKK9RkCmwfGLXal4+3LqlWIEJyMMp3rNdAtID0vx1maDUgd
d8lCevi6jvSvDz83BZyBe+ZeNVAGYs88FGrntudCK0lvJv5BlDCIysRr6Xg4NGMd
fG6k1RYI2EqwCQSRphIX3ZjiGEdNvrkUa97+/eAh08/YIUDwAczEdrlQMXRQR81B
SUBWlaW57L02R9UTZAuZ3QSXeMrApOVjz10mtc/MiyMTgmMNzEIpzGIbUgd2nZWj
7HU15LzvzXXKI9nKaKyGZw0yLjFwML0p0KDRlea3iciblEhCR1n3si2Y4CA+pHbY
GGL4PreItk+FC9NGdTV+nKxk7YJBXFy2GW/l9xxZdufKL6p6mW01piJM/bxGoi6h
yhuSJrA3Jduo1YFGClcqXY5VtEgVRiFinEqOa+rJd/8eDZhazq/vWnoPV/u24gE7
trhXRurQIL6o9jFaE5su5yD4ukMbYotjUawOvpztq3KK3ysMHCH+RjeMBTwLOhLM
CTpCO1Yjlh538IgDkS+41w9qwO+/Ug0V0z+E5/g/Oea41FJ5SCuQKZBJJ45DRj1y
9ULjRlWBc3s/ymcr/4OXbl1zQ96cjZT7fAz8Cq8bNltYp4j8klbcU5cqD9qvxjGm
8J/j6F8jRdcVk0Y3NonGf6qfM05d/lHFCiQWg7p4jPo/ka/BegzvXUQJxws+O3/6
wQJlFdOm2rJFEexBIF4Vk+KVtGMX9imrS4mpSsbS0ffN5E7jUrnWFQWZ1nAasAME
lw16KtS4OxzCJnzhg2mg2uBZdr0WBRa85DxhPjb7ak5s8GzhXUHjWvnj/I61z3cD
6I6rBMwENW894ZSj9IuZTJ54hjUCs9MK3Fh5ULWw7ps7HvQTciH86JubZGLFpeTd
XMka4aIAAhhdkz0IaP4PbDWRPbxKwHzpsgL/S5+60SL6o/b9flITJevM23KLzSr3
obaijr0WnBwAqyMnVmE2Xwm+chgXw76819hOcPLJHhfSQy+4FgFuA3pCD9CG3JLy
1MMtqUZl4nbNJG7JOmix1wk1JqGYM1AC1AjVT85cf1hKAMYex6mUjvj+P4Psmmdb
nvrCSBkdVR8dl1su/zQ6WEOUAcvxtwXHNhgdX8CV0eY7ZmoVRN83v2edPaOE82OL
luPpS/tLp7INGLAViXnxwYGS2XyCnUMgod2y0zXJTRhsE2C3C4t2n9XhNTcBFOBg
47SCIDrtqnxOLfW/pUb0CHDHiLoF0JVZOI0+YFUYG7v7IIXifb3mxpX1rHv2IlaR
duXQxk7Zm+Uy+ba/+19lrSUaSHksTV/JqywA+0kZWZ31z2AQu2jgA8LTKTCuovhf
nCGSiFwnmGCfy5CGPbv7CtHeJkUIkiSoRwgR4YNvY2Wh8QllNXkF39Pp4lr49qkm
dhrPdICMy+Ds1x1q1tZ9s9uMsCVkkMsN//2nMPf2GQcC5WCcbk2hOHcFQWBluaIc
RsfS4vbukDjUcCzYW3RcZR91ny92NIxt77PGK+rdSNUHMuNgrXrJQUI8FPUHtK6Y
ZJfl0+S7hWudZdBpFz2FqxLBhOI/3liCIVyj0/TTkTSaKw5kXtMEXM56v2VLfxLZ
P7rCpIdAxyZYTlsrTRRCdslHhvb4/ZrhVI1CBUHPLHcR0uIrsUTqyvrUkMH864wX
s72O1loZq5VkOtxKG34Tr1acsIjZ1/Ok49NIrpAPCZD0z3BbQPlObiRuPNGbVcei
GF0+ktoWbRKjkxN5EguaO37nUEOHCqHGfqUlpZs3zZr4v0/Qukceva9263yBsNlD
GQiG36IAT4fmBNfGCzKxTQ04C9ftM8PNCiZl/Bdc/SXxQ6ighWWSyb6q3r3nNpKg
zQfc5ZzAOljvM70sNvZlCc186FOOadt0BYQfSadVgV5GrBxfbVsdS7HzpHBQRewM
FDc3EW4wxeE5MrqkNk7h1MjpDip33ec6c6Qs4cdPr/xhmUx9xDh5mXr3JF9ahXfH
d2VmtVIvi8Jc1F5fr6aTs/9UFMiausyqTedeoGfTGFy43FG/qYtkdFoa+MhDT95V
fu3XHfyPuC5IeWOEdgm9j4u8LgZR6IvAwj0SO++zJULm0zMLF/cWI6rfDBztxjb7
X5ihobiOxZgINh2SQ1q6T6byy7HQSn0hdXHgx3yt72YY3wQEicBMA1UCi2saW2DU
Qc3iAQLU/KdQVYVAQTGtK6P5bK034UaBUzV+naK1SO62P3JpzuczHHktG92LB24E
5hoh5m4i4WDDVijT5DQwwvSd3ooDz1+AuamKfhsw0vzojQ0vZTvWe965uuGUQyfA
JpQUvX19lI1/bBeNPxdveV8BbbH4d9suuZI+v31ptw5yiod0yWFzGKzcklCyXk9A
l+MMx7mBMwxzM0bves1NXVkG+GYgzCzNW/1CmGwTdp0CAEDavV2VOvAJBK7NbDCH
Y53uYwyI7mbNwgVilz/ceV+tYTvDIb/xTeQhzzO6o0yemeZWQK2f92T17rbBB67Y
RT612/5nUrxtG7TZDvsjPuTn4CkcFY9gHgIF648XKFEH9vaAAa456Ua7D9rH4mVk
AqLJ3iDb3Kjil8oqaQxdwvW3n7U3Bsjk+gJJOVuFBeX0iVbNkHcYGQtO6t7pYU2q
8H+bEOtj7JlXp3FUWsV2NusjttQZKFE61hzlcr4JwegL8DWEnmeuSNh9qInsL9M7
nLEeSZWOsgOmpUlPMZW0RuIFz8vmv55NFr4VvS8oPNac6iqFmpyzlNK7mwqz/Kmd
h3p+JLUKhCRflflgPIjUjwug3HBFerp/dFRZocm+ZA7Oh5zwFvOdIQpJYdGz6H1a
Pw9nAP/Nc+lW4hXMCPx8gkEL7vH89WadzwQPLz+fO/iKgEn6yhtJE5JBUAKyqdr3
Tg6J3/qXSs5mZGB2zOppW49M6iPo0aCROLf+HkzCXAghzsdEWAFbaWy2mZDArDac
MIU0fRvP1JHKH5zLrY8fJIhFoTTMzdirEpTszt55WKoDLsxXxEvjjEopPmgvLIe+
ckxGPd8zzMqwS3SH/+4sjol0sPydIW9Vd8e1bCRPcX//Sui8W19P/hwoA8EZMIEB
WOYsrklYRQYxbFFUMCdEg/fOm6oI1ryhEaTgYOJU1bcutgJmPY6My/gCA2H0KSo/
T5XRUtqldxxEDt+4dk4AAvvmGV1n+C65sXWSn5XQt9JvQD0oe+mvOavnyggyazDd
u2ZdnrwzpBf8Nb98UwbWLVzhAyZMo4DQCAPZ9sXGEs2VW5ijbMWqXQYq5DFvW3IB
MSshM2RDc1di/LU85qwGBN2/24LCwtFVs3gY83N62RhAmW4Hn0yumtkslQF7cLKL
/g6EE1xx0MdRgAVdKxd3w4selFHCI5VKtd88L5WKhePyu1+eUOJ+4Vk4dsaIRmJL
hDZz2nHh4Hvnq8sIQTDazF8ifAEVbNZqyoKeA8KqJGe5neOx4wCjV4WufsjuKlop
oG7OJhaMY9MzyzGafbZSKKzQWOjrc7HB+RR67goYL8/RkFVBpj9BdceZuXrMxNBY
4gqiZugPuFUeVM/id8WOQGzCZtVDnkQkm6cFtYiIseGzCJv+/u36EgJLRyMOeXgH
TxCPSIivrkUj+6RC8iQvG4bgLdUmA9hxRBTQxGonbIn4IHIml+O0H76NIr0y1cTj
vK96CpAgK5WEstlcP7sSjEZ4Gwyxl2OCGJa9qkIiR21H5tBop2cc7M8aTerYpjJb
i8zKJ3Xce4v/HjTET3VrhhTDkRkKFj4dYX087a2/EQF7k7tUe8azEdEqq6Pn4zhb
9LqQLx8Np0xgVU6R5Plo7MCcabMzZmja8RQZLst8RYAZLhmS2h4KZyEvrkmcLSC3
fY9TDi6F/PnV68+qLhPCrBAmfOyNXko4bFF6W/mGuxKGDi8RG/DH2TrL0Y1fMY6Z
kPQc2sCX2CFv+BtIzAQd61ZY8KmERPFkNflZU19vWFGbE4ulaMQ/DNLwQTN+W24w
O6W3kPkH1UwZhfezgJDVt2kH1oBMWLRs1EFIL9an13Oc/KGYzVL3C+Ghif/8d7Ac
DcB7fCNBpuaDAnFd6vqd7vS+rOL+t/ZBT3kyvFUlR8XToKoC9wbxF/qfmm1ztgA9
Dinf4Aor2z+eH/lcGWY3kIdkAiZHigGc4IhrQms9KHpSpRTxxD2FRgY7iUuNCwbg
DgdhPOuteycscb1AAvP1rdcxU+yV0mHE9SnKXfKcjGTbTIHN9pbNt5l8nunI3nCL
HHRlV8kmHnAuVK/wDd3a6hmrd7Bn6FEMUMXIftK1PFn2Sk7XcjEdn6P53Inr6QMe
HlCia7AI2GdTQ2RwYMkgCCH2wLx0vmxQI2bIm/jgH+i9Cjt56OdxgTMvNGhet7vS
/DY3CskT7r/X0KgzzN3UMlzWwQXoYvCB4r19onEz15wYwzz8cRLY8y44TY4xTZuc
jJBCoaNKTNP6gWEChx5we/I/L+604B5fX2VAl/KaKg0LRV1QqTqotV2Oj6y62n4f
G4pxhPtpOGevSdq9QAAWWHQ+QyFO00dIxAA0mvMuEpko1ldovAGJJ5wbUJgrHcqr
4CbwX+Gb5BLX6LzMw9370eH3rdJa03zBJVTNsoGGB2aLOyxiqx8oCid/T2Fo/8MR
s0QBW3VY4HOqAWnc7tHvG0dGxV9Sq52JwEti9615xNZxfiaOtjEHkMTzatpg7wg4
kh7vDm4k/ZqQd+Qr0CfQz8R5A5oSSoJ467EMyyrKG1leI3qegjfXeKGYUhl3FDZe
MxM3syv3HHkQSs5mhHUvERUzMO2ywhabf977Cuo0uN8f0kp2wGy1ZjMh7DOqMJFW
U4FIEmWBqZaVQVbZObCYcyXESD3dJUmrQt/L4sLKlGBDgYgA7VksNhx10MQB/GSG
2BEUjyyTEVup75nHzO+hEoMrzA9eprPJq0oYXmvzSibI97p4WJ/zxoT5fJYtJUP9
KgDMUq0Boz0IkNCSN0Q21VBOOQf3OdXgVzvyljABOl7l/f/l/UGhj95vOOT0acAW
O/DLcmXEfVt2Fg6sKdQ/7cny0EvVaip/EdI1a1PrxkfHxdw0I1/hwWoZdLVOpaaJ
jpIEtAb+x3qN+TTKsAA8zh5Lbs6KrpQT6oEW9hBmFrCFZ1hDS/t42cw2jA4r5jjn
K9mx+AIUJUDonbkITIeGs2fcNw7Af3/ABLLsWZflLBTDDr9VdVt0BmHQDryBJ5qT
uSQP4lkqNKlIqdBOsp0fTVFLDXvw2hzLm3G+IcxvntSHh72rtmCpaxu8P3pEr2ut
nBkHIgWk7mVJsN8y0i6TgXs9KTv7MOaevg39w4uGwu3RPDp7zcmXf1DiydDfNcNt
a/9t11wvmuibNiIP+Zz8jnSdMlhobJjZz9IVm+OYL3NTsyigCN/n2mgFcZh58Kxs
0iNrECSv7OONCASKERsn4j8vqwJNWvAUum0F1NCguJe3orlaiCc3pW2grIaAjf9F
4MtIbg5gUdTTkTcM1B4APJLG3kCbrFlHETPb/a0AjLKBfthxtv8R2pTjve7F7i8P
qWMiLHxUnnVtEHuDMqkp7tdujo2pzq+YwV9CtVpagKxxsLmP/LL3376bI6QrAqDG
HeXCGdacvAXMkOBJYH6O6kCtBKhvGhfUOIweLbtKrU6q6Y5MrZe962bzgwB0i7K9
jbss8BA87AhcCph/K6Fix4O2WuevnThaVMiueHIPW5mgTLx6rPKI1l8l53WMm3li
p8KCDS6Rjeua5+KtwU1Wf3d5/WR9GPt+6Y2eOPbpKqX6/GxwxZG9G49/uVe7UPM1
PmSeg5sOWboGkZvRhg4T3h9YMTqiDquaDs70xzbbDnhBGQt/0oSGL6661bF3HgFt
5NHKWMEwbom9QF94nMfA4MjTUMT71ge97LwVla8I/5crz46JA1+dqCdoW89923V9
foUNrwJdOAfMTn+RvSDo9AWfTv/vw4VZz+paM5r3C7gAe51mIB0BL5ywwKzXp8eM
i0j6XkAzerpGwnFM3opyXrT1mRKjDU/SDy9486ascajIcq/u+/LniNZ1uOl+A71h
Fl4fgXexpn6+GBxWqbxBH1pciIzVjAj6EdE/sIVtCQsJlSg6dgNQ8PhWG+I1/+oN
Wk8oG63N7uZIAtGjOdYlqO5jOANxWHZ5kSLcq4B4kXGlR8XTiipa5qgdM92iCSqW
w5Ii7W5fC31StPbMonjuKIPZUwbTcY7/xmVr7IABnrk/1P3fBhCrVktvrXWWtxhd
LdtefDmp8rutbYhIdfwkOV2SF3Hfyl0228foMKyPC5AbVd/YnaKraVdTAdPlB9Mu
nvLaKJf434fXBYchGxYIfrGM+/3sfD4F6FpTLTkKHC5x6i7Scg4ZQ8/An2eSKIiK
iEI31QnU/jSol/TSJkNNNqibdWHVi3ItkMei4jYPrNEL40ic/MGks7Ye3OM38CKW
3V2BK0ivjI8sK/l6ZGdwiACmysbQKYXrxFvH7+HPKbpSB3T73D0Xajva9jvbyJ2X
4WJlVX1oecj1lT1xeYstDAYEVKzQ+3lYfHUEsB/ffMolNEEuk0Q8VqHL1j9wEqEL
uq3hrqNO0atrLtryEYdzEALKqnhKy4Govrufl0Wl7Wziryb4HDWoGX7mhrEwXkRL
MWmTpsk9ktkzVAEhWbtGQ2jx60hxNOCtCES3zL5VOSa9rwN4p0u0+nOBQFJ1veMC
dTZ9RZY5NRihugKdAxW9UX1UOlOomu8hOSPZvgAJKhBGSi4wssyusCqm1qIyPCpq
mCJj1h5/2xJ14HCyP9a04RkQIRuGjLT/kkpG/Qc1BSbwvJ6PMJBMxbOR2NKD+yiv
A0F4piUQGnVWZ3t4u7A5RUf7lY7PIN3fjqrkcS6nCyGNzPUg2Jajgk3cUR9Muj3r
Gp5dFG8iIkthfGr6rIZGtqarkjs1JDHUHYPwNeM1NhoJZ2OwDL8rZjxf303wOaWE
0B/U2ci1nODEGiar6UuzrQWxCrFcuiLx3XUaXDkXJelXsWbILKepNH/oaF5bzIBL
YoN9ZEMFSKlF4Dq4tvKHyK6QBIjJOYt9VLklMxRroCFBdhRujbI7CPUqDjsjI+Ud
BDqNvg4Kx180/TFrXh3qVSZhfHOu+Sb4UjCJqJPGGgIHcnCutLeCJ3uAyQ4HD6Bc
+lAhz0obg82beozat00UanZCFAsDKmGADOX01qbqiX86ziW5yCpIHCwWmTMx//84
56Dw2oEU9K34S5aj47a80+bhsB47Mwrj7rVLaUe7AeY6TH9BRtmrKNzdIWz4r8+o
8yh2DgyPzw4VU09XZDlepYGDZYyFbaG/ekcce8B76VjiT7ZWSKY+sXiXLpwdxSYr
Bmo7GqONRXjnZDdXwhKXU1srJM2nTMuuevPdSZe2PZhWMfiRosxQCYMNkdxjODUX
LJUjWSl/R0HzKW5/ZFZteM4DOFvadox9aaIKN80nWaXu0V94gV3+wfeQbOrlzUKU
Z+r0z2YKqBIi6aH4nzAb/MtxqFAlHOZnBNk05r9FewP0ln4G9kJf7QYOuVJ32GRy
WtzA7G5INBg4/mHvQDhZf7RUTMtPEFG2+UZbBKHxnWe7N1JHaWh1wd/SgGZV5/cX
7Na0BTVD6hntRWyVoAYv83LgPkKpC1E0gwTyp4SInLFyGJducLqjTOeUKiRxTRWp
gPO1AJFHAw41EpTBfCobUYwIqLO3Lyh5wzl0bKzaT/3FcN0Jo61txiBwPOcYcuVd
k65LTeMC2fYn4eg5VmENscbG8wv5/3XsZa6pr4fyu7xVqiJ28vQU6XkgZfisRHEr
vFH4AnwbnVpNOO2AFtpOOSo5bfi1A0O50qS/E4E3zq3Jgx5vaKWP7t6RnD6fkvZk
OedKwG/dOfGKROd+A4eckLVpo3J33xlUVgLMwdBno4JmK9cLAU5Q6sXGNbBnDyXq
CYKYiN4mnbtU4fn18EEgjP2pBU3RgWZTCRJ8PPzSa/p0rIx3vaQrMMRLUJjfc2VQ
KI/peGJNvgUXBNTWC6QJi5iGjfkIxteLdRQXvYn9Uof6Euu0zezCLV4jgX+kpj0F
Gns9WhFEyIa7ZaEEVfv8RpDReITcwRXH9N6Bh62BG6rlYzsoScyoaK3uPYbJHk1b
E/N7e0UPqkWF/aGEMonhc+MENK+OW9gKeizlVIw2YJ0axE1bGpseeannPW+EoZjt
Q0SVzjbI97gcm3Q6r5tA/CdRn9s3PRGhQdc+CqFyR03CjuKtP+IZEEuB37pS1rbg
lRBKAYQLylv9xaVzJGpQVqGz4o5LRM1ANFM81NlAIYCLodsIXMfyaoEYKVn4TMBL
EEmOaUozq2quez99v9HOj+Ts6Tg4lTkCYe54BAV4T4TmahmotIBJfZ3SSJ3tGXMm
rmC8Rkkmhi7FmxD/jG2L+zsav6P8UNkbvqToA2YUWadbmZVXHoQzU56/gFgmlbuj
9FT8IdHGDOidIZBe/GKHPsw1pwTlcOAtXgnnI04gtYf7f0LFhPbpz9DXAdz+uPkc
YTXvRPznkx+EBBgwnRCM4JVIuRIiuGyFM/8v1kJPdprild9olvqENWVdZB49qMgL
WwNAtHg2ymL6dDBPsqVJj9/69I/xXaIjvemJhAsAryZEgJMiVMVf+ne8nCga0aQY
pv0Sd2drFczFBXP1e9LL7V1JZpgUZjz4ueCYXhgUM+w1z2yqYEhaJU7vv8Df8OmE
v60byrlpAUqrYlxGEocUlEH99Bx/CC4xig5DAb/exchCnNXkDcF+1y4QmaOCv/6k
EeIHf7NrEw7UWDFCCPXivc2IS5eu5XawcAZFfk92LzWTCWiB9lvqCD6a76uClrIq
N7glGgjEGbFiSYtHD5SWboQtJjqJp7i/8KJKytvRRwhQ4w8F1Zo8agneCu6Syq1z
S+1frNw6XTxqJMXdt5sYAeb6zDV6n5ib3/QHWlbb6exEYhnmpfKW3ZbPPEEGIPPp
fbVyDErbskSB50x+HhB03hOOm9OZtk8sgthSwxCKNWaTp/wcQ1wgWxIx9n+/ijV4
eHQkyL66ArNW4qx5Xke729/Enzx28yes+fum8jD/aRTlWnF9w6TrTiF+j5WmlUJH
bZ91W1GdvWNjFuhO2QlwMRtBrf61jdxfm0EKrMW/42ZbON2CnrMAQHzmMAUmz5V5
DeatR+m9xfnqNST9XvdLIu+nMBlOF7j6KOnhNK/SdnFsMeOvyeW0hXMdhnEte90F
qA5LSdItdFO2+6zMZad53aUAZ5N+MaqfnSpxjXssjWdDRqnvysCWeD3dkT2ZKkYs
UZV9yYqcANVoC7ISS1Rn95U4MH95/sqkiIPYg4QQpEIGhUp3dwa4rwPx2ppjsf8t
PVCJ9QXmKlJ7BeT6VygeFwxG89KkSNDsCMVyxFaPfP9NYLzDOyYDXt3zbfD0PLUf
/vSjfn8WML+YFtD1ZNFCxEEPsXgR+zIBq6yomdrPb4WvhpO/lesm+rPVi6EfsgkY
F/G4jksO+tBC+C69Fb580SdfcWR7Gkslc+czFtBJaLZ0O3kYvjYCtTW/sOeE9UpN
uNiw1HPRLnSS9u0hGM9wEAjanD+OZdbU3frKQ8+hN0BJXfCe/2nDTRG3TvUFdOtt
hhvW/n4ydLYnnstowmv2PAb2kMMcZ5fjCXAr+VNBFIqKH0ePqSI3LiJOKty1Tm1t
RrgOHVL9EiKFag8ebg9o91Q7Qz03ivLhpvBqK3Y3/Uzd/8igaj0rekL+iPj7LjEt
N1uuOZYTVTfVmxKtQw/blk3gc4FdW8cyAIBzJq4VegfQnKjMrxAuVd5TgowS5uWF
ON0xLd2R2Kd8iqTS7Z93RNkWB2Bjrk+oBARuEZStIvXm+uxXTn4uoleU63fRqsAi
TlmnYsSEDhjQsbqNYNuqCAF60qeFn6ZD7LrA+8CdkD/OOxIrdzLnPULplaKkFRSY
0UZ9IngoLlLPZMQ1X8pzSYrYB4NjeERkVuVJzAQTeNT8PBW2h6p0I6WnC/2q+DhO
ZdlAtmgkPaoRNhMQAiaxf54WpugFrh46knTnRCy35tg/UkkYc2TMtCXpooQziBT1
HqSRY/e91QznJHhoFqXjU8gp0HudwXQCotc5PYMbvbafH+DtxS+X5h3PKx+sXvkj
t9l3+nvZy+FWB9TnEik3hx2aAN0ecmV5VpeCDnai9OjTdEw+ctCklYPIJdGyAwUn
eGftfli2hugwC3xiR4ORERsDYzVu021CbgSwHhazbu3EAvR7vUeVPQ710ZVzkawP
bNIuEvVQn+TBgxVUfsqKeGXCoWTNK+LaTUxlMOfzxKT2+V4WObG7f5Td9oOxUe47
DoT0aWTMwgz42yihkEf8fQAoV/TuTz7OC2c5eP7ONiz+hp9vTDHi9Bu91XZbD6+h
K8cC7BIvSid+hJIZxUKixBtWnq8qaJJX/vrY9UEFljhXTHnWizhXPl5Eo9qtmUtv
vZrotcPl9/qIH1Ftkt12WZ3+piG7jK0aJuuNO46F+xoRv55HrC8OQZRjmk/oCQdI
wjLPBQfvkfaTGPaxsr49zBXbdbbwRch/86SY7NBnrDBHlLxROPdAha8gNWgmO5In
GnYwSrEdhOMee2vvqDwOWZajXmOc8BOE6Kw5fZi2hL56rWSBdK1uh7H6NskG8nEm
tIK0K/UXerqT/gMashJEpSlXrRlXIISSG6neZMLKWBe7hw9kB435nm+sUiQN7kXo
5kpei5jYwEb9M4KdeL3EciB+cmgEnu+gwhBPTPe0hmaTmaLe/omnwoGFeEZvbpN9
Tomy45Oa6WnQNd3e/sQFWHj8l4BTAozDUppPjq3eo4m0khBTV3Ohd6iqen+6uRrS
WnPZTH13BcD1mxXfjFv+YpZYsri3YpSYinQJAFSKC16a+cxaNWnO+XBFXYahYjA0
BsNZZg7mx/qfd1/Lg/yz/7iX1hQ6AFCiLQFLfDT/aeKBjj6N3TBq41ViM+kF5Ena
5DqrZjOxSOZboubht49U/2ed5ru1BTZtVncULEdZfGhPreunmBuMxsvpJxilM3yd
ji+cGvlIq0hAk0wWBxuT3EXy2PtNHsPL2DoyYyeHBT56emzhEUAmifEYSPqdSvrU
bJ56ubg3FdfMsxMUDJMeyBEnvcCoc6YbUqhYD0V4fpy+O5WE9RZvdFb89AEpSYVV
FWUkMa3mWg/8+GCiWg/o7LUlM0sRo/oJ59IhaOsNkdU/PToKdba28vLSgsjSEG2M
47ODXvxeDm5t1pNUprdDDiuNMyiw/cA0ghoeoyjt22j3p9jEi7X1khqts2YPbdUY
+OmR+sANtp4Ro1VO7J0nFu/nCz5EtnOi3U+cD+pP05yA8MDltbCkC4kv+41oKpEl
PX8INwMNuh7dt/iRgl1+CWkAlE9LHn6t8oJ7wBYfy2Gs7g0Zsx82pdmUDZ2UWvZ9
GShKJjQLgz79wIIvHOreLJiKj40wSvCmy3aRseSU71cz90rbdB2DT/jnouVgsjSB
o+lBFcSsZiAoWhsjOSX4uB0wDLn5Cl/GCuM/+Q9jaH7ykC++zwRwRZofRPmTXzqk
qB5VETExw4uB9sKK6XsOORn8KHPaUpGrm0oH3JfhRwK/+g9CceP5PAxweZ5z96oq
SmGbeGLvgn/VkCB/p+cpkDaBVf3lNDzffFOp5wjIAYWFGvKIUtcJe29m+SIghI7t
tuUtLuH8JTw6y0lqe87ewbDyhHWfahfrA+y8/R+JAyJEt6Yzm0jVS6EBpAnqudJH
7/YdKb+O9qSOO2d8M184/eeywOciVPOyUP6147L/jMf4DiNnf4zmf+9mPOMQatEd
YDzLBlzG8I1L2KL/pzmPDr+LWG/IfKgonR3egDpQOW1R2n2kICWASVmbTzuj4pL9
JEmD6v3DKOdbdgolXmMC7yMca6EVAiEZ2NZo+Mb3TIHEB5MDkhgue0P8WxtYhWa0
mJcSj5Jeu6SRtqafLzVnBiBMzZTorICmGddVU9tkEviMXxeOlxsNpgckpyS92AfB
2jWYT7JRlnOvH+S7XulfmsJDlZHq2zo4ezbnYFw8LKEt1WUWMA15C4kvjqGQ7+eZ
1YlMGCvXNUPVjGDcK3xq0F1QwHjP4mctbKlYsKio+BLklqONA+Yi7nxdg9ZQQBuf
fvKo8ll8vyg9iNbvkioKXaXBYXIFXj1d4Lwl8MW/cjOEAB0EPraW0ZUONNa+41Fv
aJfZ3aEpDtGe+cZ+SCKS3b9NK3W6z2T+03T/o9QSSTLfmm43jFufJ8AylKOOcFGk
2BBuQP1qI4YvEoYocPMOpHoUbT2La4hGGsz+JNeqexAVd6Mbty1rqGaoPwvX2Azw
XEfr0EyJZEORZtrRtD0ID8W4tGE5XNriOAIkObg5FbYAmQ2WYNmG1hvgxDvya37I
4CHE6Q6fj3I4HbKHCq/5+SfqIruZBWiE+4Gg8WDF+sbkNjK0gP57fLe/JNqzRDSJ
l5urQRXMgoYhXFBwZj6tR2pPFdQ1nqyhezGkpZTX13MCkUL/z6ju7rw3c1lH0BP0
XjkGbfZpD6+FpsEMTOZ1mCPLxfu+Td2ayyzjS6S+DerNc9VnH73HC8XkmnbJheXg
Y9PCl6bZX+3u8pgRkvpXHK68lxy4DQWQ1n9R8VUL079b9QW2F+PLH7Y8z4IGHX5A
Kgw4gqqOOiBwwpyX+nO4F0cbXmNvsfmC/6WruTxP1IPz1d4BeI2fRiKcJIVa311I
ThgSTbDpc5n55PzjjpjPSBH5ffNZEGlD/PTiFpnXJg+5oDEbXx6+bbH+zKRcQwDv
HnZZBv05Tqbd4i/wpZhrEBajaEpHm0IbRF/jEFJChvDvcWjqXm0BjyHA7m59whyq
2DNpxSrVIu+O7cGVPhYvDtLsRGdCOBNze6Kl8sPLiGl79GMH5JwAF8SnPntIrP/3
ZzR2wzIglBEx8biGVfkOghjozocBYhJIVKGwgjhF5zLAKOLvoguCyeFn9BIJSE9N
1oq9bjpUt3CSyQB7nVFoiP829ckN4zowQIEjAiw877ZLYdDbHDwY45dxKhEvgJOq
K+bBsfT2ibcQcTOmnpnksZwJg0mV5fnCV70kMCEzujkfenB+7qq16FPaR5dHqbFu
TNx6q9S9l6GPPYgSIbrpxakiie69jd5e3+pwOi1/OtQYRmCiEjTt0DjEOJJeth1E
Sb+zRzUEKbgiXC7KY8jm+daoZBoYlk62sS7lZ3eU933av4mud8vMl/jTxInQv3gB
5aT3kRb5Le2NHEKcSq8mDaDDBxHRR8f1x1wT39fZGyz2DMNpFj0lRec6H7QxXMpQ
sz4xPY3ta1+6yWkCva/CHP94CZyEAi41Ftug5fm2zZZQZkEZ4BeRwry0w5A4XjQ+
LVXmF9HXMuhQZ221VELFtH7h0Ku4QBiileZDM7tcnytnTA/TXz5XvwuK0dPjy7iH
0euWmSSw9qM10VI0b3saV2BhRwLg5rBP666m/IndokmeSd6mPbjoRudaOct3Hvpz
CpKmxIDja8FinWtXytSEhApUzHgeHBYD0h4o3crPNYClzNFITTDyPuektmf2YRDn
7RfKTmVaYuOSfgqZHLjkDzZfQFrzNSWxWmn0sq6swm40wbURpff6C85eymCu8M0s
Ruk2in6n1g8eao6o6YSFPP/5Q42PFzofbX4YC7+4zEzgsifo9s9X06bY+5hWpdKU
IiMX49Q1SU0ZaIYx9VI9t/L/H/zclYPnz0LSBRlpkutoKZAbw69Q/6J+MP4TYj7I
WXkBqiNDjVD93ZWRxo3qD25BukTrUCRSP11oCQq+4Q7nTnSNUPSHkPkrpDZ0LOKZ
zz1JEWU18pDIlX8YI1OuE3wR9Xg+SoOpMJ32p5C5NtJ7iEFXCYLI3G4qt2sCOrPR
8AJu1I9NIuDRFOclDozmV1unbjNPRmzE0kjXD0f45zVS7BdrePTEhR9jFJdMSBmo
6sh9HnU2lzzrEmr3gZAgwpUMhfgi537vdNCCqXS8YDPAVxQS9t2TAbeMrdXbldSL
FFhmcYlhFgOHC6jPh5L38ODVurJIsfGYcKDIptiNa0GI3bbG2F4xrDZeps5ZBXTD
lx5N6rOXPruK89nf1CzJAVterDh0MPUZIaQL9AsRuhyF6W3CEcmge7O/cIQHKWyM
DoJKGLesNjxbWL+klSxXZPtgIVgyhNKs5oOvYTWefKCEkpE4vaSS5qWGMAJlm9TX
IOc9mpjlpgVJklLb2LvBddDdsZ+l5bGhgVmeFmfLdaLK3DQD6MBnVit+xc+cbhIg
Y6BfdRCH34bNiP2DRMfZnl54SRcDk0i7+s5Rjby6v3aiQfxI/yHEv7Z3xEnCoBtA
hgM//aymI8gSB33u7WNtV6/8Rnq/AyOEgIjf6yEAhP1cmw+nZL5IalmYpqxauBoL
WU+9Fx7qzyZGfdeK6YIPOkJ4S8063vXYlZlraBiZkIT6DuMu1zHR7SXx3V8Xl6VI
WR2vhdVntd/PpQFj0fgdNveUv3PsHPoJVylTKeJn+4qXMY+tLwHENrYUpD03/jjR
8Yy9vHnjUWrjACs4e/FTpJ0tGUaxA6tcv0DWqXfSAgUBGLpTRDEXO/vCENDBpLrG
hYI3g9EjWOMlJVn5T0a35hCg7GTQ46oLETi1BQhJjSDnr3pl+F9kVjEWSlojWgJ+
Xp3lm/gvRdOrtgZJFcVJ8OYTQ2KTjIiAGzQAa7G4b9TMOPghOX2qHMoqLtolcfd5
Sku9Rs7X1UJqaz5/b4GyB6UbfldICdpdcvQrTxU7Kan+uGqQOi+SmBZSy2VEVLzJ
1n/NMjf/zjsMN3MXLZcFuBhSU8OqQqR/Zc2WIaR7VNmV3lS6/L5W5lymPjKOFl0W
IIofuALWKlGimTNtcFtxEuda8Q2TBYlBIYFWyHOqr2jfogjY26lkVRb0wMkIxBzH
bsedFpG1mFAEDyux5sX8X7D0Khbt5lcnnfUCTzvPuOzAXoCHM4BMIIR+qmRFb7sA
TgWukiPV4oX1ekMKFJbWXmpjHrFavKsSbu+WUHKTtvguCMzpOP0dNYSaTEYiY8Ko
aPBNz4uc3wCgBUveVjRR2Jwlh0n+HoJ+b+NVfzYJ80/ISVw2JafelAQtNPj6ySsB
5RbqoGV0FygmsXvjtbAfLuLWae0UuurjRUu9boSoHS/pGXffIDLQtdY65dn9RH3g
clKIX39ENK4BNGFfLpyDCwug9Z6itiJQBnBpMMWJNm30Okxf0GLDTft5Amqp5/YW
ETIJKuag50E2lSQBPXFd/rNdZS+WVGVtyx6gMd8v9lJc9Qj0I5qorcBaaalWXLMB
kmJAt82/f7/P4lGlwfcJfEmtBEMsGpVbhda1G4lf5j1gmxqB4DvSMnKsABwrYnq8
ecnUkP50TKxSRDW84TtkdsGUQ7clycepvEQLnoRntxrfbYRvh0f7JXvYZbKbZavs
xXPGbQRziYiyXlR/4mIQzjqIeBHjqKsNS7mawOFkhfQf8fbWokWKoAKxF8uNhS+N
ny1ozjWB4TAW1MANisLRLN7nE89KXxFkFiEJIwdHSfHmp2ZE5HAUiiTL6hrEm8dL
sxNnRDUNrB6n0bal7VxfzpwFkNdMbT/FLt5Mz62j9Sg90VsIkDgnNjYZMlNmAvl5
o8kkVLRdhh9EsfXbIlXK6Cc4V0O2QPI9lr49jJD7Y0wyMotKlyzJPWDHsuy9e93e
dRdhfOUQYRH4Dxhr9gaQ0pwScWVPuj+SCcrJCn55NsiYa2kz1GGbocfVZsGvmQPx
HYsgdHmlFpStpnXXypttmObRjkopsLwnmgfxR1Sjx6RLmhW0vDpPB4WRA0idwqYf
47uovBsmXbn5wOIXE5ObgXXPnSa0IyblUqFHZ7gv+uG+bsg07NHKHyzEddGiM76P
+pd4EVRrAV8LW+TATy4k5YeLSsh10qtAWYP1ujHKjwRcz9KznXQ2DSSom2ENhOA7
EiZ07DNvyDDz+O4f1q5xZVZWPGl55Dhicq8JSB71jFZeZ3dYkDxnmBuDQUFYvNsH
ypYnDA5mZ80ZZFzTesTw08cihQ8X3VHt/C7QqojFqVuOD9VsokcWV67Nf8sLRRlI
GUBUKLypcIiScmDNRYHBfHtaRTjIAFjOLXnOjQM1C70bqQZbDB493qQ8NNoWtA01
ccPx8YwBO9vCVsl6K+tCXduUH+26hJ1xCKTCrZfnBYdlG9X2OP/NhvdGeThxUNL9
lnmJPfRN4J9S3Tvyu0H2F0Dl6QqMNX52cU9HNvYtr2z0sQU7DbIsI8zUmLaXa41b
intNyeMKGoUT/a02dqPnMC1u986GMjxSyH4fob0FCMOSqMqy+TDzEErJmLVZkYrx
LXVIsYVDNLFEBYO1Brt4a0TMPyj/KYDYtWb7Fky+UJ5nBx5WKFO7zBIjFbbxwhtZ
a0qkQl/lBD6ETo6wqnEux+Rc5mxGIzVjr3cecwHtHQL+bH260i/GZSsCmnRCvddT
88K9Xb0KLjd1H9Z9RmvE9Kd3ilazaUHB+zRs+3GHO0PfjmA5rccE/St0p7qaSR9J
AKZoyIBXS1Yp1VXViHMloqEoYt2dGtrIu2UGgCrv/BCCe4BtTTzVu+AW0FdR3rB2
zqGAisQjoUvnGEWt5e//roiKGB/7kLqmVxJjT9AaLNeE2tBrqg7UoguVlhUFU5fx
54dgCn9a7/7gt4UwYO5HSKiEkUpXSZskiEeO0UKhmbQqkbcIvVPYYBlIEg6UwNfU
dytydYyniEHWRHCw1SloMwtptE3h4qFJ10q7oc8NRImbQgLOO5IOZu7fIR19GiS5
DnINBHm/2u3+pO/vQ2hHxkqPSMXebR2IWMZbKjhyqO1eY7qdbuJEvP0+jWP2YhFh
VvXA3eYM4rCgenI9U9bU8mIrW0NrFh5qgkk1PMzhtoQ1oJhY6aSwe8ozU2nw+L3x
Qaw87jjdHXzNhk2SEwJL2O9Iga/J4F1TwdQ5hrajLmLKlw21rGTPygs9fdm0wgKo
d+J9EZQFTfp1UJja/YvuHkksLDTLdwfZ6vAzLqK/fxWmQUJYETBoA3/LGeqVlwVP
lgWteJ/VNTZ7zkIA6KwOgIfdkZsPqrJ0AEiUBLng9I74CcZyumSjMYiwj/qtl4A2
zQRKooeVOW6372x6VgDHpz3kvEuLliInFoGspG6cAzxUHr/pBQWEoMSvJzimg+n3
HwUJUvU1OcmTZLIC4/oJvH/NrXgOTuy2gJ7Q011qzkAeqIgjno13/+8EpS90svqA
7ner0K4ShE+0/IwMRam1Yqr5l4eQNJgBt8S0uqJQOGDsf3bViMtVL51osc9o8dse
tdV3uhOnF0J8wDKNB7KHFt9aA5sbYCmm5HgvLamvAFzmgCSams+R/aqPbhZHGDrD
mpdq1grVjKxZmcDdvBlX7QZWBWZMEs/Y5IqDxI2cKKCFRs6xrOrzb9VmCg0PZW1w
o2Wxzy4XgmLkfT4YueHMEljSE1nQNkXbfLJeTyiYA8ZcCx88kcdQ3KXxkwxNwRZR
0bZ++oG03Ttv9fJIYjmX7tC3U+ZfHv9/cSY5rvfk5DSonUP/eS/dOTYREFLTwNid
Zg4hqopnb2+lSwoQdj0Z5SsAQIxZE3s7qdsAfbBIXiek3z1y4oXijD9zKomQqSkq
JXy734rNYrLZZMWVPUanMpQ+bQWSe9HyNsuJxDuVwUp75zqLC9sv/p1jpNubK0Ig
JMqimPJHv2YnOrDW1FF7eUlEViW6+nPDj83lgM9Xhvc5qIQ5TKk+FSabgG+i+jcQ
Btt3kQaUN4C4Cj57vpVkbgbXvMQE2HL6UVe51VYMK+CeO3tv0hX8VfxVr1UH+QfT
ZaXaWzXwF6Qud7VhZAoaxCMioL/xI6UtJq/FLJLIcXKhavM6j3pp/vjtQfY/OPW0
bTGbSgqM3RXvwWb6zXP9rEoijp3kHEAGl1+5HW9OeutL0fVVVh5iRNYAc663BGzd
xaBOjvn47Cl5dHcF2X76G4J0GnnswGMgb+7pfO0KZmKrmTwpCpKSQ1aBCIb36Rti
uPsNM86fl49DfKNLSttDdkvTHTm1W+Zc5+pf0tbbMtUMbBMdg+GJLv+i7uFUa4nZ
lxciK/NOpd+ytKuOgQWXCKCPSKze6r2XKAWKpKSFK5sJH9cDdaAT7Oic7ue2y8Io
Qpn3PrRr3Ka4rtA6OvZOsU6u6Ighs/lBXK6+SOmJMclDRZ1aCcIOPjWo5qtOgkjK
28Zhr24VUznEiey8DtZGwonBYz0nVl+MGX6vthVRq8EKwYccnzGF6KHpC9nMpwf8
S5tJiAeF8E3j3T0/UnOUI5icVsKUIwKK7xov/FLfLpvS/DkMUwcb3oQXJL/+hvoW
JsQkPAzLsV60ZVOE8Y9bbEuBHnijrI8mL4yd8ZTGMDyhsD0UHZgBWw+do9F09uKV
b4Cq2z3ZBZkqOVcr0yfTpmMrEgcAbuHiS4/rvbbRHJU2FyAvLDcNqtFgEO1RjSRN
dewoFxU9E2x8YuyXiTLWeffHwzCX866Ejt8JLDF+sC7zU8Ljkwsgz48A3M2UBeOC
f6H5hKakzguGKv2e7q239xFoDgMxmF3k2rj/dBMIF26xwKQM3uZNf5Wh2Gb0ZztZ
91vkNUor2h4mdRj3ieTXGPgsjd8o3mEgNtOMzkEysVW8FpOMlU/G8X9n+s3nV9jK
u3oNF8atMRevJGZHeM27woE4F3hdeWULds68XZRvsX1IO1Zz33zU3eG439G1YL4R
qFiLK15BYCyG1gjE1yLQBcJxyPGUJ5V3XRejjdB75wghWbPaQImTG/XI2GlyINC3
iL41RtDMY7Lgnx1Fhm+YIkP4btXrI2KB2mEwsBlS0TeU5sdIYF2k3OOU/mH0XPI/
3Jb8XPhtGoc8ucQO9NuCwMte7htF78wAyHtPIlLY62AOqjYGVOLceJNWAehto3cV
duyfvh/lu3YhJSB6A4UbLeCvudo579ZZ6mLUKq8wzkocqoi/jwUMvDaPhPo2mqsd
K2QQOTfW6Fp6HUOOqSEYO2NROCXCFPGCGKPLodchorru4A3WSqDc/KyWA2rTALcY
1Xz9sKamAspaX5XKcJFAozkMjDCoe8iL7WgIjDnrmAXRuzDOfI8fEzUk6wI4k5JU
NUFTkHPXSXA4oATvyD082xmVUlpuC+xos30dcsEUf+BLclhGg7WW9xxoCQ4OAvpo
NMIMRbNor2SndjUNOu6MZhlEFWW91jMZdnjoqrI9PsvxV6uGqJH8fe054IhAO2nm
UqaiCYd0AtEfP/XTpbS+NXY5G8EoeRf/6w/AJ8JONTVhhBJHk5GSt51CbOy6K5ce
qrG7996R/kr5Q6fo4axnT2r5fTcfETUeI4IY+Y4OvhE6dm0asj294pr6OtQ0Xxp1
SETSMXHfyW4bvxOZAW3+qD8/Xae3/QMCs+5nHol8xp+GP+2R9p6izzpHu7Ixoiqg
Oj/5XiThOv4JkaIdK1b2Z5ygV0GhPmHdIK5k9qLqjwxpYyeRNsvlCqb0cXOpd4b/
ZM51ZzpQXmU0sFKctf6UqofupZB5mFzjCJyViIrpHjbMaEb8lEZjJGr7zJUZXe8i
XhwgQfcbEifg73XlcLf7gqnGkiuqPLfg7hxFLgS53eb2RaVlwUjRrPCcCv7kn6RG
746cC+6I4CA0NYWrGW85obDtMO5L1UUaFN/1sk0jSqW4yAIvHp/V62B/TJHvP34g
3yHPHAEMMMu8XWP33GnP1/QkZn/d+BIwviGBid70Zff4NjVIHVYSjoh2FFcVhI2n
gFcNNr4Wl2XWpCqDdge4EC/U2+RBGBQm+lNeEKJSyuuEbJwXxlnpHsXfJ/j6ko9o
6kHG/piT07zD9Tq8hXb6P6iES6fmJsRc2/FmjmgAi+Jm8uphDZdZndoGohVrsiI7
pcBOVZ0VWgRZ5odnPdjsVtfBCxo/k3HtqJESJJu0kc83Sua50ysYc0cF2vWn9z4O
pZKQhi8l6UBtLllxo7oNSSITgx0ldBLcCmcJr9OFxbuJCTEjV7xbVxhRtUTJeXqi
uI0v2zLbOYQeyod/YiBQv5KIx4xOJGK78vNEX9U7yDs0x/+ANuvZmOJW9kG72eK7
tOSUrUS4+6mS7FG7AZzGz3jEFl4cH8gY0/bb1di62RlCYGIyqU7xfurCDriY90mO
cw25DE5aWgkUeKs9kCRFqPpheNid290WELC7KiljOjedlGg+fy2nYKXkTgg5faC3
G+I+ynTatpwmMKN8YwzNv/3XTbn7dfuAKMkzoMPp9W0aiNvxqUbnJh4nT/DeAwmw
tYyJOc0BpiGGFCHnsKe5EMrf2oJaMDq0JoLixtX365wHsPA/CUkd8cqryNVUkIrW
N9kYhSnpCOD4FmIFi5i0vgcfmZm0eNQASZ1sbDElrzPoz0V5GPbp+MJchDzRfoUC
dhYRTqJEXx0NNyAGNF275hCPyOkGC8Fc22B6dM6/o3lC10zNla1Cp/nswT/Q3SyH
8DIX4Ii/Z9FHU84QdAT/YelCNX7SYUJTS9a4Md5BczM5vNYmY/1CkUaMUzE6rnxh
G5cbvVv8/DYkfAtjVNAtwqjGdAMuhO8UdVIofo0JC94rW06gZnxFEdwLZeOKOYWD
o5y1mYPtyU9HrT41KF18hymVUBK+RzmpeSv8wESSdll4qd97KRFpKbiMDO6uiAmr
vot5iiKu9qYGIDLO2x24F9LbWOUoaFG0rMcIUX99Eqv1oUYf1u1A6vFCUZkJ+PZF
u/YvJ9J4AUR1hiXyL6KSqQ/CAeaa0oVd9oNMAYQXkU7Cio8N7QDlwTh2Z+RNz542
ItHBQj3arp/FbixCBHC8W8aV8KOd4hquxvYDMEqq3LHM1bDe9yq78JfWy0IsG3u0
oPSjFq2+gK3KXyp4eSeIogQdRVcRJr3DXndfdbm/E2vtU4KEvM5SMhJRDVGMBBWq
57Tsrv78V4LGjLdrNd4rx2VOEk19mWlbaAjKx//SkDdlYRwU900G+gX0RB5KYRSj
Fb4/u+Puo8Mt1N9XjNjKjb6aVZzzw8GnBOaUzUgGgynMnWNw2MHUnFnyvgIhEoLp
49visWOCC0+zFj2NVhKzGrz33GIWPgjxDektpWfdYbpVef49nf1XOFcGX77560WJ
vi/BHBjxDX88jWQRHi45NNXb1om7O05pk9+dDddj2Zoz546IrKHEvE7JVnv6I/Cb
rNP++ZAKBRIuLURvNQYKpXeaKxY9so0Oaksb7q3Vc9MQ/sIwYjxUoN9/2v9kUmDS
TUiPxylIBUQvTAdvExVXKWtNeAcm56pRrt+xp03TNxoeUhP7TUkXv3855aWP3b3n
eBqyWU1uydHFOAQsrscZXPrm6iUIe5wcmWERqRKqnO6FGS6E7c+tQlnDCZ+5/Ktr
MZlBKG40JZCVZNgHteyZG8CMlAy0fbGnkMCXFwpVQ516x8qx1WDivgjKipTnWYIj
clUQvgX7bq9OitSnQLV3qjv304tc/6sJqcXgfTVcSxuMintoZ05xlGUtRfh0WCwy
DzztElhx6hNjaRm4fNC23qqw0DLu1QAgr8BgOgM+W8jcrMK5/BQD/222LLIxeGoL
fWG0d9neDGgQ0bT1mYHrhw1fcEgn1zYouNfFD/zIhF8epV+swMnjQ8u/pGuY0T9n
axZxGxq9X0UpylXroDWLCwfqUCzEEBpx87OO5DhNlxJXHKIXpDmslo6LXeuvwdXD
WjNqCmFkx2umvu4Dfadz6lZraZmphnJXlCQB/QVBiAvFofUiQys9QftEBjD+LsNX
aXAd762JD4kCKC9hb9R2fPVfLXTqGjXUtMaXsx238muzv98B6tD7G4s/78InOojl
+c22U9TTXso6Jhn5sgcTQK9zJ8i92syeSSiyuHZ9vel9sngM5tA5dGY51XQN0SOX
VrCTmMuJcwXEkr06fOnYw76BogzIDAVsgexlZiFdiEKV72TjdCP5twv2/R63UcEN
egvRy6zxggKeK9vqaTStA9GoBuXgy+bpZ08NnWkcPhF5SOkWxcXtuwfOidDPAAr8
P8G9WRqAPVC/B+dMrMxUwWgXLJCWiE/ERfhorM2IsVT4LMKYLbvI9bSZmhO8Dk3O
zb90y/HF0eNqJxuqchGtPgmNK3X64G7CNLQ9FDwqxmKZSQVc+UuaoprPm72QECUC
+fY29e7HyfTsjnquPLBLZwxKgpqhRhRgbBHhQGIA4Z/4vihQnZwgjM/+3mEcXXDR
5Snr2BJqIcNcytCGLefJ6Zp0tRDSMP4fNsnrmVi3/DImFX4Iq+O4icOB1+YFLVcP
H7xZjfK31apHBdmpGVIkgJqI4IcJUIGTON3k0Nt/w5PWZ8hDoFwVkOi4aynOwOV1
u0646qDdKw1Q5gBArAvJTWfA6eou95k6jlVyJjWyl54MFUiZxr2JNRnzS2Pbz3pH
xxeFMdh0ucNw4trZBVsY75mHxmlt/IXU6qorPTQr/5ZyrSeKi1VdbnKXqbX+GBFk
XSBEPF2w//2V8c+OuuTQVAQQ1N7zV79k+LehF5OJMn6sNBNjqg+JI9ObMPgsG9re
LsnJwohI9xvS/hahZgwBGvjStd6uSC5LyIcV6jqgepdp0+wJQ62NyXFUvbTKX+Hm
1Tcro60nt7CmJwfvWAZOgCpppnBNU+KV88HPEmwEZnx+LmrnfPpIgC5F76XJLoef
0veycms8sr5OnZiV5g8Ho4rcqZU7ayRGPstHN+A2S2uIYhhoTLOhvb5X3lTcWdWT
KDpi7/dTnllcxpCTQPygtxZiyNxBtHLBYvtVX+tdHsxPYzXW+UvVKwLjngah1cXa
1NZDbWQYZwzXMpFB3sBAud3abcbceoXOKQgl59eRK9GlCVK6NsgNZdfbLEYFqTe2
RQex51wVxZCCLwz0HoB5BsBsIr2dNhw7AUU7k6Q7psWWc6j/u0e63uwmUDMVcezK
A2uBiMCHaBcGIVJvRe2dGd226+RGdSTzOflfkJECsSxk1YZix3yoIfd9V2Xqm5JI
FnUq73LE+5jlfpkSHPX1q2dLXCM8odcO3QthZ3nuTjX1Fe7EshkV2dfGpDRI8jX+
mkK124cWZdHNbJSy81wD339yu3lnJSGdNCtBi2UUmIzm4aPLInwX6PaqVWcMiPDW
yX6x2ahiTXwh+Duszhiriw2n4ZyyCnzaCyRNFa1yFVkgPE+gTzIo0TVBSVRE1jxB
EabJLvelJD6B7NcFwW7DB44O1+fw4Qpp8nsF9sY98nj4jkl4JWFgQo8VzMv+RgE+
47Z8DT+LUno9CC5ITbqWnzW6zwPAFSSrFREMZklNfgoD/tu3lcK8jJ/ENJRaab+J
S1OpRnVbrz4kPdGv/MApANVfU8qXNLpTVSIAgtvd/IlpgLvRmI+60P8RMBPx+qFT
ADk6vcGWB4lvK7iXQf+E8SD89ggBhMoLS+wW1AvWbvha7rOE+A44CSCs2Q7+B1jD
0t5e74vBlUzKTLFJb2Ki3vPUSlFrA3x2Q7vuSfOTGRqSzBgz+XA89K/6YvEMsHa5
xI2lfBX8n/7PMBrOTnnXERMOVrVea1dRBxW2HEVNghUrLpxxSQ0XV+l91bg3rXwV
1H/NEysvCR0BzZZRLMIlFBvUd56aNXVHmLDQFppH3vGSDssBIDeJQq/bBU0zD6rT
Gcwk2KD61yIfRBSKMqI1Fid2EPCl5+yM+t1SGfNOGzAnrdj55bSJZaz+druJuhNM
kczXiP/rgck80g+2oHnyj88m4n2yqviQhxJed6u5WNQPuIHS+qMzP8zDz8wRnPai
0qiKwSxubeXPCvKy24z+2aeuufluLgM1BLsYQgzm+OpYtiBrVOYVOsXIqyMjepVw
oNH7bb1QJqyG0kcW5iXjYVJzyiGJeyshUQpICNIdQXynT39CMjLZudRTjE8O8jOi
9HMLVFYhZ8KbBbYAhPY/NaNewFQ0wRY6B24zOk3LdXqj/Pf/e6wa14rRjx8VsM+1
HFGv1qhKFzl2qUbpYHDR32hH2bvtv2Hp8WEXuN//KoGGOIZiqFrMxhVwz/5cC6y4
+J2+LIT+LEdb3q8w4RpG93J5W9lR5L9h62lP8z/xgfebtGbT+s9DBxy9MKoNh7ez
kPVQp+QG1J3F6mPOhmeeER040g0Yx7aAs/F3SLiLhXplmCC+FDIp16WS9fqoxfRP
ekAQ3eRVblB/Q/HuwREWorabbw1eppnPl0AZGTfHrDvUQ6REDBqToV412h+6iINh
5qdBB+Ej85wJGl9DdhH+BJ/IGzNbKwT6pov7bDRwPRSyMs7My61U8fkCVNzWWjui
6NEWOxHtRvK3Ry9uneK7RWIyxirWDEpHlLYu4kIiUiUBkYcHH9CuDZi0K493d0pL
kCiEBOdYGbRLs0p/h8El2EanRZkua13K0B5a6xm5MBxJciWDFXq37DsVSH0s59ev
xYT5bWi3VfFUmX4g3PUQbBm/FnS7BUU6bOr77fvz/oVEaz2BXOWToVm2+1ory/AZ
SAHhcHigDtVr33lB7ugQIqoKhhs7qPBsK7ZsQMGmq5zuU3UXib32fgrB6P0b0mDQ
GNBY1+iXRRGp3wgik9n/R6fO49P9HSUIA5JY8399wUDl2XFfy0a2SB4horVsFxlN
BpTFw1spH9nNCsI/f2A6w3uI5Ihpvntp5zt8RFBxMJb08VSUlCHJl/jLpaCVLpq+
N1liedJjS7fr2N6WJomJR6mm/JTV5VvozYtQOSYDRO2bZ/jqaCo2RbNP1b78X1/R
JbO0OJue3Bz7MT9zyWo7w4wG+y+DpZqYG5FJ86Vrq5xxEIQ/BOOHRoVN1sO5U+lJ
+EnX3ySavjN9uXwvXOvNYWWqZimvGHKMzFvV+76I+zMfA67qonb4k8pY9jw0uApm
cQfPHV/4GT+yf3jDSiGx37nm3DR7rCIV4sWzzbkbWAthFeAb5jzEu6a7scHcqpJ7
tBPR6GOgJDbnbHwPsps6dqrmF0Y1Sxr/ibWzfwO4vahdSbQ+/04Hn3xgu0yiztSf
Y9ZqBQ/YgJx7IYuUfm2KNQ+anuAo6WQKV+yPwiY5OS5fnu0eHBgXw/vIMzQuh0gt
eQTfG2H2GQfH2+08DxI19PJSh98yzZc3jp/wAg1H+cesmf9lgEWQQ7UX5bgOZU5T
Vho1fBcP8KJdkhGVoJT161glgr1UGS887/kOa1C9e9/ug8lOSXITeKXdPCBRVGWO
thIQ6kvFFhuCAbeI06OW+Xg0x45sGCcEtPIq+Uq+vJCfueL/Whw5cxcE5OiOyow7
6mCfb/8N+4uYQNgzSkIhBcIA5NOA9ts5Fi8itQssGuKrunFTpagJ5LsRiSMQAVvw
zAL2ecaws3h2J0Ds7yJf71MGQ0/PFEizZYZPQPAW2m/y9XwAplG1cxrMgHCdYKJP
bSuiIVLgGJzCgwg5Kx5+BcFFLNpQ8d3OynTJSnBOvIRGGLfQyc3RnPOpWTGPbomv
dRQBpS5RGL3J4jgj7EH+7nynvNlkpiOAr1mSpuQgBVEz6v0cH17/3rlUaPOqJbNr
2lBALBoF1JkimLd6y2VfzGmyxhHsC4XZ9cercRRgTtykb7RI6N9v5eJFqGE7Hz28
OjOHuicuwGUgI4Sw54oeTa1Q0XFtn8IFCCve0VKzBxnB9R+3Vcn8ij8LPKf7Lc3Y
OGRzP53nKmXVsTd0M/eqyhBG6KcPPGPVVNpUnvjpLjKcn048nItGhFxFn52j0G08
1M/Mvj/4Pqff3N4ukc8YUIR1vihf5nbEiqUZSv4GNJXxzWAPB6Ix+z/Aqdc04fzp
9IYXieS2Nt5lSdFxM8ORC4cipSEEVEhHcyrXMm2e04iFMnDR6w91XOCIeteswh8l
QeMlpiw+S4N7mAd3mF981R+RqBaVxXZJ46wW6H3ABZ2UXIWljCLB2Z4lFyE5W6H0
Qq4pyZi4MYuc8oHcWKKnNhyvAjafZkRZEoQZnuGAdw3mEk12CDoaZv3/A75qIF0M
F4uJrC073eKOoXiSqE5IUyVE41HQJNwhn3qZBGcwZsg185cBb+hPeVNk+7SdAUIX
a3rq3Fyg3bAsUu3juOlMlO6yDaz41MDW1epMXvTJPH+ZCvAFaGkvwIOsiJaP4jMB
emrQwfSip9WEpZfLkKdlI9Ho7Pa8Frv+5FHwT4TFvvmNr+R0pEs49dWY0QJEsaR9
+h7POBm5PLeoV+BaZrpdQoxfmLt5Os7+lU4SOVLPxMlzMllED4AKRvZLrSLyLB2d
1g1Kjt1HJWt3eGexFrm17fdxHPD/4GamZAGFDoCcCytYdfLnul6BwwuEWgrqHo/m
C52/r6bBKK6BNc4n7KpB8l8Qnf/SSKAO8vYMzPLRw2is1lnJMhMNhIpkLMauwDUp
6vU5TYAVpKov8XdVOGdBZVNj3NDU00lWAAeKeCIXscgc9UZduIYXIDf3MfhBtG/R
kmezbp1oF+xCyAseJnn1D6JJovS93865XphTt1cwBC1bibU/4rWopr34oyBuL3bj
oljnzcCa4UyUl6/UGeqqBH541PEhTDclwBjiuJrznWxW+NiJpiUKYmdHaz9cbOn2
w6epESdz6aMzR9yclHkM22sIy8/I1ARfgkIdnzGKRHzpaF1AgaKlEPxHAS0xb5wZ
9v5KXuy69L4+b56sTU6RxmTbJSpGb7DrjyMHJBMreoLeZeEGdwuU8ujSMNKQzVJH
NXr5LUC6BEs50hg2Z10cS9xkb6gC2zg4dTjFVt+t7GQvUe4xwmAAa39Y5eVEuGba
w0CdJVnqYbCxSAym9hm5TdiAfVKsB9RRA7NV8XqLpCKKrQrvutWj1r+PPkfxf0hH
l4YuMfDWjdc5G8T8O94FRFtrv1Wy/9rXRST2n0iXttcbAughhn0t2kMrtuaNrFno
6Tg6tJBiDfs3u8Q8YEOeqt3XtzS7aQNrDCVDQtCbsiW5i1xv303lrNz9fIPLTZKU
yCM8l9zP49qLQaT6+eTr9h0faLLHN/8whAiFc7KN6NLdVRnMGkL3TGZWz5dGm/Jz
MrXo9kXnnaFpFEqpOVXeFJN+3yXDcGq12EUTHpCZx/DTmYk91qPv+TOElEvbbsjz
F1cuUBIJ8Ey/VLRjuAJ2uPChMkRu1elFBPuzhew/CEhyfDkQ+IxZZ8Ee4ofXDj3P
YqZQ6bx+W0S8g5NN0PFMqknXm7NhFUb8HR7o6D+g/1Dcga0pXSt61ikf9mVPR+Jg
2xJ0xs2bumpnYAnpLh5gVVAhbdmwbMdcxSlH3HS9QPiJ7Zxt/hjijJofrc5ezLDK
cUsDlrNsNpi2W2Vp8A/3vilNcLuOD883KjHO7HE6P85BFsDfp/GJa7dFqTbVIuQO
1OUPMyK5EG/Lkg/CNtI2gdeu0qXlY3fctuiJLpR4qmPIqNH3tyJktIyZVKbGM4hd
bxoGIfUbU00daN40dK6mP3Ma+paFMVeyyTbTkvoa19PAfkBnJ2dnYSzhKf8VHOVK
7c4I+iDv8csnZPCS8od2sTK4qzZvkRgmcjnBJHh/1zuDfjia68+Si9iEH+V4N90l
HbIsTaT7sYAn12RhXNEt0PVKMWzlII58hrxf5TVmSVCxW3K7C8SN2z/IBz44bg8/
83woVyTt/tHQL7SJAEXQhrbrxj6AqlRfLl8IBIzDuy79qTvQHz6D5GtVsfcVfCwG
ylWqaQc4brnmG5MWiiaYXaOJWB+MQrqUKT4zUiCgJ8cj1Ds6VJ3SYOCXA/TDvx+R
u5xKrlA09U70oAvOTBHszo8TBO7Y5JHg5fEabVrwQWYjapwUA9BAZ5Qv/a5oE8nr
abAT7r8tV4LKTO5wOombx0p9a7SJNrNXAUYLFenMIrb6k6XW4jlgyuTow5oh64Qg
UNfx4R6NSjDfj4T5pmjuzfwZW/mgko41fU+KkNTARvPMyq4hHj+fIq9ctkreo5nf
JkZ8G6oPYA1BrlnimEvr7MGjV8683/o/8VjVjptY5zYSxb6ie8WH6NRmTmf+bPAf
/QuB4ziv2pGNgojNOmML616Aff950XOYAjfucN7M5bA71ocQWL0APeCpJrUi2/3K
g3enswsSbiMgKCxSV4OnNo4matZBGTo69PTaJf8mbx8wMVrOD1g031hMFdRg/GC2
AtyerVsTvNM/fFsLgpZtumQ4hl/BzTx5HKQwbGIA72PXEIUcOjGy6EWNTJ1gWwDb
DqXcP8UOBvAh1BDP6Z4vKEU9iGwK1h9n0XDpaE7pLl4x8Zqkj/aFjPxc7JxZb6hZ
kSatg8rJJpkTcB/7wBYXNmmQGz+tHPiwcHtiw3lXTpkNxRIoaevlTa+HSw5t4Uam
j3Rn4Up5xc89u+Oil+mdbCQqd93RehqZhHeT6ExsxoXJllLjmyoYowJ0tJSX9loM
MROqWgD6TyO0zTun7Sf2ILNayGb2jUZ53julGXAnLFkEY2woCjokwguJSvcDM+MC
JLodpi0CjIg4crBa0uK8WHGnTi/UpbexGlnlqaZCCyiMaImG5XW8NDo4qPe3+Tpa
R2gUWdSEkNZI4bBOGL74z7LDllxXzA3qd1hqfM6fqszlo6ICXpkBVFPjOuLdvFKS
JyzX+bN+xNtLGp2x4flCsY3kXUSbnGK9D89bfhIxLQiRxBQo8GW9iDWT/FpZMtIW
AwhMr3XPmrfuc40Z+tn44fi0N6BLCKRlwY0BF1s+BgEx+NLPK71U0118j6s5VAqN
qbuDxuf8aiDkcJ0xUtX5eH9DZiDSJwbu3rO1gImG5oI6J9Quqqdteskvk13xKAyo
e5xWYyz+L29AB/Iyl64cJrcwEoIMQHBtlt27OCGXg98VDLZjaxkJCLlRlA9Sep8K
8txlEWPw0zNI+yrEBJHCuyav9pPsoPr1+EhyAfeXusMrrlTjIj77Iy80nn4L8bCJ
5boEjZF8YHncLlaSUk6XJOFehgAh9r3gudNBKgHOETxJFcEGyCIwAGXLWnhXlo7J
ke4n6jQZQsPRiQyW46onxfu1/uQz4ybkTJ1ODp8qiPpompHsIHeTqgi90Ui9OC+/
xJQBQUA2lS4W5oYvjWjdnNIKJLICp0IaDBgm65H3oGShd+yNxg712Tu9x6lqA1r7
IoL3eXyZWh/no0JynJPm+KuZ/lEvHJ6tjcUe12uiHpSCkv4BVhnD9DvnI8iYpyQi
AXWPfv61BmD5VrbETOAsqgOigXq1vj8DHtsHCeN7MvOAnsXWSrsMQVfXwBmw5fWS
sycplI3gPsSWn5gMCPa2jkaWPhlmqAJ2rvUCH7pMKDV7LSqYyicDYNSMRtudfcYx
G2GY2oSPU7eAvhPKB2+ZQtKZRlP3KLQ3ckmj+AE2wAa0N5l9z/1GkV9X8qap+Rbh
leL78qm2LXdoQJjG/sz1LHV6KkUdkQx64SjLPKHpB/OD7PagiBHd1xbPvOTu1YF+
a26zptEKlz5kYeIMPrBsWD7Rvz3/2xPfh4dGqA+JICSMY0213fna1bO8RPIfOzzk
YcMLKplzTeuFJ/yJGx/eTqwpjCxrgtKfFYR8s76iVWCL1JOQlkdEUSsWNeN63TNN
cNJuyApB5/kHHSeVLw1LkNWFF0gfArG8wvJVy2pyHPtxuhuJaolpYzD+0uz6OW3r
5VeK0FsOFTmKwmXEMZSkZwiVY7cvx2KPYTOIpUac/5CqWkMz/mc66owt2UKMD+gZ
qqat1PzQrPiny8xnUjD8X61ksThBbm3hp8SNuV7bIlrLpwNRFOh8xMoY414D9Ocv
Do3ZWtdNTnzcyjkLrl2YV/Tm7ciPI0e7LjZNdTBgoKxvwgzbco8twjrsoz8q84wl
8C3tSUKhh9bq2QKuATtYn2nv33N389+cioPEboHIHCUQC25q3ph7MYWxBlrjHH+c
mOoOp8xYdagwSSEk1d2MwbI+xHbGmXRS26UBqvR5Q1I/UYTcwdYXFOZ+i1ZZ1x8I
h4Nkd/7Z076J/JyXAh/nzH6+tt6XrtDy5AynRHFH+EnnILvDIZ0doksvSlRYWeOF
xRX0eG8coWA4FXWmyUkgQ8OG4UGHbTPUAq05KUzbIUzPtkDqpY5aRYDoErSG2hRJ
BGL6nsLAGMNvgRCyCibXhMPovUpAP8kWsc4ZhJHVdFTpNnTFnm/OneRW4V8Ssi+T
8xl04Z7rp7Ma5miA96H3BYIj4x68rU5ezzu0bKgGaeTzv/79y5qso5SWIfcl3RhE
BSF7JwS7Xcr799En86ycfpkK7SNRtwu128aC/NrdOYFVa64IEC7Tz6tRk4RHHN1c
no5/30ntc1ldQwPtdrVZLY3GlEEsUzK/si+G8UzebMKxbPaSytHpkIz/P+ktCG6Y
zHZrKkxePe1DQEb7wpLKSDni/1GYxY632Q7ga3cKHVBvKaHKHoSM7NoB3tIKiEIN
EqLZ2VM9cEiYogLDvz/mLywtbiJS4frXpvwcZwk6RqjSe8LSSzJsz4qSf4szF61B
eFfvfgFKrTzLuOO1YEBzq3FJ3vY+T1EKThP6opTQLPr84GMv8aC7AEGvm7+eD8gN
5QPLdV4YTiS6cjRRH+fTz+zuyt9Wjnls2Mnt9zP6o1LiZfRi5Vjk5jQSAu+OF3Ku
v/vvGD9QYqX65o9cIIylySuZbLkV9351B0iZB5XLxr+YRBSDUXT1OCXv7qHk1lMH
Oka6yHt3u+IgKixDeIcoKOGeU2of7fpz20cAaBKOdE6YN+CHmQWMtxxXU2UOPZLT
NIATBJcWfDph4bp3hNb5nze28UUBMSXHh/Te/BmEptmC0SpgRMgBs2ppAOfEvBqR
7lEdJmgGMUiEtFmeFtZEKOIRZgH9RxYltpniEQJFLaQQ+KUZ9dLFhVrA42oLXx8q
Lt4+VGX45JOD49QvVXhv/5wGYUz6fPyXulsSjrZZxn9rYdNynm4oaBheg38P9BwJ
LKKljX1z5rtkmfFG37G018rAVW9uGLPGCBgjbNPFpY7VXM8nJXqUm7bgHvHjdI+z
3k0lPXJZa4xKzlw37PpmguKv0k6oX4mZ8AmOrZrmva7eh8olE24O7h1RKJEN7dN7
UXDSeZPBbPck7YgaO5JYB6QQOYdYftw8Ay2AYpsA2rck5sNH/m+38mW0XdjqhVQl
Kghk2KOQTJF9IVhlcscf6xEmm3H5qFaw5cLczMkZc/wFzn9gA02B82OtvdzVSk8W
/OrnChd+tvQFUW+d3dCoDgoCyD7+XHaieLaWjGZQBwj0yE3sotD4VPaZGxAvyBJe
HAVP2JzkePTAqpyusXmfNZeYHO3FhuqpZrWk4s8ZR9nN1zprzgsdIoW9jamyqGvA
3o8nRf3dMtYccGGIPJ77BAgZjJOfodvdMtPAKjfkVH/VGgh6jyo+PQP0V3Mp94OC
rL01GCaVlubA80tpFR3giI3DYs37Cuck94RRLe+CB3I576DhqzmCx655KeH4vFwa
gYkbLEnz7tuJ/2BZ+kS4+o83E4+vpJ+CU3cx2guOhWROpR1N9dQ4nEvw7Q7+6vsV
ltGru9my0874FfjIOlVlktbl75axOuP2ozJNDkNOSGhPh4vcvtxOk3Y0bhV30epX
6oD4gWoBV7TzJUwPtvMRSPKCB/6Vj+u3CfCgpnrQEARElYBGQQk6SrjNH6nZ1m1u
C3qnVhAPrBWfAKgasKfg7pz8a0abAuju+mouyuf/eXo0U+B6y2hochdNFQ3B56eC
LlxHXHgxVOYXymd2YX7x36gxyzzAh9LH/xao0bYClA/QrWlanrn3brFpeIqjLR0A
+nzJkm+etcpGze84kwUItByD8IGeE4EEICyO7hEHSvoPfxSqXiGTL3gaAx7q2bmK
/JkX8fX6sIaaWVXj7/gUEzzq/IW91g6w6WPn7L34/4u5v4q2rBKfzlupZHI+PBSQ
WtvMmRMrnc4d3hpKjWAI8BkUKjQMgQO9VSy8/SZQXcQno70QlorAZTwBJ3lQmWBJ
31i8h33yIVzDDM+RqMxwFXz4f4cqhsdivnjvA0fdkVnWLtexHLzWnh1UzG0JeW0g
7sIFC+2xTi0vAaKXwXRQulZ1uJgOpzN6RWPgAylXjqENzdwuex7lbPhi+DnPp0R6
fe6Vxi6BU5pUJvM3FG5tB8K7uSwbJdwURmyTwZpdh27eSvi3p5ZPkOsUbluodnrP
gTgo7Fv9bqUgHYDtbAHLDQRZQfDZKVGlFLkP8v4THsH6HcDF2l+UdfcCd8yQiJSZ
C/r+CvWoJHSMwWpLl3dlmRy27M3vJVngkLMO9YNAPWUNTeuBA1k59J4/U33fB2sR
r9SJdmzwaUYMMikd5aE4ACEhHIQ/nUoeEi24tmctMp8UrV9HnHxSAdyK0q8RpC34
FDwy0n/YLyS0GzR9oddwCO4KyV1ED7/k45OFL4gkHtWBsdd7VM+7Oufb45WkxQir
/61neFGB7xlMm2oyzUONVRsxpj2TjLNupWJ+8w/L3TF3iXDgbvaOL0OYvcl/Wm67
Wx178DURoS9nDO+UYQO6oF2F8YyNoLv8f0XEbR1YJeu7v5/NhSWaBeaAXRoEtT/2
30Ww6+sS7dWrkWOym1OXTas22KImDGFWAXHMRHurC+luQNE7oxaPYkH3/EfCe7Ll
SWbjZQKtFoZQmpd12XI2Bsuhc+i/fEkZ8CBVQ2xkRikiGrsDbV/sF0ga9e9vT/5w
YUTeV1T/mMkxtbVw//wRJHCT4pn0HcixyQAGcUHJWjDxuI4KGu9UXoAjSKWQnPe0
mAREUVQGidg4ubZ9JGt9eGimIStMCS6QzazolALeYZt/32tXxdSbIswegpJ/2cqB
owEBL/g7M9cUY8CW2ASAOMwBWxLLJYiY275MY9OFbRsTxobTrLG3yVI6mgRaDEJp
9ItmqUGuyj/6Q+rlRY+oH57mwCJv4c0ay5ddtBS/KA8wjzjIwrcWgTNMmyOhpjB6
AQV+1YlZYMNZb0JbcJGSirRKBAtXvkNqDXRhfDGwDlWgJtqULb0LqERBWBuAxzTf
RCKp6F48nif/I1Kulnr40bHhXUX3+RNXGwCO2YdZuOkjjCv1vq7nAnwSPLuM1Dih
ctnNT63HTdMf2ayU+HdWDIsmk02NAntw50CRBiVoMVZNP0S5vwJ6CN7WrfSVwkLx
p/3ozmeRbh0UtiVw41CqP1w+4bzTshJXw52tgcjSy0qFGPCEB2d4ff25Mr97Vynh
sLHT6rbLtGflaoTd7TwnFzzKZlcdOgckgmnZUGGQ4q6d8DUriXSXHsAUxS2vFx/F
TQ6yaRy+l5CVF+HbrgSTvdws4hwZF4mhKyWJF8HzViejSQ0/oJIA5wo9z3tCyJaS
E/sxgECqo18ldCmhv4uNdvnKGjNgzDTsVjp6IYpxNIpa8KDWL+mj5UvW9TPz+d6a
RR7haoclz7S/9L0hL4MqUndWIApt1ouEGYfh28pPB7TLzZB1wouvVaRhcixatWhv
ls/lnSJOQ/EMQ4B8oeSSREr7c0X6qgqB+ZDt+iyct6rgVhH5XxHBJmuw6t5d4bzu
pGay+aOVmi9hZQf66nEUhxhZxHd2l3VYJTY8vPjpyw/j00oW9CglwYOFYpWmBTt1
3qi/y9DzjPG8DMK21DnqSBCFXH8gN2OsgkkKJTVmbCTBhONLW6iwvtZ5P9XObx2c
tKz2rgTJ3rLcGiawY849PIQYBPP6C0giB4k+o/BxzayKmQM3WHduGpud73bIp191
9558cyOoYEID++it4eJbFISnVSAJTk2bJPIrtRJHq3ee/feJ2Xmv+I2Yo/4CsEJv
wsXgrIcCHKIKhlsdUxC9WVP9rDYShDwtDcjJamY0R/5Et1iINzqzEws6yHRO1UAe
0pkqkPHnbbcp7H5pp8oRNZPG8OPHYRcxbMyRZLQt2FWHT6os9h0VFNceta1/WoM1
j3jF19ZuMPAiTf3PqY3k4KIT7CLLlMRUVW+wvcYb93621Ej7Ae6r3XiNTRT+5Gjp
aswAyGFtRmUvjn2NxP09bz04r1AFjWKNg1JPcyrx3ncvggpxdjw+j+CtrIe3M0IM
MXQ/UCT/Ot1HNy8yEecLGTZd6XGhhZ0e7JVr7wTy6DJ5bbFCcxVsIfouQTCrykHG
K4XAlTJd2qKiQsvkVZeRaFao501mxd/bVrR7wzmz+lKE4/x1YxMPqgub7J/m2T+H
nLonaoFMy57HFMvbZep1h60m12ChaUHE7xlZt5HPXCVF+QSL7UxxilFzPvWyv62B
nnPTBgu9yos2jHrlvzcSZQ5Wgw1wkEIS5dKitPGbkz7OQKavpsGN7ZLMR+afkSdn
4AIiA32Evd6n3iP1lWY6RKTILk6LaB53PIj3Fo/J5Kvl3S+PXQvSn2zBIX7/5GHh
xoyUR13XOtxYRb28VoaQE4khG0hC453+g4nkL5BbVKlAoc9yhG3pBIZnrd7Yvxlj
E7WibfhHjc8Scg7F5AeGh497gJkCUfhNkgSCi7NpKfRp0zmcmIVXD4FdRqOgCgjE
PzmDO5rQB1H92JkT+UvLxyX9SlurV0lUwqToF3zS5mCMvwCx89nFibvcSYA2gTzd
ufODrOra4QwhDbu2LWwZXgtIb06rUa6kMjXqHuoR8GKVvrdF7I9+ucwysQd1KOod
52QbqABjxT5iGVsHOVt1SIE+IAzF8/Q62uoSC1lXhhF1ogIOi3+rSw6PNcjMsNb9
YRi5BrtPTsUPdW5Fdsjy9sO0j3IQoOHAGadsFzSqlvKad/QG2cEm3V7laBfPFBmv
VegoDw4JhYD3T24mbu+ln2kcAFhp8iOjHo+8aXt9Yy5hxyMrdhh15r0NRMkN90BN
syFRRiTRp/8L3iXgk+ZzrbPBci3r9IKq4VBxovEEMLg7SaIt1C0T4s7xtepqb8xF
KLi0lxU6oI2t80S0XCIRwFOMVchfUQCLmfht+R0LXERmsy/Knpj/Cwy0Tpi720k7
PLmXUPYOjz6GjHdDDrEDBAEwlarzi1IjivUYmw8nZS2A0Iky61KO/IYB8MEvNQpM
Av7MpC25lu9eiLxXIVg5f/vaytJ93yFPBUlpEb5GobUBgR2A3UMs2/frILak24tk
+4yhZ+jQUJsgn0zdf4nnmNCZBWiRrwDSgp+HSg1BwalDY8R8iOzjhEesiWa4lfOr
AAbKjG7eMqxXVt/QwZv7ScxWHggOKwT+hOUewy5XsKwuOW06z+YYaCCdFR8LJ3BN
9T5AJa6j/zJGhqW1tJbHRtSzChNMgyNR+m6TF9xg7cCFtLvz5JPn9MHbIicfvlMA
kJBXrWzDCKjNsSvUEVr9BytY1lUiJPbXGu2HGxgG07TsGEQ9XQFwqhxte++DjdZd
Plz4AA3kpXBcCgmJohXJgpdgOftWw88fxNRw8Alpf6med0Rq4Dpx0I6NP9Bi4OG3
ChRjeh5FDraFfX3MvyhnTH6Jc9CeUOOYswx1TTugHlvUKssGBOxOselVhlR1yZgB
IMh2shgUW+I9nm2ZpQsb3AkDDP2sJie4im6COaDz+mTw2w0FpPqbfp2SB4hFonaj
YgSeVvUWPZ6wGd/Bl+MUWqsIKXTBRVisGdX9g/dXWMlzIYzFr/9G2Osgg0MIfIMy
ndGhpsmzaVi7QpdElCEQCImmyLAK5GdvgxA/ooMek9TxgHuaJ6M9K33jZC2UhL79
0c+BH7qwBXaTwrMNUYOmxZ6GqOW5/KyKs8fv66EfVa4U2angzNaJiukfraSVX5tc
I9+ABA1ykzjt4RjP2NVYFKvIM5rx8R/lmQv/Qil9LXhFA9sylxkmLpGz7siE5ne/
ITF56YkPVU6Nh+rrZSDCzdgVKPXmcPawn819hjcuZiMDjuxSTIEoVcZV+OBPkVVf
JX7sD+OY1hpU2e53UHyqBXLx/P45UeKMnnfyoUSXimJbZwaOywn1yi+HG1lo3Oul
3jPazwUKJ/lUh4OaI98r0uNnGTGn0nLUkUk6HZ/PEpHjk4r062FjsR5reUWbX6VE
50xOxXUe4h5q94+H8XRpdN4/O3ilfs1sT9XBUlhtFTxkGlN5NMg+prcWekSNE5fE
hVqs6O8HNdUqhjlVbxu4bkwxh1SjrTNq0OCJCOzovSHEuaR5zp2CdQCV2fTdEB2B
xvxs0xqNa8gZs1+yTWkthjESnOy7dJPHdnsldr5iWKI/RqdG4QE8nS+yqvS6SNqc
EaxvP22nWq/4QFKvnLsoCfL7hzvefelbfZw2wkQThr4WQI2RrTwYjKmg34lEmlLR
Ex8lrXoWIb32vJqA1xafFfFiwGIZgkB+nhxaz7iLyVHJ4JE7ZHF8/COQ3+YEored
Zqn3oAAW/QtrH0uou+RZ8E+3OsCq6+nhL+4UYWDgM91sj0KOzEALiI0tukaxVX1u
7LLSLqJmqyD5b3SgvFwbjHDewbJlLcWSCFpiB7P1txxRs/V0ofn8PB8Ufg0wqqFQ
gbjgoasFx95/kghTCY5dEV1hShKdNAL+lLW8pcTdwl5wtcPOr23giJx5azsUHqux
gDB+/vQ4U7l3D0iDvwLmEMXzWZSRQItsy2CRHjxle1O1Jjwd+UKyF58KLX+fvnN8
PDhhnmW6fNXXBIWA8tZguOJZM4RxS22qB1pevUD3AUfnQS3qgJJKlWTHMlwM/onY
X4WVHB/hhzlaLePksJTUMqdx9CEKOFRZnRK30KRZxRnCae0SepLOL7iWeUGOzmo6
UBJtBSDayWLrz1/l6Jx+v11ssNYg6riNifGfhau6A42/owX7yPi2f2yRwvnb9JS+
ghY4Z5eSxcEBJRbyMqnsfK/csA9VEm5t3mPDAOEAr9Mj2pIo73zO6+y+nq1+Np/p
6ng1egEZCzlATcax8f3pqGf1dyyw/SOvyo+HFjgraS53v8EoD1GV8SVs/OLdZdml
kzm1OxanMU6+fnPQvz030GdyhOqj1L7bCiv4AlfhCXgOlATiowrjO6DPw86oldmm
ecIO/EGd1gK+yhjWfMc7opiV5hDcONlkYB/cCHhSPKZtqj52HHwX451ql/ElS0BI
NuvMHFtHizgLQo7hR2GGuoW4iVbQOQNsbRJO+1d/n84g5Nr4ayXzV6hwrZLZJEd6
I31M+v2c+AyVE7zLeANnuMP+BPo/1Yhy05J+ZaV/rT3ZL55VzHhYz4lqaVaTf4pG
mLpOXEhXeS83E2rBs0nMCr3uK3QDUW93+RmuhaM2HgR65FanFA7JNRUXOLnOR5if
snVsew2ysqD3Z4q7A2HxIBp4IvtQE6oU7+/7JG31giSqkm1ut1ZrM1syOYuU5Dm9
0BIf0XujZ8EJm8DtQdjbLQ0YMZVIlfcaevdkigRGbG7XnMZ4cnepSpEXXeOyyt/h
/PSi4x17qSa4vU1gyOSZT8AuTWdEYjL19TdZviNCuKecCC25bydnX0AlvaeWlmGC
w1T7iITOaglNd1hVi+Wd2YzQQES93HQ/pf8d1HIRtNCR+BaCxWvf2d4QJljn1KqE
+M4/tfQ8Ydy1EFSByBxpRkdAZSpYUUUgRSzwOm1GHCkZ2is84SU8gE47KAlrj9aA
djaySjoKPcTV32ajjCxfdSMnkCdlT4Ttd90rwRH00gzct5KCjWAjbqdHSofUVd7e
Wtda3oEoW1hXK89uAVM3iYajFjDgGMtMUU1/LGYP7f6zJSrveFAdcTLuKx+6evgv
C1hqmitBh4dYKmK12bY1EPh8VOgq75obwiDJ/ZXeAAGwa2q001KHxrpGtV81zaK1
xpq1BzjVpWY4STMlagHifHw2/ByAimDSjo+6wzFQ8TcuhjTnju3cnE82Xuig2sjh
rrBbYHUPB6+jYSt8BuWQ9TBTzJ0CYGVbH8QmNixrDEaeN7hTBglzmUiVnHqCA1XO
t9SQmH5rHo1jt5VigkxudbtDmrroFG2uxb8M/2geRC+636RYiIItpMA+8pM98aZ7
UiQVko5SEPvDuUovx0tBcO6D5XewND1XrWod0ufxW9g8+N+DanLu6oGQ1hiIbqJB
doCvt7S0iRofs43lHNZWaasrXFYR73MmyrvkCpTBu5UisjPhUHVH+vT+zJFZtIZF
IRHZ5e05ybLCck3Nes53RECalkp9x2VQc1xhM1+AqZZUJhtGRxz85QPwKGnp1fhE
V0GRmyIyE2DFIaIa/tbF5rfhxd9o5yTs6iGwIvgy5D8ieVA2nQPAhes1wasX29KS
WEZCBhtbYbxVZoryFuLXvho+xZy0BnclcUq16ThF6B7lRSXFyZ1Kg9aWVrtUak04
byJZ0bXvGfyaewjPnP9T55uiRolIK93rH+yoaIfMHZLsMkCM7ManJEyYTxIqcXBQ
aJlRa6kQJIyx+CCdKrZwAkp2jKUslShITRytidcl5YsxCJB5n+UAgXwZH7xSeg6E
HbOOrqRyAlcqL8t4J74t0rwDKu7pjL65y1qXSbT9eKhtuJ844k0LZXLgkqwE3YdR
F2LaVQMQ00bRp2bcrlF+2GIA+dT8XmPFkGS9mRKWreaCjRgNlGvoky95GIlR+Kfp
yLzuqbly2ES0qWpBaia+OVYXYYtdp1y2qvZXDOkbv/hgcB5/bnpo34jc29vkuAq5
Rbi0raG9b1ks1VUTDx/d+Rou5zGCbzftDvt5wEE+uz7yrCAR6hxYsaL2hzZIEArq
dbY+B8tXv0PW4/5dxA2QuG4X5NnsEhX3q1ueRWrPEp965mvscikhmOM5ZFkWQt8Y
9vvchRXQZIlXL+BKNaeQIBnfVe0rBCgYiN83s0JfSTR3Z6wxHMts6EpIaERfCgY0
vRuOxozvsVeNavmdgUdDPJy28KSwlyQFAn3FZy7r6IUknd6klrXgSWZ0WxRZ4Tai
QqrP8lGoVqzgXQU3AdhP5ndwi7Alt6hFXOU0D53lg6lzDPiaM+lwsz9Ut6kD82J0
mrVuRUDFq2endr2DCWLg6yN82GTWoLb+t10e8n4/fcwtT9/6sIPsqi4mwbdMyMtl
+FowwNUSKGgex5g0H0FlI9DxOT1ERj+lMCN/IMDg6dgj1SGZmamexHJE9+6kTkjx
t+Nl+xZq3S+W/yn556f+MHDMgwczrgpDdRh0oKOOqmUwDjM5lJRzg2Rtw2LdDthJ
V+Qfe0rEeJxEKkRrnT1D0oh9XpGogl4I5/GykfVZaYgsnni3d3tPjvsCz4//d4ps
5NR5CFI11tjG9Bl3X1xvX0B2ij5w2AlvGyibm38vbuWNvFI7WaChN1IQY8Hdb7RA
EdA+0brjGjJhi4wpwyIRhAwglvmZE557x6amOLilbCFODvhDXxwmJDp3Q55W0Ba0
VO1uCWgxZdo7zTwtSAfp5glrCu4rSFXkKjXXf6Tarp7wnCC9lMuYCvksV6u/5ToA
NxP0mVhFNkIPVjxPT4iWRfIZ8Y02nWHoJ5P+jlB/AuqwbeSZN1srezWeh7pxTlc7
DZfpKwrhMFKx+UWWWyFuf3OmtJ+5bVowDiqqe3QSfWeOmhtWdmV7tJXfgPguC3Cw
jfYswAhd3pAq7klqqMhlm29eeQJeMwwCm91NZME4zTDImGG/h8rI7EwZZM70702e
bd30V960mjULqk6qd3zCuoxTSaJsU2WIVamsiOB4k1qUhwZrWcu2qXze6KE/y4+g
O0BxPJj70KOxPCf9X7fZNZBANopusqDUs0LEhTbYSG8xKoDW3aMbpEKQgg378apP
F/r1I9fBKrQZjHuGkbExSfZlK+/lEXOSlzJifuN/FnEtQhTXGBFi8SRIrDczM2TS
vfh1rikQTn67mpwOJpLEoaVTDZDmuqOF1yytCfDZi9nujffEraavHqIuSMKwhhNq
AOpMk8qvxzXOmVMXdqxSg/4V+wtmTMjBEOQOzeGRDOND7f7AwzYj8rMw87y8kc4y
g/PlgPaHvfzja7uz8HkVubP83BDlxgseqfmGC86F007w/F/Y9hDzitl47gJFyIMv
vmLigvoK7s7AV5OgElgkK4dXUW/IhFspNR8LCZicsm6B5KW2ppSmTaO4OUamHk+0
8zKYDnB+VMJV5DZtgYEWDcn2+RkSqRuxa7sIInvUxoGYtuuMsABC/j7i8o/EWVtz
XwNoYwHC33FpYmQwSFMBH/XpfV1J17PxQ2gzdn+Zhvf5e/H0aYdQwT3B/1a3ra7M
PhzMnvyNU/yKkiL1CCU/gQZ5nOLn9UVWYEJbZCzrWH3k9xk6EJ4wkT2hYvVYXhp6
RUjC2K213LZUStbHIPHSZM25jfsp/yxHLngDui3s+VXbtkQbok6FEGs5q/2+UJCC
bBzO2uiGYRzDfU/2lGiAaKDhCdlxulJRobqXxahn2QD1x0k+viDqfYm7/N7kn3om
tgZxBcX6ISlO+fHwYRpseaHG1dFA/CLyb+Y8zHNdao76oN5LdSrNGvZXXklCfRci
Sq5Mhk+QftBGGNQiPjnVWKfva5mnwYvoMYFQ12jvXC4OQMuX3/n6HYEtbX/8+q/L
IwOdrNCipYMaFwXRiIvI2NRvK8xkYIe/zAH2ZAdSgWM0EtSXL4D2I2bTwWZ8kvce
toJgmH71QLBBdtZcHCOdumsxj24ei6yk60uKrN5RlIzyt2PYOmZP2Ii3Dh4gT53b
/9/UK1Qqqduq9fqBWvToQMrH4qiWaKR+xfgUbgjauWt2UGUP3b/kbPPi/tAEUIPu
sQJpyGIzT4+jSDWkNN7Gyqunj2wfekxDqPv9TbGnRuABvt5cXTAyncuuQydmMBiV
j/A5ge5uXhQiPmp4jJ1RDxjTzWGc524WaF/8gjfs/OmBt+lr/Xby0q0bMegt8zYx
nLpWRBaExEHTmAwS4c3LspJY8cqYd0+cSXuSHD6jrtAwJkTVq1UC+ZFG5ztDa93U
LULI76aExL3Si8Gr2JqAea1ubvZkiqNOtvd08jNVzYRN+ENlUPUE4P9/8GJKAB8J
uK6r0AAbKN7lWXoAhmhjfXhYuhtvYu5YjuvShwIeIP5Lbp6ehqqzIRs+m+GUKFnp
GfyzrzbGJWIfZYNy5LTcS7//s84qouGDBJgeBNtZ4i4eu+DYe7HB6CH22PY2ygDY
437yaCFJuOwEHKtFk79QuzWGJsvtR8HyQRTzP3uEKo57ViKpIqiYDV/udsO+Lkpx
g/oWPCYFfIYqskdWm2dJ7CmxKknEM6WwxnZwqXveHzJfbrKoHcEfKasIu6/2DkKr
1wfqjGs9BXIcb9BEM9tfPJxgIu0QNTaSHlEWoICAIfAPX9+OcSvsHacRQJ3yvVdZ
8VfhIxJlxcelAQHG38yZmI7/l/Xic+WhN6qUaQJMPvEbfLX1/O5rWrjML/vP8JA9
IONhszovl23jGtBv86m+bDTcALwAdixzlxhw8vBeesZ1/D724A+64hxnASlBGpSO
jCfhGzViRUjGbhrrHZ2/kazAs84uQP/ZDqOIlzmGz8eUGs+1d7WH5CVp9IiVuJLm
m5FnMAhXbW+FH/BjtAmyY6mhVcU3V87qBZhX0vSzraNGoMa7GMxGUNFN6MYXpAgn
mRl/AMHVx54Br1uw+nmDCQX3OGuX91IV8k6SSi9cgn6NcMB0BEJ2xYr5RlHClZnT
8BWnJsK0YaPiaL5RcfB3m3/jZKFVxzzMdubYO4DkqD0qDv61zia0p6QVE5h4zqjD
cZde1MsHmD7pc0WJvjTmFj84rvaStHg1MW9+BIASAU1qac7Z2y/61eRyBMKHzubf
Kbh/YM2jKiruCCRHQ9rBS+N4ShWAso8OHUHqMRMQJdRJC/o691UQHeF821Qub3Ds
Kbpdn5R7C3Tb8R1nufwHzJq3ktcklzxJCRZzzo8ZbKIn5xQqc9SebC7PiU29zYvU
50uoZYOktpZz8C5c3IVNzeazvv06LTymswWZvV0lPejCR/LGAf7BczCrsTm2RlEt
iUiAwuVY4Ow3kU8cbGYLf1EzuMbKOEJ4iitVl1X458K5wgpE4EP7ymWEnwtt6lRC
bHX8KIamCVNTgGxAyYJ/s+KViTbP54xC17cEMEo5uWh8GksO6orsiZZsUSLp2I3h
wZKOS6Q7ukzJaV5VlRczuRdHWAK87gZQ/GiMMzp+OJPGi9Tj+l5+nvxr8/MuFOIY
qzXokmLnvbFcIiEihfj4JqjuYNUaibzCZ7RGCh3UqneJfgh3OASPySyjAfKt/Dao
PRGX7/iwmzY5PsSlCVwJKGjoTlBKKUbx5JTHz+fBVNWah7/4h1KE1mBrwLltKPEG
HquKouHZEiiPlWb8/+ZPek5XVnga3dKTxAe7qGStVfvf683qUZ1EAowv4m23MM4O
AQAz1ThuZ8Nuj4fJde8b6suzK7vqRlzdexmzdkQkd4G9EC1sJRFXNRQX551HIbrk
VYytbuX501bPTYAiAUWYtT9YnoyLZ4HifnB/WSODUBO4lYhif+56F7Ce/vP5MF0+
kBvR8Gw1J+y5QuDfh8LwOd/R7EHh9ckokN1/Nt2KoifjrGUH7rC72OCQO1BFr+8f
jEheCHoG4XLIFnJY+f03Ve3PjAAQxNDVZWCv5Bky9FTvWPM4K0wyttmD3mpBeooQ
jeqHKHVCTj0B6UtwObxhra6SQTLUy/v3ArZiqs8nSiB3DbOUhFe3Vd5KX9D7f2fE
A+OYf1XQocfa7bPuv9sMblNPDJa83bAJ279/znFRpAAbAhQfoGdpDkkhBEWyc34H
Hl6bgsfC3GqiFjBXES20ilAYYOt4hL1i1t+wi5L2/Yo8KZYNZRchqtknmQg2ikau
6mu3y7jsPQGVfVrhzEANSC9BrlkcSkHtCEArFwdLFibAi/J7L9AZYwVTXTIr2j2i
KqzsNcfspbp5fTQQvyOX4QPvVQBlxhMOPo5rdTe6QDxwB/32DGQXE50v0suLzHPh
zjz8z9sRiru4RSkGEdWKZJ0Er8mWw6RrWrxgbFDpQMxOEhP4C+qdSM7hSuVH+RDt
JPWiDtLS9CWhzt0rWuBs6AhhgbhKd4dSmA5u7lHjEUKaT4EsmD6VjvJMC6YP+wbh
Yf0ZjZmW7nlW4YYCNI5mhVGfJRcDTTx9ed8Xs2mlu6jQq8P8CZDMYkQCZnWi34Yl
yUIuMP+bn7E1ZuSERyqwyGH0iWaYubcGd0s/LWm0FLvXVw/PLjq/fVX8/YlBCPCn
C/R5WM9dYqECScpKm7o1AANSFfp8QZQlhB5Faz7qEVCX4uk1ANrPja5wlAlvRaXd
GId+dDziupsd581D2hRDCVhlydbVng2YKD401onxLPhAtMgxxPaqcufirxX70KVk
0IqLn4R2K/Hfk4rNBYfs9x+ranc6Fvhfa+tqcj+Cu3FZ9hzKUpvp13k86XqaFNAK
YcXf7Fh8Z2q/ZmYwg1AnRZfUiiLj5gfkR8sLl2G9Yhvb/cvqfYqC34fWSJUyXZT7
uxCGJEeIeVwv5joWzUogy0vIl+vxwkZzhVpKHg3dk1kFG62JsRTQ1A4a9ZTS7x6h
gIHBRAL1Bnq6tnWrwN3ndfuvw3k79CyKJMWYxCIiTZnvYMF4JaJTgwruP9yRfTkV
75dsYOHQID2aiEa6z1sb/YHEH+PLwsDrJ0M69kizJWDLhfgqPl/jwPRErtfHHP7L
NCO7Yw2fApNNW/HGxmoBBKr3ilyv4W0RGcdBm/hxnMu11jNqIPQCSPjSL5Psyfad
il4n7ddPef8Pg6BWSPu6YXxrnYMzaahKHz8K8UaFH6h/jd6xuzxDz0k0DIk4bnIR
GbHP2Q1ejso+7bWAWzjbYkYsVMc3zW6lx5SeKqezG0PcVZKsAFz3wCK3vt5a6FTT
peqw9dIlCtlyeuIf153vv+5pnozJvFBgL1jnUlAT0MGj+bb0GBVtj0XeVVWLO+rz
E1QV3G5IRJHyxN6gr30hc5+KZj+7L16rr0e1FcmfWs4TS4W7nODlJJF9pN6MRDnR
iXsEX+/SVDRKcX5p6It3yNZYQbUGc3zdFmteoK7HpjRE63j1fiVeCj36IbBPEj0R
vYYP1ZKhtvtu1VObvipeLRtGntKLJWqZ2YytfXTKlNjpB9J8zgJNthn3BS/I1O9H
N1CtNWRQexjSdQOdhA4BSGoD33KuH+VANFgbnevUPdLcaFg4sCokUSzNbX+JmonK
AE0C3m9iHlwna6y7gNgaklEGZ3TgkvucU8EI+G82uUId1Ip902pPlfGWJS70r/eP
NHXO6j1oXoUT4mcDW4Dm1r+5Qwaxq2aif+8E72/h9dbJ5Srcz8zXHiE37+Gr/Czj
yn6aK30dfNf9txx+dvDWGh52U+O0Mwkb6C2wNhjKcHo/HwjGJ3OwUW7iTAl7QXv0
r+MdPyPBqMdDRQo6ljb6KBcPTLn+yeaHt7NAjWGfmldoE725c9gdZSvONbqbwJGj
m8AyTy3Ohj33zw/F726kxm0esKiRgTD4VCTEbIVWwFPB57ld1BDpN78mPL1aQ/Xg
JxfRcn/o7wp2kNha/zTWbBIKIzdvP5ckvcu4ALptDkxWFZ9emAO91Wk7hc6v0Qbe
RNUo/EuSqJrB320MfbgUMqL1xbG332eHETkTiNkTol5hzbuqd1kXEjTWdudw52S8
AZKtzMJjZAXunaUfr9e1jhXDJuK4LoSjLdEBT2bt6AUuCLDDOblT8swdZScUiKAQ
CO/Nps+eg5IcYGn5UnpgehkYdAxydh+2aINltfhN+IV2/lN1WuNZL1pgB/1RGqZg
eMHoJMfJ3IsDHKvgaAUECWob4zmTNklc7Oy4dqTHiXYt4R+LP/P/boT5v63nCwwd
XICH48Td7ew/ztu5KBZT2/p5VeLZiYhn/Ag4i6yDGaFKHQNv11JZ4qbNNP4Cd4jD
+JvpQxLB0kwK4U021ATz+2PRJFZ//NzGa3PkJn7k2RvmfNr9L3Lo65B/zk/+r8Zd
ZJiRVTYXQLTn5WEKO1rqJJrVulTu45sUierJYC04iPQfEAzvyejq+VgO6cn+qw+z
MNkEJ/ArSUluOoau4Lwmicg5g9P8VQRzmwLdJ0/c2Gy5HKLBTnYWoHl8MRLcBV9D
gkxbcye7JW0YA9M8P0PkCNETOSq5DbilFfjwOPJB9rJSaRTWxmQfUqFHuRI+C1mR
NifDZ6jol+joH43qw1xbF+kRps4DuumIBXxKueTZcdU6q+cBWLj1ObJ4rLB4b91b
0Id1VM5EHMUwDeneYuX//d2b+CfmB4fPVgpA43oU/i3vI4UO4OHygIAze9atckwu
ciKyPicnb1lXdgpBq1Iwk52ZZwh/2cpbg5ymd5ESHWslRF7M6gZ8lJ+oOGEEZFrM
TXrDfguMHshzRSIpKLWT+uNutGuegEHxJLNwP02qkjuIg0ufPUZuIWTdQ4eEHxye
rDcblapef1rAbWBwF4mdJJ0o6HJZCypyJvq/ULED6WUMSGEjKNp3BM6pibbh+5oo
jYvxktafaVLh/jIleUGaV2Mdzkg9MyuUdz4nj5nDgGqWA5YXS+aY3rlKXVl0Tr+v
Bwsr0aHyqAb8dFXWz4WruEzrTGHJf5ep1fAXwHOFy1VW+C0GVB1NWWcnVHLbKfIs
2Vx261B/jje+vALJhvfkgvrjuqQSOOhiusJ3qj9UwGTE0dS/mq5krJDB4V82ImqW
/TSufosVRoVyLsBJvLeSuQnmPwwlS4neRXy01RzL2veltkskBqSiVQX+B2fLf9at
3JiuQDMAlzmkZ85TK0cWg4jOITnAr2iXw4lvDuBb5vpQ6/adpPqPEs8q7P3JR8i+
2jS1vgYJU2nz7J97WtTo+JQmCOGBURS08bLH/kLVYEZnweGAi747UwV2HEzNsqwq
tPHctiRaUzCsCMxFq8Omxwh2xDuz9LO55IIr1uT1AA7cAx9sstJSgZZsim4VKrsC
gOOms6ddzGk9q4nuQD+GLUd5JxRZnCMaiQonZOdwiqfulYOtzBqah9sKT1IkOr2L
yjFqYeiLXeec5Er0F3BNgil8JCVKStKfkxVvTovLUAp8puKbVJ4FEUwaLRqiSFVD
tiw3YI/46P2j56C64JC0NzsdI/H23ZpGjLyaRfJP0TdTiXfc5iKYITi/2VBWGM17
GQe5cDaoo1TqYXarb7ZLnRVJ8uXnjPHYqg3jAhmrkAv0e3BtB/f3yc4MaQVFR3+N
1cA9kLLQlWRM13Zef7TR5uIeyuN8EqP0t6X5VnAR5eIxNIRr3QM7MHCI5344tt40
T7tiYXZhzOav5ZmLTCLkz9zoB0TqgQFy/jFUXM23AE4Nw7hUvaQn4ud2ceGVu2Qw
KeSiv4emt7s4eVIn9v6A6Z/cNdxAoWoONq4BHNfUtHYlxvv+y/7TjwMY4SOYJqmy
A7Gw22l59adVmBzPHWuzY2TbLmo8u5Pj0DJXtOaCOnrU3Hq4mFcAflWAAYRj1muc
`protect END_PROTECTED
