`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eFv+yDVxE+N5ok7iuw+qSaInbD7lJQnjTiZN61n6+UgxXj8ZsKNSyWf0K5asYi8L
AebnCUjS25rIovtie+rv8qRH8Uxt6W2bPPWNsYaGs1DK83EuqFyDvfXP2PKDRXhZ
PDQRi7+o9dxKGipV+p/2H3ftPb0ZiMZF535//tQAHJ19Z8OfoGkopHPRAe/C4vMf
UYmgmKThgEELHef0Tbhqvg1CBGmNO/oF60VlmUcJQVL3njllT7Sj7LS4wqttpp2z
FSjC35OJNZ3cRBMyJr82su1WUB3m5QyMWhxGe0oRFRUIlCDBm/FcC7ulO0axS15h
K/WXn96ayNfXwo+52GjEs11eJIS4idwPGoRJRjLKjCOCtiWPy9vv5gQMt81NHTmN
a32dfdoZDQUCiTUbMEAz+LUPv/y9weY9scCQJK/RoBfDKvNwVOUzJAPcuIzjA7Wc
gMc0X9lfXuFLvz3mvRO3u3Bcuhf5g/OyGZ4f4l+/LHm6S/wDYgpHvzW1dsJ//N+F
/rJPQSgVbemjdwYjVEcGlbTMOa8ZERXDfcOWCzLzmREq6wCMapcyuYwD/W0hORSB
AbWP/IQXqDsdh/ZV4Xbk19dxg1/EZ6zBWYwknlEQHHVpHgEnytye4mB7QoaGzJzi
XN3FBtWIxAUQ0r/iFZ0im5UFFPe8hAgGQ8taR7AbvcEwPvUH2xD9xlgtIpG4Q+qj
twFcKs0eTKkLiBx6MnWdhep1fSHYIrCWTn51tUL7+LM=
`protect END_PROTECTED
