`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
AgCUGjhYZOhTDRoKZqBEDhRQz4xHbSsCBHASDQbQ8C3QtxNzI0Zm4Kd7hxkKSQln
omrGGDbB3mij0sUq/tCFvdg5jNCsj2ksBMMkh2hLiyW7Edk4nKd+swJ85x2vlbla
rS/TJQyVjOkP9KbbDxUi/Q9pKyMLHrkS5fqMkmoimiQWN8PPoIh5PtL9SCK2u4BF
ptn6O9HHdxCYsCJbsFCCvHpdqS/pYfzZppwgw6s+4SdHrnRsPxquZmON++ckW8Ku
aiesqcu+o4R5T/y377vfEy+0CYpFC1iKdQtoLazSt7dXOWge5ujHmIWgGsPDxVxp
K6j3MaqdxgZEnwwwW/4e0SQwMv4WseTusEL7e/25u5LGY0i7XShXxMzaOJ9MgBx0
yQLsutPZxOMscV5uQLz+1E0YkV99IjB2KYd0YUSSmyX6qA0oRmu3aMZw6zT729GP
SdAVGEbQQmUTensWNYscY7Ye4iK4aQ7T1ShdkeAXHhTcVM6omsYJYbFxRINUowzF
BaSrn1b3qfBU+Z9/EZgwiT6wt2kpFYBpH44/tVV36eueXE7WAjzS4zgkXQjCgR3b
jHVoZJYJtwoHdyxVJIyiHwxI5X1Yw6SYrUJ3oNRl/o0pZ9MTlhGXS3/Za6TfgyGC
pQPqv7hUpfNzGmbbX6giCJ9VRcRsYhm5jx52fxq8hGuITX8cMdTJIzpc6bmKuNCs
PStSDCBPLGpnIfCMYPEoxSZ8GBzo3PYXQDRSXcH/J4MEoEyPOSsDZ4aXIziBwR9S
WnKk1/XiPqmdGeSwNIAeyQecJwxDpVsOBZ4g415rAqvXEDr3nCgWJa97He2Y9bdI
6uHUCh5+OU4XWOwis5WYTh3ZO34CNjD5LSJid+XilpzTYG45a/btHmrAbyXaHys4
gU3EKilTq3tNDaYw3i3fpW03Ku7/ln+Orl1MSKZ0xCzj0kcFv6MpFARsa53K+1eM
hLBEUnGitaB8RryGkzfGUA6tvTjNRrowQs6fLafZmXW8Yh+VsVXtUSU6iKfg1bRk
Dl0iiDRyOlJ8qZZNN7cWBqmjS3vESHU6/t6ktwedk2PV+IZN7Q1DQuOhWKiS6KZZ
IhvTWzyY0n14n8ZYSAsbfRIK6f2j9EVk6CCShOYIE61RNVnvnSucVW9fSzv5+ZwD
QdVkYRDVuAr+YZ6L4tpE1gARhyrMWgdjasav7dRt2MkhUXIW5RsDdmSf0BdgLGkA
8sGhxdNZUnwQ9RfXRbWiTLmtm2W3OYHpQfpPjl+28rbOauOrjUS6It2T15ZAyvG8
agcKKF1+1inbG/8JDpTQrOSK64pHXYz6Sr/h3zBJ5rjAmRdWID4NlMVO+KQ/muUj
k5GhX1dtM0pI/Kbd2yOxQsbEVTD7ng3bYQQJ3+dyZ090LHVaR9KsE8TFVVmYi90k
HJBsLmbh/V7lJ652PmZXrngZtnyLLj0Kr9wmzzA1672S5wf9idP29smAyOhN+88o
M4UOu9JEvrCJ4ybenXSIA/KA+qpml0cCxsLGH0NXsVkHxh3dqYGWPlAh4sFDVIgy
r137hmF+3NgI6ncqEGyV9w==
`protect END_PROTECTED
