`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IUxQa6RmIPcaCJd63G9Nvs7pFSMgevNgnL2veklyO1zUUgtUjqZQgJJZoXaOclb9
ECQf8kx0MS0uDPNOt+U8UEWNpjDc5x25vbZtVpnRlJZH8PBX6n9sbF7UY7dDbckS
h+HoPaZdD2T8X4veSM6yan5csG8Tb8NFQNnTAQy6XUzWrXz+K0ln8hGYJJk3+lf/
zeZM6hbFvS83EwDnR0Dv4NCqGuhcVOLQtEaJbM5CbPuRwfwnJgvZEYDAI5DKQJoP
WubhePADkShsRDOyfCi107McOGo1MgGLFGgyCLYVwYx1qe0oSo8NRfbp9iVWt/sr
BDmYVYagBur6cbmJt1QVhreWNReyRb1S0OCnKdcpDWQZ16RQvBmJROFybI82NmCw
tpKs3SmY3RdiY6dqzjgyrw/Kvj90uN1GgP+IPMl8himrEkPgmrb3fk0q8RMUPqqa
ghkRnng0aTdwSqp46VThiopsmlPelCsjZ31vdP9VBDatGvC0nK2jobtOY1GnZEZa
oM3JDfVetnQreOl8GaPua+oljkV5c6uwFneAylMdHexeuCx3jQ7Evf+4z/mzvdqY
EyZrH5xu7F/NMmLUYXyE4PfR2koqQHVUgDg+Tzkkq/qeDlLU72x71mze/BEaNt1q
TyDvDmksuoxA4DF8BsAN0keoPx5IxEx3NDn4iWC3mSvC6CXF/gXfk2MgSzV1fMlL
qAYQZynGULKS9byoqczB7nitmCx2xbLtJc8PIjQdB1HYFYFWtB6RghHyF/cVDF8H
U6iV7n9p8c19dwhHvCf9CVx5kQah4HEl5QXOIKiqhYKZqXAPt1qbtUjLd3Ye6dD3
+8+oc/KoG8MUdEhQiMzUCvgttW1reUQB6UhGOxY9suGjZs+XOpZKBgTHn3VLtCk0
H5CSC3oMGiDswpIawq33Q+Q+rniR26K684enolere6DVXMF8QdlUoJvBdc/Ag/cF
fWKx3C+6+fYm1zI7zx3Pa6tpPGflaldLat3A9r5Jqv/eYCDResNMtBsNZq2ZhNYg
u5xpz5PBI3CO+fBdzj2IAeWWgnEK+Y15lAyMiq26nEiJVubfX2yqi5P2gskhz2Fn
z0z1QkKtwD2AILMkIPTHIeAhxNlFjNGVo7hAM2Tl6ouwIbpy1lUZtBGLhwi6xnDX
yIoq5VYRSQBtb1iwgI+TgJ/BBsx1schi+Xrwr3qzh7UjlF4EEKF8914NDRRgihDI
DW5ZSJ5GkUCsN+YQlwMchI2vuL8nAimi4wpNnJiNodGQZyO8ix5tAo2iwZbLQeUT
5zk2ivg9+ZjQNSQlDP+J9EsFL+Al3GdshSF++Fn/BroXCxI91SWGDEx/9NoqsMHu
opEry7328oR8iuUBUgzJatR3WqC4ZicVKoX+X7VXhWbmxkMZtYPhXhc0mwqXuAFu
80B4er1jbmUVfJpKHAt/+CBq8kh+JZLoiUs2Uey+6cKlCAcHoZ0YbEOl3hpk3x6D
ZtgHMzNHAnjNXzAFMht8j4CuC4PhCU8jRHtKmqGulFfjPrD3xZ7Yp+i88jH7e39y
R47m/LI+oULE7Wl2oDeMfAbNKSW5Q+BchNswxqE8TCqcudoAkD6z8QUePOe5DjKI
aPBTP4RmpUH910YUy6+/kexo2s58hIjM3WbFhOZFsxxH/dKEpBoYlHPbz4qDma1c
OyjUqlsN98JTw8oEBPk9pF/u3NHTa82HjrRpeI3qOd81a90e/R76LDyc8KLUMpSn
/DfET6nEVSpmWtHF5oTB5V8VOCLLeKNhCLDvX9aMqDyWTgyCKCKXulLiYUoGfIgp
ldu1umKZ3APY9RwkEGO8c3ox9pAuTcCQNlQXCJokLSdAGx93vZU802RHUz5txbCc
gMcRqGu54SsU4zw7YeAKT+y4Osz74StAf9+NXWNEdrAfAynRJDCvQUiybmR36kqT
pnb0GSZwnHbx726wFNG9tvxEkst7T+m+s3XTzl2FN5Nmp+fpPT/Oy2YQcjK+LJvo
cu3aw5tNFnsvO/kL05TTuF2kcMdxJz/fZ2Io3Cgf2RHXxVOH7mCInsymXJEaeb8x
bsuWh7YrVq0DqkeNcNw6xkrA0JxeQu+VhN3MidPNfbV2iBRJaQnJPpPheTjjlHdD
+TT8XSuS3btZoQTnw1HT8ICArOOuQfNG8VhEckiVQ2hn2qBTNhxsVu5HPejc31FO
fe4zO9v/tY4IzQXzDBuQbI6I4KOQcxwC9/hi69umBbM=
`protect END_PROTECTED
