`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
5mId+pgkxUs1xQZWMQk3frOU2Xtg4kKY0y/DbTFmgwUeO51PLB00J0y4+PQ7E2XP
2JobnTPgkQRWuDUgzdIOmW2VHLgwCRT9z+2ghW4VNJiEbRew80VkcEXJsgrmRI+H
J2+QAnO2794aCKiiXSma+6FvwGtNLCBxD0vaD3n3UUpLVnLRaHFOd4jrl49Q1SrS
2SUUDcM8Y/1errK5HUmxiIVaqqUok6v3xJJCdrBgHO9OYYXZA6AdCNvmwhbGO+gn
apZcZR9iwNywkbIB2WA/PNW/td2rtysSDi+C4Me7kCxNlaJbwamYxh2w+9VKgPFb
kKRBSEpC2sJq7XwkLunXbNXMiRCi61+bwvof9TzyssJYCI7eIlgcdKQ8Kdeiq8or
SiGenggmI8opzXKTgkQMz4wirw3F7qtKZivF6bQvl87Gvp561dJMadkO68Y+JAhv
yGuxWPJxEJwhpogbcZ+Ofj66r4s0anARxdGO0CrhJ6TbHL2Qqx+7MmCCv+3Zv15f
U2A1Q7VOQAZkJ539PuYzWkAPs3t1k8kcM6T6jBGyNgPv62/ybfVU5fmq4USc0aRd
i1tnP1J9q8ATHCn9pWvUvle5GZWVLpQnRDi9LQlvBMeFtJt2RPIYSMUauX0gY8nm
1vn/C+4Rvd3/Ku+yPIlcN/JnvuyjYE2NmJWqg+zS/5dLIw8lBUgGJ5+80N+3S0MJ
3PxpeItUnaYIE67EH8ec/FjXgeVRkKCuMLeu5NoMY4KQ3wIHCqfhqroIEsish7Mp
yFfFdwyQCCMFKPWGOOKrfMV5ToVnhIGK3XBXrsS7gRyPzq9brC6apUVY62xAcPDz
6xFds/LcZiqR3uxmhXy3ep7jUxy8ypQIIhZUG1CCKQer7vyXz78deGka71FQgGtK
mwboSWsa7Nc4SUP22mTh/BBqAyWJ2KVAqiAl2IF7Uy0vCZiHFNtBXNRKWG3vMhJC
4tdfli65PFZl1KHbdYsC3AfrQNbcVUM3SevmTwmVZ5L0fWkgIKHiQK5waUTHmgTN
8TklQjmjvesMBO7COYUtKCfZosvMcmW4vBErNW7PkLHrnX1ykx+pkrJ1orUb4VD3
/CwACR4uLuqOubkH/8203q6Ts9FJfOfkdrivMANYUOmfSiWLjvvRNClxfkC7Fni3
U4hPTAh57QGOKe/sXdjz+kV8v5RVY7eQML/RaS3J847r3XCOVLA81ZD00OEZW8TC
St6RnKMcQxSAEYZ/XgIiw/zXTvB8RJMZt+LRi9T9FaqOy6tcWVMuDZ+3Rha5+Nb2
QxmRrZ+eS/ttCguN7rqZCoQOhQ891GtFaqpwpS7ik/nqknHHF2pWSIKpSEO/EF/A
2Bre+zbYNc25yE9Ffr/L2uwN7xWzQW1a/9yqAOy1ji+YZ/FHQUiq+rbZrLO7e19o
WcQGdG8gIVRmjjQims8ZhsFma/GAy6mQt+PHzdEjWJ4b+ALQSXNUAmqkKRSuF7N5
cGeuAO/KF5eUp8Pq3+PJROm8tIroyD7LeUApk6ddQUcqgC3ZiTnmktzxsVZSC0/p
SQ3MM4mQDxkJZ2OJbm/EBCWuDSacEjENzv7IlfcdeCRdz9rFJZweY9X38dTgpWYd
C0hdoecrzf6uofpxhOwb+Yz6MhVMTGaSLrNUGIxKROOa+kZ/qDmImRzIV6rqu3Q4
IwSdXBE6oOBGWr7dZI9MrJQndfwjdp3h202IFxJ/mbkEicNlK3YkZpFilWqSR/dB
+V9DvPSL+gGhIGQYyUgZphVWsFCEBQQLfjQ/p1g6EEpRbRxvHbuMiRnUCJmRDW/I
05n0fCf8QUJ88jojYKmO/H/3OTh/5/rwPRfh/KAZhQ75OJWrL1nu+qvmJfWY0dWM
EPcHScLanWbd6M/sG0QrvDrKBQDYjE9IAUj6NZBbJIzi7Qk/yMM0WyFJvs0A1S4X
bYy2RuogWm9y6jdTG7R2JLliPuT869dBv8ovM/ZcJrsV7J+0Mqpip1NPW7ysCY7o
F7F8ZT8QNRNdhil2m1vsRoxzOrIzYTCVzFJLpu1PPcpmNqkXjiPZWE8PfFRYdCBQ
jlMbddtc9su0vNh2mECtC1mODNpWN9rHsYzU+iGM/Alfg8naxBLz4XGHD9PT0xnH
xyYGcXwc5UIEiriKsBVZobS7PjRpMk+nnBUCgRggI6grKtNzz2htK3zTiNgSD1/9
2h4dvDbLqVX8GPGvEvAJAtr0MxtQVT/+dbwRzzdL3AxtH7SrfTgLlcNmpWkyzy5h
xZWfT5pohCf9s9uNrEeXsfCwBp+rB/9ULzVjftLMd9dkbiapy2lR0m+Y+6mdsog+
CWFUZC1jalUKLCVkxdHmUarTvYZNspd35vPOQI5L5xJB/Q/YtRvP7JTRxv14s93O
O86YtS97Yas8QL8Bd6eDJhAR8oDU29QD04SCeHbJ4Qop2Y5EFYtNDLRMBkLw4rNM
4/eFiY+8FROstZwyZQz9Otb0d74DJC2o20kiEFWepMBt/B7vxYn9tdaaue73pdmD
Q4bg1sVFJGoBcgmvGp5frGVFHDYav1nri7e6k56lSD3+lccWWhv5o6Cxhk6mIt5R
IicMXiBjY7qQ1rCz7o/d1PC8ZT4YLkF6DMneGbfAe7FuQncev0NUYiI0FbBln7Ob
EMUsJrOfSQjXxKpvCSR5tKscnF466izQ22Q4kuVQ8zCy7Fuj9UI8z1vWsDw+21dE
8k8KLPzEiosjgSGPfc0E7bYPLaFxDpLB/dtwh5Q48K9s3BLMAsmHW9NrVRsvmkd9
YsffGqhy/uipl8QxEWVYhgYJmehNWqzer/V6Lkz0sTUucvBBChXkZhPGlYNcnCgz
ruaOGQ0k2xe27kGAP5wZXuTKneuhrhpUPKnLLzuol/MRyacpC8pYsykt9cImeqFX
WB5cR6oKngef7HZ3WEBfM8HDNjVL6/J4BO5OmF3YiEfsHgWHrcs4UyQHrnGKo5/B
K6gkrIV1/PBypEAkmCNkWYR3xDu6uhMXu5Z9p4CBmvzlrJUUkAtjowJXQAQk+HV9
Jt9yKuJb+OrcSyv/QH4/U7KNVT0337Wac0GTXOAex1wwFIyewOetQFCDcOVkqUS2
QZglhcH8sinGSuGEkg+6j28PNYTkhyiv/ElztGZDT20YT0Z+1XqOAqxTFprxiLOL
DbcbMYmuDEz0fTgPlWyzk0toBUKk9UDFUW9T4QXQf86LiEaDdy5hmFr2QYIvHKYg
OcC60QfBpiFPtQVN6W+PSLUDTkh8Vi1otAbxW8WF1kzjkI4J6JLe55Mviu2dDL4n
96xxAxbX82lHhmgXrhhnikLCSwxHJCZ3V0QsaacvGbaCidkX8mpoJ6fQ6MTi8AoW
EuvWbWJA6drTvrHRNhGBJnsb+3Tc5dMxJN/mNrAZ3LOYLh78sJupiQIue05kbO46
N2SVayDmneL2dq9jco1s6k0beCj8XcGkvgbPNcTj5R3MyhbBZV1jPC9g11o4bMkm
sEqpznvCpUnr6RthEDAe0Bzco8p6A1hknC6TTM/3f7T4TwQNYNU0b8s/mbEZ3l8q
FJIMsBgyQ8gDv+u4AYrBh6libiXnoUMH3SeeHGvrlqUR7R2tbJYL9xTXBQ2oodws
V4dNKjI9ZQS/RYaDfV8rRdr+3t040B2RkT6LD+nt6f2/c16nBdKoS5ar23yKpPL6
DDGHMT/3PNVb90P447A/zFDVWv8QA3tvCOUyi0kI0Ed/weezeAPqXgrPpGTV+cwK
k8tJZU0/eSAa+e8ehDe2oh8bZ2bR3MnpLndBVXa539Rvu39TcJWccALjduVEjwKj
TqSg+yzr91grb0V6WvP9n+9BpxZtniSUbQuaMkQ/QJnU0c3FWkArNx68d4w1U+Da
5Rm/6wQ7A2j+qpPQbxulIoxPKuyBc1tVBxZPidGhvI+gIPXRnTsQFOwlbFEw0Fwp
FT0ehxdMjxOApoDxXXYObC9UgYRa691ZpkzybFdUqqdOVoQrZCKZHD7ROleJRejb
HXECGqAdTga/Tl2Nh6+IskUdFMCLVrWRL8MO8D3qSituMR+hM2lI5zK+qZGfs+0R
rmKPuOzpDqMIrFzucqhPcFEzpzyVRYNYpWdSS94LMJOoGBrN8cvrzvxTXFaeMfZq
en40KNtPQGd3VAs3y4a7a30bhlG6+N10WtWJ81kN3L7QxFTkPigX1pNv6EfqL2rA
dPomeJJrOm8A8iPASznsHVO7q1obhH6cT/FA3vj9xcKWgMT5qeL5BNCgDSYj11Zb
yLssvE9niD7VRlQJP0jLrleeAGQKHlJIggO5OxM2PGWJTPCPACHixOg4TRtm2pbk
OJOVb+/gcktDUIZoSbMBJewLkge73QtPmo02lwqvEdZqvSEp9AW0yBmpxkCK+K7/
DaObkVLoW0NN35N7ujSWU7Tn+AI1mB9ypT2navCth7vvrHITFT/WDiTw2YlbUw0u
BjnZp8Axg+vcfndqERCf2MgWKkV2vLLiXKYO4JN6aSFXm/5yXxUzAPZ7DNWaGvK+
EUl/jq3EZLXoTWzErDLVUjn+icVZSVA4S9j8MVrEtN0+QXWlatgatXTpdgac5nay
0/ZMrqFcRyOVegC9+JrvRNEOdBxSI2F/2Zv0jgWG9kD7J8F908fCCI+uLInecSal
8qYpC8KuTnfFBi6umW2guTWCR+xRxFP5Z8d/+sD8MP9kunVWPvgDLKxZAESmvxuV
pn4hwBPV+jHGLGgw+C0+qeWLBK/Ata+0JwSxCaH0EtrF4rme+6Rf6XCccLub9+Qo
+nYvwBfg4NQjIrVyWjG58ktt54VfqJehAHzO/Utw24WszKH1qcVbLWGBm2Caz8d2
aMLQhIrw5jsPZme3homCP6YiV3IcJG24LYnH1Kv+BOXCDjjUoue4NyTsqmQ1mNvp
yGSvjYgL7IKc9q1n1doH783JVXUXfQd31vCaDUffVEtg4GLY4Jxxrhr8u/J5rH/t
P7EWVRLffyB+yl19J6D9edwKmrvlLINc+2PwzNRIGGvGbVaMTVRCRrF+JOWQopTp
iiw3UI8zePM9pP0S7C7ujVd1uEXAo0VSBZghqWbvyQpAMp2PqVFum42tRMptf8t4
JkimxCuHgAoa1ErR9RiPuYWilcgSFHfvOPcNDV9Rfz+kWVKIbY+dzMp7gWJiYpNW
C4hofikcUt5HbQREFToGXSvTk4GMkui9Od/bdyvWZ/I26rwclxa0byQRB7HNrO/h
mBdcA+vGaBsnz+cEwK9bwZcvAfx8h4ZjeQAW5qiWesJ3QbRXThHu8Iou27DsYiPR
nz55i5uyqLJM4pNIBYdML4s7zp3EPqRXK5G4ECrjg3YtgGVUWM+MHHjmY++kiexq
SZOhtd+TzwpYIdcLb90X1phx6sud3nfy810OvNo+d2opJ/n8YhrnS9N1og7G4l8t
BbvwKybeQ4GFq7fo6S81vAlMTuZ2ikOvL1B+PuzvQOpj6F8OdkFqEJQp4DGKsYet
3xoZJUniPDJikJScdQstJ9pZqrP4lMsCvS2+yyphjhOYYwlfPs3zIqPSTdNrozeW
Z7ulifqV41Ft4yFkra6mQGP3ViNwxvI/04wM/RHT+Uy1hn6u0hOTKDwGsFffhW0Z
tZbOjKiQY0hJiRgf68wBjwY7r9SSP7iwOI9Q38U09GjlYBEJwMnJJ9RrRpCAljKQ
bZxdh3/+T2+emckUxQ7lcQytN3ZnbKmqrKfMznsrgbwSZaNB/eDpCWL6/Mz7WY5X
Rknt2zqNXIkIHT7pDcmrM1G5p62z53V8Hl75QN40rbvmKGV5ItpTqfqoLkqRZhrl
vdCr5rlHvsd1VfEw8l0E7Ld4x+f3gGmyauIHxJnh82ObiZffKnmI2jIrPQ3loNq1
uBMrpmMSsh0sCGYJ6X+p/GMLlmQRtuOJK/3TMyrXnuM8LCv/MpJadnqVSflBSIjH
1dCR/Q67uKkFIWvjW+MUz9PSfKRJxYBfHMtdT3A8FyXcMjT5KEZ1rnYi7vn5EBL5
7VyGZBJ7R4WMljb5ruGAU4BUzSBlICLZMDysZ2cOVn7DB9yFX5uoBapHXpuvN6qQ
veHhCQlIHTJOxaGWyf8EWS++xpkF0juhA4KnOMbkraYouuLXpSW2IBZ/16G02RXV
0FfAfOutddXKvnx5D82gzvxob9dQCc5lvdR52HSm16ho6doU8woDUgodF2EQV/hc
NnmeNNUJJAw3gTfrAJDclQ/eWrnZvRflOem06y1s2UPGQOz1Dx6ZUtz6hnv8auYS
JaPT4h0W7BoZRN6TOCUTKwBn+yXEQHZ+ZG4kG0wQUeldTyTe2Ts/QEJ4R8KaQajk
i4RB72AtMJqIq8GKhdLBv0AE3Jdg1EN4SGTi7hbHjTXLx/FzgBsjqrixOFI/c++Y
JlbhWNqmCWkjs8NvEVjLgdQd2nE3731QyGqcbh936Kj7st9SZ0Px3vBg/gZD/iLr
SZCtseSXghtzTj44uphDqSb08z0t0pU1FLbNaRds/+V+RVsbXv6Q+R5Nes8YFBBe
GoyHujEga4jHece4E7lL4WKQ3iGVIB6gLsZTm2kZo/XCo/YV6TqoLaM5cHVxGlF4
agM0wnqHlgfuiV33/FdS7wub/tMyF2xKTlBwYTr11I6CYK0325HDD2JPQKvF5EPj
jOM5WLDXyHo8QyGkoqb/nCAp5UbMZxydbELmMolnc5gUz0oCRMcxvGQvacAI9Nwj
BC2eHj4kAJbtFzuUNC0c6jVGjviP+aMjTeqMI0xO/ZFr2g+T2qSLrgR8GxhE6gAu
+akbjxYVzoKG4vUvoAX4X5UUZjAJH8VP57fgN2C66aVEGYivGVIR/kF1du5geYxB
Z8j1rcQLEoGc1zg18kXPqQHZuS+kk1BhbTlsUwJJPIqUbAc9TbvBTUP+K2/uQyoc
0DvY7caYSegWbocRbdTIsZlGtEosRPpxoSkhKEGodWL8xfqzFv6w5XW9ls4fTWGc
RHr63toFxsyn7glpa24u60vRd1vdEylFZc8NSsGm8vwX/MsIr0T+oLd6ymKGEKSh
yn3Z3bPA5HgybTC+pziEgRknLpYXCyvU6Ztd/ZYsohR9YiCO+MTUp3t3i4HEoAHq
miqGXeZLEjXY6hL0rriUs3ZkViwxPD/Q9J7rF9YzCFUM4BKSy2ZC6Fb2oeRSolmZ
vjxTNDKvUW5zAt5b9tQd629b4R5wbXceKj4vhI8CXeQFbv8iJYfkEjRYSWR5VvkA
wGf5Zfn/lJnPFKz7dlgW6R42C13peCn5LASvqdnme6hWxTyrdVwDotENln5PW5Jv
/cr3JtbMKYhN79exQwWOiih3IqJzXVGc8ZFZJWYEzU/TTn2icpM04uNNIrz6ZAvn
zvCK6nU5upxsZYNV3ELITSZxjDWf9pNeqhkMebhgb3PAc8hAvy7dwdeD1hwZomEv
93QLBgKTeJV3QTHqYHVaZfxYnvcyIckYzuM8fa1McYqO5D0fAfMBeIvpcHCFRKHQ
akhTgoChokcqo1xU5jQVmZaktvph9nDmhLJPifoy0OZoOUXgbrXLllg4hOmuZ/jP
/lTto1EJwVsHXuem4Oa+eE1xesvSGPaFZCA54n6dlLabW8sTJJqIPKkKrG/0fKNh
BQ1Jutt4bZlURSpy7uhdWGJmn3ZbYFRhp+7yPyWGndpGsSr+GovgOcjA96f6YkTB
7twRSE+qbVx8OIKb0frLCegfvmFWdwTfKAjnXTSfq3dJIM19JzMEq+2Djh/uoeEt
yBG87KUOLq25B8HmmkstyJCNdnu/kF2UEyRmwk+OiZx3UcsnguOcx12DGvnmDXFx
qgheiMu44TxEResxeBXj5BgICmd/H6U9ZhsLXXBcfETHAtRfdWABaIbCft3L3tb3
1UYaWm2+Ms1m1uRaNXDb63EZUJVcr8D/WMxKEASnNqgrKDsRhQ7LrcpPnaqlVUTO
yCuHLbw9s/c4eJ9BIPjyoPFWkBeZo7GwHDtLMMh4xVhKVm7Ay5uSLzTPixbnU1Kq
UjYW2jOk/yCca4XgVjgaJjPHEliE3k4JcZnOToQkuekwKdZLqdvEt1tldRSZh+a5
YKpzICu1Gjl1/wZ1ATcnhO1saDo9vTyACn/+TZvaOX2SOQKNbbKdeW+k6gsTfZS6
yRw6VlJVu1uqUWqW3IZQstUWP53d56RbZUhout2soABr8bErR3rl29JkmCYRnHlV
qaeVmUjYabFOdtIKvRemYmXJbKyERt7iMMBw9HlwN0wlk5Sl69/DyZS957/upGsH
aYu0ymW8pabFVJc5DX9+10Tk64XG/M6StSRQacQkm8YiFXSFU6jx0/r4+GUkbdQP
GhCJon/d/kDLQZQWxcwB7H5H2S38uXYFjPLfzX2b2jX0xs5kX40a7WOmK3Q6pb6M
KUuWW8xQfjn0hIztrYO7kjoKrLD1NT+ahfa/aS+Skoqy/4BcJ/FmRg/m7L1m2Dhy
xdeg2/gVfr1dkdi/ETsrSlw092kA6YJ2BZDo/Vj/5iXNMRl/ay05kyzZaYaUOtsD
hpcebpYEmbw6qSlSY0hmm3C8YelL5oMNN8zN4GI73qv6UIepz27vLTLn/tUonq5M
ai7YmZhC94oLWK9xBbtskM/8Ez2FJFKC0bbbrNnDauQimqYQYFMINnBgv9rl6B2E
qbaTDkpqwv9nbLt3puZyRbksnYSKpTDI3jVeOZBXAs/g3uYAXJ9yosfvStd5V9/e
Efs4e4p2ldQe7fcVS40JIjGQboKz8EildfwrVTQKPZ172SSOqDaW67fO9Is3BwcA
X8jcl2neBqLr0bbWI+jU5Gfwb7iJLvbQxaCTV5//oFXKnO7upUV5/H4Ajpf98BoR
RU0lzob8uruG89g1MhtJO57UNUX1ldGklx28S1BnPo4dctzQcOfV8G59TTrxibSj
EMrXnfN+KSuJia4RH0RIUUFIPvAcktxd943MZpRmtAgdp1+1xzJfg+8YB/T4iqzK
x8ip42s1u5Fv3Jz4/lfzHcQqAskOu66Quo8iIUyFjpvzid4LZytQskRjMw2KQiRH
TTA9ImNI6K2z3u1vy3dD6oOw0OigOgxqQpSoOPWS7poQulH5hHzaDFJw4rirKBqB
8JYmNRoDCpOnU7FYXxgpKd2afrJgCjd/5up/3KvQnhp6XA9FPj3kbsLiuqxqftxE
SN11i4PnBt+IurPdhnMWl6jR1EcI3GunbiN6qKvVW1xcXzM7fDghQbLRDTjR8xak
tT+olxbgzqqXM5sQpSBuyWUBenDpe1v1CdAhSHzKJ0Wc0LyZYyAGdLwMVW/0JzoY
f+GSvwThPhCVaWdK84Dhidw6WoDEsDUFzyMtQedZQnx6V51yBXRz8QE++lUAbxPe
P+7fbfMUNy3RXtFIfM1UmnjqPTYc2sd+4DxffMeg77yFCuNLwSvZD80hvfL70Fub
R5ly1DeqoVRfSudANnjRtPmwfXBPxAThnaAxdLenPXSWuOBOmE1LElNItJGHXVjg
BO5VKCcTrPYGw+eytJzpZKEUUJeBkVwIbBarA5o9cHMShhIkvCZaI3qoupADdTPp
V7fwG6grBwARjRItScltXjpjtlCH8GomDVMGlNzeATTmqP+Qf7ueWuDs1Q+hWG/e
zqYfTV3qEPW66tTZOUbono3N5yOrbQbSWAJNl3JXk+BQvaW/4n6BDOutlJRoReXo
gYvkwxEbDnawgjCMjKu3TUIVyvcbHr3YzNpeQErSTeApWh8X2eB7wmj54wFbqrUM
r6+fJ7ATKSa69v7Lrv36kgMOUZNR6xbtUzToY9pgVaE/yF1tXOIl3dygwv5+3nv6
JcmC0TDDEdhRd3ryFmUgbf94ixRwBVMESvy7GxraqBjIDJJkPUtbn11eRHPEGiiT
bYyaXcN+zNijEagPgm3O6k6S86luCx4UPBB2Rm5b+lk6/6xlI7dPvo6uDPuwD5tA
D61aoNqlu0Qnw3gejgnP4bjh+xAEw2fa/tCJ9aK+3fJ6jHAfutjsfq/UBuXtkk11
MXsS0iserf/egeEELX1VlbDNXAsnpiN/LXQ0pO33BCNOCXJfMU5dw7OksixEQKtV
4vyaFJ4WJy02Zbu6XeNnf4odJ7B7ay34FbdP99WbOmGetXHE3EmCSfPR0xAV2QlE
MHLmS4Z67wes5/pG0RD6bUYUB9Z1fJBVF9/fC4xuAH8i1GKsLRAxkJDSMCrOq59E
7YEgOc30MXxcUVER56/76s7/R6LP9hsZ3h3NthBl2kopwn+H4PTYftOPAePTgRp3
9GaJMxINp9I7IPeY8jB5uMiclqbMeTdKXI5uCwCC4Zs3AUIgtLV48EX1qh1BvAQm
l6VjP8jMAX8wglqFD3c8LlfGYAfl32lWuOOptykJhZRhmGbmRSC7O2Gz29kVYc6M
4OC6PVBkgVQ1jvUqCqoRwLi8RsqrQs8IFCtMazaoRZW+zfevZdhW7MX1k/nu4lIQ
AZX6NJ8UZ3m+kFUOFlPRD6tOPOCCMr+A8FVH9XhwO6Pg1ZOtq1BXk/xU8dl5FkT9
drxgKPQ41I26ra8RyLUESxO7D1M5NHrCEmoNa4FSfbsUaVUTh78SkhKN8KU8gguF
rhYSNaN/JhICET3+yK5qTrhR6ggUYRUDZcUVIDtP92lSaMZ5+6I6Yux0C3z/vOfM
E3gkbZUyuB0Ym36ECr82rx+Ev/HINbKTfAzajHCGhmS/4CchsPDgMJnwyJRW3OOk
SgIpw/rwBcCgTdQ6H1VHJy2FxdML1Qx19V/9MtV3cS3p/uObYiAzQBCKGEhQgEYr
G/0AsQWmFhBWs32Da4ltFQ8qPGZMsVRt5xn4C9R+6Nrr+oDwJv0EoR3hEpJfDTOK
DMcjiA/BC2UmWs0lcyesj8lW2QD3qd5x1xbwzH8NiGCAusd/pACww/if7Q33zTVv
QlGBhHw57BN/So5wa9KlPfKx6VTjUZTAQUZGCSqqfX+6OEToptekR+6WeMisE9K6
ca+DttozPXpehzoie40h3rOxo5nOasE78jVZkNcOdtjnnM/nHWQiw87YJcGvC34G
D4NhD3Ntk67fsV1GZrfb4xL2M3Z8qXPVnBLBOoYLlOMtH5gfaN/Vh2MAtPrOE3Q5
23FaI2bPvSB85fiV/9mwXG2OckeXpaxDZyeFfzlFCmKEL0LtnKWNxYmHisjZ2O4F
lYLRz8ko2aZzo+L0YhqBa/vLV/vjzV1dbnTkjOnql0xzweSvYU5BKgOAV+QO+R2B
PDmwr24OsaZgA7iWPXK94C337zaQdQVSGW2JcVO/sfW7XN6gBgDmGlAlBcud/Rd8
Ey/IUl2n0bgER1yjFcuiSUSTXmOwhEND9+o/2xckf58RR02K0H9Gw5OFX6hOwlOp
P18y2y2lWu2OH37HUuKSe1azmb32q52MsqdiVQURxqS4lKMHNT2pzg1+L+0FIwSY
QC6Lbkt9vhTdQkTR+Ur2e6Qht/xaOftBfmjpRoCm/piLUd/L2zocc60lSq1Wth0P
q9jsenIkz8szRpY+8CxzSH04vNttZYwJX4Y/4GUMWxsyciVBXFCXT2AFJ9BN/cBG
RG+8/4q6xCw/pzUITYkggnV/dKU1dmw6bhqklALhKo50ETllEYusUI0kR2AjMKzp
eHYJWLVjIeXGQ1L8YT3SWghOn/Yj3SGA9FuIinD9Ig+UGYsxMRYOjLosB3KjlwLi
tZPNs983p1zddlojNVqEK9CTDCHo+JQi6zgns0xlhO+SvK08Ltz9VqtCpMv1u71E
mKTWCdSmhhk9ZYYqudOmtt+q67sedlWBd5fCPPriVzkiFzih8WxeDVuYlPByjBCl
2Hn7/b0+Ev0e56pVzlrWxKaichruooXnfwQpdjLi7oU3LV3sa75F4K3JE5lQzP1h
PhIb6reXAcxiKZidCCyD2vO9QFumO9Q9zoJxjdUTXbwHEgVOEYUi6bOee043v/JT
R+ziCnw/IwSLLy2Rsq0AV+njhanBbgQRZaMSLUl2OpIY9TUWum4P4aQdwNP8D3G2
qNIjLOQO3XIM9hV7e9HomiUSFjJxdty9LqWerqb7pkEYAeTPUke0Qg0sEH8b1gDQ
PH/+aqcTNX9AAPwMODOWHewsj7iWmIOg0MNHozLpgD9i6nQe2gd0RbJ0fUF3tuNM
9j/co+YonpZZD8FW3Us1JuFeHGQdzfxni9EutIJ3OCpGu44j2eWKshCj9jCRBuim
WOUPnb78Ub4Im8cI9QARYUTGpLkB3UrRzwAttOHBNoD121HC1se5A9fIYC1RL/+C
hVr4YSvfqDkalkJtM4PMUd9dbmhVqwwQjsVvxOkI7Bj0jikFmcqzHouxgmMalXmP
UmQ4mvkGQ5APrYYNCqHPvygGnO2Znk3ueBC6PLdoekp2fsnzY3MAc+lAScNq8VoM
mVRRLjjKmlwWLRU57m4f9bBRG+fSkITQ89vH2eYvGh+iUpmQMTiD9Gha3eOPIhsy
oLNTBh+TdGyZhZuutBLs8HjWJ2zwg77aCMLa1Hl7beDWrQ8uP0P5m1PT4WZ7Evtp
Fya/BjYg96KJ3lkFIqdnaO06iu2B+tCvgqKIwFhYF7oj/0rxYlz1LdSE7Pz55x2R
gXPcQBVFMTD8x/V80qI0nX2eNE3YCNyu2xZKbHVunbJ6J+vR33jXkntOY/V3K4Pf
U1uyxv3DAIZJkfQvwPt/NkcCJNfXAUj2QoCumDfJdv4IY+BzwsfneMcLGi72zG99
faEQuFKT5CnjIXS/WjyS2FXwtlQG6aUD+PSjpRXidgJsVjofffTI1NgZTGOVM3uM
LGxvRvIj/nBLhgjh4M0gRzN3HsKDEQahXc2ItzB3htFg51GTQbNMy5/XGAkAc5he
ix4eelpFN6lraeZldB0ub5L+bkFZUOUiSw/NLWJCTjjCEuUEAwfqcYlLcXpo0jsR
WOP9Uox/dFt1OIrpxXqcVGn0qY9LcJoVyUWqKrG9Q44rG29dabFw2LwGDVYpqCNZ
KmTgN5WO0xElhA6xR0TiUyNEPTJQTymnQ48NvfrnK3atRPttWreY96wd1Kd3mvq8
JQmzWAX5DDWzZ4lMs2408NAPNTF1u2wYskB6DRjMz/ZkvjxhCXTbGWKVL14RZ+l5
+hreYhOISq0cbaqtIDBVqm07bguiZFd9Ut+hDeq5mQNkk1yg37hBkBVxVUONO/Nm
qgYyZ+EAlFw+1U7sqetB8adugOn0Srk+9nbTKqWLt3zxGWGzQi4ACzAGCU57NW1j
tq4HbCkF6gtwlS+TzDe64T5JbSfGaDJFx+G/64i5YgS2e35IhTXGhWiVAmy/7W80
dQHM7qYzIauE5aMciNpgBIFI6D7drpPkOVj25BS7LRQBXX8WfOt+xMtfi4hiy6ji
W8meaerNNucm30NC3Q4ywYuuCUT18KBRcv4JYPz0g+xj/x9Gioh4042MAEoEs2x+
UEweNunXw7By3FHzbBlFEm84Wk+8EhgVBw9a60xk+ojBYXgCGs+bdPRZCxsfnqAi
8blUt9LnO1+GsM6A8XkdUGpH/BjBlaGg//W7NC2KOLPvbNYyVyBfMft6KPCkKkbv
43Pj+YuUBef5SaW5uzBnSaKvlr+ZcUBiXiIYjGzCAMaOJQjKqi9IgCNm4+sCFcok
clDZ/iI5jlfyh+N7/9msqz9jutl1m31Tc9xFKzVimbLqCvgNl/3Zfgw9rBzj9s6J
xNOHrNmGNHUW2QGQpgVEz44NpaG9DGRnNdl0j0LpNe2904VK7Yfe/Y7XoFYYxO0P
rMO5P4WC8oIQuuG0ESf63/Esf9mKan7Koa00hQN0bNrGk3MfT8wfxqoEyaie4MSf
K9XWJxN5uegqgE2/QKUSA+54NvIluTClELx2oxX7jBbVvyMCbU6xyNSqc3pWIBWB
XxcShnZ7PNisNYydI+aJlLNA0gYiPURfP2muzWffTyosJ803DathLMooUOJh2AHi
hia0X9xxy30yp/ByITbN4pV3iHreccmq6f9BoUqNo0q64FyNYiq60SfS4ekhsfgA
KwOBLQZ8ue75EDF3W3R8OS2wKrGPLYvzcE2VfLIY1INmYG8cCfOesGckHJ4qB9nE
naycnGeQzPui+3PqrxUXjtgkRu7RXKueOpILm5WCXMh30dZJOU10hgwXAHGpWI40
I5A7SGrd7IF+pf1zExS5wA1E3CfwGnJrn7NqKlC+qFbk6kMVJrEiPDF5xDyf3gP7
Xf+wZ0sSoikXXCnhuTRu08RtmlL4Qrkn9ZcUQHsBDFJo5UZC3HKptO70JPrejPlt
zJQ6haTlWHbKfDHKQbGh5OHg0z+wIEMl0TxQkqRJtZ/xV4vUxf3j0IESRVaOmZ+f
V9RXHNhH0TIhxWKKVRzrrdBZMBfYQScjUd9zld60nMG0tlpG+dnGgfkYpeHKmzOr
3DO8js3cAB3kvPknLvBOB70HkEglgS5yYswNi0zPweYf7biBrCMGhzzaHI8AMKBq
pOKEwgKdgwxtgH6IwnUFZd42hVLsU6Px5OUvz6kVVWEEIXYH53pxlLLbLet+jRPg
GNi8NA5t0guEz89PgiBTE8Y6Ft/sxIbg+B2h9cfqkce1a2OYnrlKmclu3OmLToVk
mXGz+R+ApofReJemwC/JGmcHpPCU0Xo18PqIEBtXopg8UV78FCD5XxRn5yMtzvX1
dX+B+JpjiN6tNERmuQ3FC4CNqnwS026lWaUvL00Ny8Ihh0cBCWzJQ2+IZJ01++Bu
zI0Ia/1HUbufBwS4uEK1QVklipFqSz2yTJoQfVw7EeZqH6Uf0FF/+bKKgsgHlBpP
FiSlYlXRKOBhfCvhnTUHbFfzSV+CNAavQZsoRiKph5oZs4eyut+mtBJ39yg15hgJ
/PHREg7zYf2wYGL45idJff9Gffr5NvJ2+n7ZDl7M5zf3OMnx0BGJKzB92okh9h0B
AoJzNsSOcek3HSB6Won8XwhqyU9kmQjUEKkGHaMmwf/VDvgHHTQDno1gQWYNO0Oc
+pUPccbM6/LrT4uyRhThvmU7wj89KXOiFSTLZI8+A1Se9g0rVhjXzfsEAsKYkOPG
lRp9opvMPAg/3K+UhqRcWoC27W95G+W2rOvtVjvRFazycs6IWH63vpx7l9AW6BKf
4tuvJN5ogbtlrvxtOZuRP6lGZyI6wCsWHu7buHxuirkY3S+UQP0GZg8YPltPze+N
QUK++uli6teYNUf7UGuHt2KMdmK1V3BaOFGzA1aS2RpVHA74iV64W5j+R0duGf7B
1OVuq/ZCmQZadW2Y2VSYDc4pLKb5xmCm793iI47/FanBz74Yr+MpdeOF8kmdWQ8c
0j0v7YNgMIOy9hcMHR+HykH+idoJzZVvZHmTey3PNKIuCggzA5J8D2Y9U4FGMaQM
UNrzKMZgkR6ctSWIoQbvR9Kd4azX9r/HpEqWG82lYAzIRQkXUyam/cExpKbw7MPb
vu6mnPZbwYMJGdbu8pEl0pqh/T+wz7OsV6Czory3j2ujRaHT5PfoeNLrbVjiyBfd
ouG7lH6eFIM/X6AIr+E9Gqf2P6sseGW2YNGbdGCxG1ksOBFbMw73JH6okrxirGUr
YYHZm0c/b2i3NsNzardf7JHWsp/es/swBDh5G31tqQ2gKAtNJmyjWpFlcgchIYnI
KR9qbMnr8RAZnSXmj90ID0b2fnD/YuxeX77o+EkqeGES5yoXK4uhdE71p/KVlXES
vG8Rn7cxqvuEXDuPz2THmh7jsrmHCot3P1xW2Xl0No4Uv+RWH4gE/jE2bMxwudes
tYcHNOfPVp2w0e47+3dWhgi5h6kJkSRa7MNIgke9ddWaMLMoY5eL0z4RobleemRo
B7E1rj35QfbQipyXK7w9qMBGF0/prsn3G9zIv/BxnsbG9xlSPToY+NMBMDZB2/uH
WUq+Zta2x5W0o83KYiPpHEyNyZnS1vkJx8xZ4sI17toDiZQTP3RBybq4OemgHVTb
7SJv3gBLIY5nLR1BrWgzRrrA0B2M74Z5aQ6ZrFQ1B6T6HXyR2UGapQpycqrWpBVY
tkeJgM/0FaMQTzhFFBfMrhbFqgwEBaNXZrMzNQ/vn4MfR53+UK53euwLTQp/WyeW
uqs7Cy91TatZOXNCNSj7JT7YyTsyObJvmI7l9WlfhInxFxVepzqgyJZPjd5vjKwj
65Ntv+scZ5tZ9linT2n0N+mVrULC9uLby5hSESupt8dMIxTkMvmAAfO4ICamAFD/
cPce5Ju43Wq999F6cjdRrK7pGQ+Dx7SCgQVevlGRApu8EgdfZ1zxh7c14/hnGM3r
DJkJE7c+3af6QK9EM73fXk1qN6OToukBeFNYcg58hTZM3Py8JL7j1IoJp3t+UdLn
+Q6s38VU7QN4f7MRZkSLqH6rQ6eAPhzVfvu1q82GXddyr8WoQlUWkQ1T1kfyKtoM
7HW9yLQQWPtjVZOvAOwv+AebtLsADCD+cwBTh4nH8aLs9Jt16sIjAM21qlLNt5wI
HTco96U/UzU7g40BO9oJ7XRhqsiCQCMkubDoQTc14bFjakjYftHAvILtRrr7lOR0
StG0jFVmF5B7CEVvP4bS+H6aOHzG4Qvi5z8ATew1F98XRsKNFtgTWbYX0uX1i0Qv
63Y5E2+xgkn5b4DxKWzm12aFf28f6RScfneJgVQ3YnuGBvnrkEvZP/bGZAJjUn6M
1ScS5vtRxjTcARLkrA9vtEUiCxQUqMTQeK1PSZwyZ5C9Pz8QDnYj7aG8BwFv1mfK
w8CGoqbx/PGusHPwEtaD/6uQ/JdsA3JAton7hzfzh5OVdSfO03mYIrVNIfkPZ776
8VC7zyM6+A9jpZPI8AXy7fR7zCj2EnTRtfAE5QDrpXqE8+wSIRHvlYpoftVylvNO
dXzseg2EFSWoABy+shmKxEtBg8tQEVKu/YmhwUIoIgTBam8feN7WPyE/Wt2+7ta9
pxeAPhBu0WStMCB+gSzDt2D1mPJ40Xme6TZ0XuRvUM+6ISHZNIcEPYOlBzzgQ2bO
9EA2LVKyVDvafkS/LZtlf6Mi5ajDiaBJclvpl9sdliaAbhN9rVjveUdvx4B1vyRz
VcycpT3c4m82hLx8bvgw8Ueid344rKGpWqNR1YUt8s9+NbVgHNV8DuJfHpIYGZQb
RFKUraAArL5/fIWW2LZAwk0qGRN6KXxiA6hcfO2tKCgLfm9sYzJSnCfKjqih1H97
ggOFfRByZZ/ho08AMpPYam2S/VmT1S9sepSA2o8ZzZ5IdBxl5OD0o28GIHeZOg/q
MQdIstAvr2PZ/BsbsVhzAY8E6lCdiJoVjksCACe9DJMiDbWJJ+z0SBM9P6yWk7q9
es7wmMvZZBN1TIgMYXcMeAu1kgk9dA5M4ycj7UtHr0DlBk2ojBusksm1V26z97kk
DVHEIeCwy6awN2ELPE8rw/qKbhJXmHS3YVpREm4KY8vk+gIHH1GzJR+/ttnVE7pZ
cz420EqgAvCUNrgsB8rhtfQa86pGQiahai8jKCI4i+kBiYrwMLrFgjrPzNnJrj8a
EMrgthUiGn0JzEAslZly/7h2/B7KGOIVNeoZlinqUb3bziu6yqvVhAN8pVLDX1xN
PhQ9bn1ZQtpF0ODS/E0cWTE1BRyrM10CWk/109/6QRm63AJcDaYgyAKV8N9WahN1
otZcxpJEtsM7sZOCRPA26GWnPJ46oo9i3KFJK5+zVaYPWPBkfdFdLwNwqqYdXC6O
QBn26oNNMLF4KaVRHShHS5VDvYYAvk7RVFcWT33UBffjV5xZvVcqvD5BjELeQ2y1
w+a0oJ25eg3/g4LlpK5BhvIK7qqh2gh7zbnJSxePr6p7aYRMBTK+rShBqCoIDQ2S
q3nCaQbVsPxC7G62wGjJHU068y4gcENgbnhNRVEWNKflpvRIKip6ljnyzzNYDQhz
tyeR9bpt1/muA5L4wHRnWjWhBO80LJAkJKE8L2jMPL3V3mr64aYtihVPRK7lHIpk
g3wkBFI5qFxZRWrslIan98syptLuVBgkRDRzeaMOLEY8uykNDOLpEEnbXvAaOzcG
EdEkrGAnBs9UEejFsxfXWn97Qs1bbGS+JxjdbzenfBqdNDh0LVdx5I+3h6CIiAqc
bXs4rElHTB9uCUXgcEO+9P4u8bFbiyHV/Ku8lI8hvkizrWIgQ2nGmNwscrgQx2+K
Tey+Yrm4R9xJcJXNCiGqVSqvi2PHxMp4zWDH3yGnX4WzOSqUsNL+PE4JvoQM3NHt
iHCZuE3ckI+M6NAzhkm4fcviwTRDwpkd+Dolhy7bCZpvMIUjY1wAT/1jkPW8Uh1R
vMgdlQ+vIz6zfe6Hb/BhODoGr48j0UYxLc4zzyHuuswhcMrsjqi6kFvEia6ASkCH
gEhNCL2axSIfv3lA4CfLHM+G29MYCribR85Rae3LVlXx+Y73yysrUO+xJmvh1aMK
7LGHmKeKR+l3oRY9jkgpGdYa4xYVzQyMxr0uXXJj1954xMEEV55tun/KL8bJx5wR
KqjvAwF+i8h/8T0E13U3ePKi3bewZwSOtbEVSvmF4mxoLzXH8yU2tffP4X3uWZfw
zT0CWGmPk50BdWwMe2E2FTCc0pGmPGBQkIzwUeTNU4m1xwPZFC0V1olXREpL9MUM
D5BbYzkXcPySFPDZhK+WbKnAcYk/mCRxrDyHcwyXki0QYij2dr6mKyrds5QUEGKa
03zln76ZoUdqyEgDa7dZg3SvPXPw8J1iR0Kx2KpHsynoaShN0aK03drtxsxesoud
pjnmdOgCsizJRNwy8FP34MJaRuvF3LOL3uTY/ZbC7loyr2dO1o59890UeJQRaQNv
+IC0xqO5LYQncFaD0r3ZbPq2PNFXpSlj/kMvdzFnmNL2018TpRTUx6ZFKazj8uZX
mzUwyXxdwqyyH72L9kxTHEYHJEbjl2wfek+PYcZeaEcucH/59G3rIHp/rcLf42NQ
uP40fRxdlf1XfirPhNI+K3tdOrS2hqiolgNdGtSNxOUDbuTwcb7yh4m1bo6/btlg
az24fx0Aseg+zd0GyZL18gQXC6WPk9bOuE0tTCffuppBAAo5axsYNG15Fk5vVXXt
omdw1/hdxOEvodEIQuxpdAFWxZIU7oR1K4eRf1BxgDJISsqDBG2DpIEdoM0/3lyN
H7mjgN74NGfSU5FM7lD23+e4WU8xAzh4h5bzQx8RhHaA4dbStn/mrGFqkyT8DQX2
zHXQh4oMu8hzTfCrm9s7aTAcVcn23GsjrsmqSBsSoGsoWPnd8ket4kOz/1aNHjmw
IIFtL2vpnH5ysmhSKCKgK5sMo5/nF97wP8Yx1KAfh3hJGIR4nn/OxCPjCtQgxMVa
q2qMfdclb9RA4wLAoXfm7LFQBsErrG117Ss73wkKCEcDMfLGT3PPQNQALv+A12Kc
obnLr8oEZIskn+8i9VOp+alEyMr2SLhxjL9Vfu2aK40YqbyTRw7SZDCKu6agnXtD
7dehUSGXrI3DCysPb0cO/QgNp3J26wdaqeHS5o4Hc0nyD9Guho/K7Nl3GcnrYp/h
DIzDhXO+DLGaqUNoO9lsBGvaL3H8mupVF0j1ALZIfLAHkEJON8ShLDzI15TyYWex
HfqACkygFtJO6NOXNfDbxg4TrivuhJIvUwcIA8ZpekWuFMBthczHBXycb0eYRBmJ
jTJvgJ38EXijf/29T/MQBfo/nBU45bkIGAhFcrCy6uT21xci5IMHVumLDSI25AkR
U44i93qgyXo4NvYE2SC7WAzL/K0vDhpmskKm+mIrhaji8eyQlmzeXEg+GspI9iBd
9upOKSiEn6EF5JzxI9sr4EKgFfzjO/r9utz73jp1cyKEzf2be2Zazot0KkfGrzB+
LF21iuL8aLhqorfwqYoi9K8/k+3EdlEhKA6ycxmRTQ35QSywXjBH64VaIWjVUAh+
Oia6DUG4Aa8mD92QaXeYPvHJbp9ivunqoKrwzRhneiuFS/5qlzFDEbw4TjMj7uTO
6jNYBZzoDb5hDteW1qm1E7U9KVa6RD7x3Q8prC8K2dTyNBK8scyGyAMaWdS0yu4M
2xvzhrlCyiFiloDqXn716kThclLaVQqRNF8aLt3RQJ0FVGqSOWbKAAAfJ4qnIcod
w8GYqWaJ/tOLcVFaELaKve9czeFfid7grvwx1z3n1dW68nYbS4cIqr74e809jm9N
t9uWsdfIW1Zbton0k1pDEACljIa6u5g0hUxM5EXaIAPGoMPs3/07Es73h+oaf0P4
HkgY5LrvmBscJsVrYcQcJrF8LRviOu2W5uHXDag+WPYixJqM6ZKoScRK8gNDBdDN
9eZOIiZA6mfb4oY878i6liStkoiXUYMuZfsUAYzXkZ5dRipM1ONCwro7XrIQ53yS
8ePeJhz0+r0SkSKF3DHBbfx8+axrTZ6TZyEBqwhFvy0aLqwnZvhbqVyOQVgQ7OyA
wJrZi3oMleyBDU2o+QtIUI/HTFT3BLIKzjwkA7hkk1w9hez5R8v4nFVMB+erHpP3
6ZShtMTJDaGiUm76TWoNcrJpXDJLK/RWjKk3hUDLB7a/SmgSrsVXYNO/Z+6pTbWE
Imxn3LbvhtMCV11aa9ahfBVuqKLlX+kfY+F7XV4Ui650e4Zz/+XQQ6o+uKnVr8f8
teoGT50r16/XKCAuUgEQ6x7uWhAvNScRBfcojm3mSOrP2kCNJU/SVlhLJF0Gw3Qe
XIsg8/tdcV4h3A+4E5nXNPiahHlVJqMSCJZFZBE0vVhCf7DBeAGDs6KXmF8om6W/
iEt9iuqre9WiVU1XE1127NaEW6h3bKi/tHSs4ALXWiGUvknycleK64Z5XdYcBfEM
2e+YmGGNFIYH6XmCCdRwh2vk6g3Y/3L6UEnUaijEg9IEDxCQ12zMkB9q03aSBDm4
aJYAiyl7xTBcNcMu0DDHwzbRg6FmpSpGgcT/GBmJxxkzAU4q98bueTKHeZedpfcJ
VxRh3QQ8KCYW1odEyAcRURxarj7+fIGuyPXFqgMGMUoSRNkWUV/bBtAltHaRPkV0
9zPbWPSvxPeqEO+HeNhnYfDq4az7TfJmpHsAQCZVUz2TbXzjeFY8d68db5o5VoIP
8EYvz9QSQkp2y2Fg+pXvKTDWoeaG0WhNmunhjW6+42EJi2RnnEcSxEiW41bstimR
Y6akr9oPE0esirgSK+Zz88khS9IKfUAgXV6G2rupiEXFUmuhbrCCp5lB2J3I/ZN4
m5I7VstPDou6B/mKn6xDjNwX2F5v+aktx7veqf+78ZqITdLmj0y9HV2jJTPjHj4z
6K6IKYBKuacCuNzzVypHTL76VBdPCRXVxFAYfzR54m7v+JTzypW3gXoL8jMq3gy9
0MVm5m5Vi85xI1GgqAPWUQDwaNdbbg2Nx8/f0VA74b5XcMcKG1vApRE43SrLWw6q
9pMQCKMdIA01GhwvFuTAQKSZan/k230PjMdy1rqsqrc9801x0Ifdm7y5Pqftvk+V
L2dxvdzgaQtW7HYX1sHxmQN5kebuQeCzN7RjC34s7vOSfp004Q1R+JHzbmewxDZs
QDu521x9iIQlReOmBeLDtqLrB3GXQwvaFcdT95vmYsntnI9HyQ+9kZALIaY++7T/
PeneDKLFAhBMKzAcdu0TOXb4LT8WiGy5LoKKr8VhRQ0Xx3QsLaFoWnUIZYfub6hH
XKLl6LwHnsHmhrHBbrXOPa8JMexJzCKLGOpj1u+F4TMN96E/go9T2Sz5sJWg3xCv
44oQVNNwvR83K4LMXFzg0KrMjmD6aXuYgpiSOSXDdCmXMM2v4Ocl0pUOqXad+O8q
lej70jZEQopJcUlOmr477IIsAcI3Q0PV20vjRxRyYaphVQ+Z8pBeBVm+UOSxUCBQ
xGxue5NV/znF0uj+ELFDFVvFJHnGZ90sZOgIQA8hNYNFi6jd4Mlg/rFjnkV/yRIT
oDGT6H+AMBKlNO2dn2ran7pB3dnkO9EHObdEO0U5l3sdoqlF2srlah9eXdcnEjCb
B8nsN+Vy3H7J5EOwyjCSt9hdkZI7/OlnOrdIUHM2Ofg5G1h6LHf6bOHEBK2stK/f
er1qeAVcsD9BjuVgaXjVsXMP1RaXp/uS3xdhcztyRkQiRUcid7fcrzpEuwTUK12N
oRxHpjtdWfChuZ/aP2IjRaziGWeSN3lY+PNUBr2eA7vudLjuV8p7NDsHgX8aTcyk
LyFVKA4TY+/0vIm/waQ08C/S6RI7166tLQ2X6n303sdLR0e9x/heXj/iYmQAfa+V
3AXueFqPvug4Qb+kdfzMmUJAy7cFPsasJX9H04XU3tAjA1LgBntxQrNbNgy/QhDl
iRiGClYmqQuAbiNIVppVCCa1pINecgYN+6e6iFZYWXDdI9zsVDN1wfGvvQl+Gfl9
2V6JAaPxhYl+OPJSR65XdTp9sbt0seLTUzbdYEfNQZjllmlH5PSRBFT9KYXuc7nl
IatqC/V9E0zOEU0mBx0CEXrw6cjpJ+Zvr7pcG7gr7C/Wt5Dv1i/Sol4Qzm+WO/57
QpkFPudqPaYIGrClzxSp+dzZx1hbqRnN4pY43HDE2OYBBVXOAhbYRXlfT4+ycuxk
csPtUE4hrBbVvohWusNpvPctftOnkJbzDJKB6NMkLy+Du+4FXqgen2hpCXcZWzC7
hz+0uGK5tbiMoClecN+qS291YzRrGxDYvWm5f0Y8zbT1kZhCIhZg3skGp0kYxc/R
RDbiZppXSRufEsxBMPm+QrjRYoBCkWN4XJlpT0bSdt5SA71YDPWr+9wiPx35r9jW
IKBxMS6+sAGKFDbqPx/Ym7cZIaP4qmVxLHF1lkPKcxGYNgsaD/kwk4ZNhyllPyBO
oKeZX2/KhXQ3wph1vOeme/oFycNMTnADDmQpHfepJzuznMEyN1vz0Kgt/QkX/WME
C0PfQFM8YahWHa7db+Q9w4zkImFQLt4cQyuQZZGEIQYYLH60xByAqh8nOTh+kize
LrZRLFVVHT6y8Fp0DXS4+adBSzlzaLVA9dF+2eua7jdOpF80gE+vhbXg5zR50gP2
s45XvSXb3ySS14wjmnghxbbzDryum/toI1HwwiSwhvfusLGqLBg7wPzAkSzCoQ3a
fzXzQXZl7khBtA6uSiaFI90KBNjRKjP3Oalm6Vem6YvOzDaCo+m1i1yzF1IoFiOU
jaJ+EnMX+AtX8PgZOHN7JPFUDqBgK+5R9ha/XscOocHSaykhsSZADRLpsY3fLtQW
5S+VYsnEO2z/EdVCBEFeMCFzSkuML6flvrOuM+JLpKWWO4+Qr6RSrnm+2iQWVdk4
vzsN0FAwMgYu32J0XJsqB4+uIqwBFOz3vU/jh82pIoDfq9u0oVvMLHl6+zi15Xj4
RruyKtfWjJt7+pSKZGMCeRb5vgAGUCiQLJwvYq/K778Aqf40eA4NK8A62Q306dV/
gAgtrRvE1Cs3vTKVDeNB9HXHsWL0g35oK3gOdJLNbU7+VainLZDcPie0idv7Na7o
+dfkkQXsbDy83n6Bun/ofBwEQXX+Z9G6XkVaoJQnY1aDT2xD64sieBo9t2TFA619
j9x079oZ/yyYx42oY+t8XIycjT0FZCpksYLjyrOIxbXanIG0kKECY9rD51oNgSwy
9dN47DNc0d/bTQdqVQyE30iRsZyKJpMWChkvo8NuBbGbSMvJ5bbueqyDHl+lBC8Y
LNxWbwKVQixvtgvdwgsEpiXmOiPZ3U0Ho4vC8NzY06KOk3AfdEIdfgO7ngYqCKp0
ywaTj8JKtmZdEsDOEsK1uf+jOys99F062ArRsWSIt82u1EktFZ1iMrhUVFu3lzQl
2WOkAFvClO0gzEh3GaK2NghYvhiaMKZfpA+4f0/LaVk3RYJLkg1RgI86+TV2unk+
qKFtSPwTAeLPISv8Z9Z/khFP4SRdLet2I0YlzFhoZQ45ZWfP4R4bLlm77atGhbA/
HFwJLOIsOJTyRAYqXFjqCmPEv4f+ssU/gRCJ3VlaD0yl4hvgh34evkT5YK3FODSl
3ien1a4EBR+vF5sySLltD6VWk2nYhJweTJwJMkEIVAOc3QKdMQ2imyEheVLPtkny
VX85YZo/M0qAFlfAx1c3jdXTWooIqfRPbZ6GA8RcijcXkS5V0Gbkga5wqEGQb2Zj
FHyJj1uwV5BdzTgSOK7K/MYqcdC6ERK7Abi3sl9r15oz/mS6DLKjx7rptVC5sSu/
D0t7C+8GS1oKrdyhrpro16vK5ndgeWb6L31wK+z/HbHJ4LvPgURqsUYLLjp/CX/1
he92s9R8XU9acZStuIfkcLjdn9ecsqe80oYpFn/3vuobb2SAEmLCmNkiGb6O7Grc
9Tpim9cEY9ewtdRk2ZV04p3GQAy4U6I1DRkwV/hsI5FcUrVTRZxXuq284oy1lmzv
nAXNjEiDKpZQXo+a8fmRm/jhN2m/JLrH7cQAbYAYxFnZR5MU/dunPWQRtyv9Vlrc
qcVlBKjUYBzrHFbId2hQ3DwtP03W0/9scpsViaPieXIUwWXlQaTbaw5r9oNb54Di
O2F8N21Uq+d6Ba/MR0fCpklvKoRU+kQD4MV6pQtcNnm/v3/pIDfHHNGN/cl2Wo6S
WzWI8nt9Yome0u4gESxseGmYQtLhQ06pHOrwPcMQcg5XncHYY43K286YqROMOyNB
CcY1YJ5lPD8ITUS+H8GznauzvTrkl9K27H+0d7NAq4icbd/JfVbKyI6XXvYy7uwJ
247B9ptv4y0V0VXVPU4Vx6IXSE4KAGYlaO8rB2sxcOzlMuu4/hFAJD79FrbDXeqO
IS9jvATdeM1RveacQ1T3MQSNn0EooThTcZ1JDB/i9C0VIDEEYKHBeHBCTc72Fu61
GqOvL9DQuS8SLYZ/easn/rJQ91Kti2dUvtLouUni3Q4+wCUr8b8+YxerYKlSlQA7
kUd6bOjWcm6v7TIh10R3FDmM9IAjTr00j0YQN6NR0gpIhz0niEm7UvvAUv1AvgIU
kcpyyOd5ntdaUR1Nyrh0vzp5cQIw0UWY9yjTVMdRQPSc5F/2ltRTbv/vQ5EKNlhV
kjBwHUEUyxLAQ1tsStDfE/ud6mOu9ZX0kyyM+ohGNIbFSMBgnOLzYWy8ApCawTCK
8yb+jjSVUXLNz5M4vWgtJDJAVDHJ4lGh2PfJ0FeitLMcEHUtYF9DuPmppdknKVog
XKq3fkYjNuJUWxYsTKMGRxfzOTUmJdkeQSPyAgPBkEypoZZLad95yoPE4yfFFx53
21iE8kGl9PSVarnX3hYcF+qbSlhGuUqUSTGcaInwpctfPZBbxzJH78Hlntqtwh0S
6oqrmuLb4Dv8AncArMrmhWJzXeAXilbeW7yTEjC4jBJO/8zwciK6uMl9NwauXoLr
tl+u5vi8Z4QSOQPRQx3KAOyqTNlaJVmWWWj4b5fX8aBRL+V1CnWceG4ej2FpslXy
lWeqRkmIIcUw8yB25j3JBpV0W498UxYf30JybNN6d5hPfcyG7ov7IN5X7rf9+GTD
AK7WNoC+RLzFtmJ6cb3pyK38XFPjHnj5c0yUoyPXioWQ2RfZYTUL3AGMsm2UsioS
h5ppvY0uvnuTMBJCrqtlboPc4sIHE8CPNFzTgS/ItgIuu5Xi0VAalgXmNR55CUsV
k5T+yYgpdpu+THeK89s0OiLQ7SwxE/3sO+Lt25CGYb6fqEjiOaDqNp+jNkDtvXbb
arqBJiDlptggd9MKd3cFQtpRrxrAgp3OKvcVnztM14RUWBVO678wUFrF3fXCv0dA
78Tp9Ok83e6dwK7JRYsVbUmtrqrnaS6mn/iYAkN9hJRm0Kz+aclsphchDiLZDgqJ
sMWoiVgoWnjUFsSKPQjuN6Rxs+ikBeMcctX9hQlcVBuvwwOdLbLumTkckb3NNxqg
GIQGR2H0h2XdIGOjdgc9DJgB1w0HGOS66H7yQh6ka7MK+FJFMZuHwR62Q3A59CVn
HFVlnfxUf24zbuyVQKR8yg4wADmQOlrTZRMQFdxsWAI33ij2JZCiFfizUUtNe9+8
ZwaERLg3hVzCqQzFC2XeMHku9YOFGzoLTPXjXzaXZp7EldtQMBkigm/nbTpboWyG
eQ3BRAyuIdazelIEYaFqcIioe9/HXQgJP1GUAfFUmLtUMERktfqTm/0+p+tG2qqG
P2xMbNJXOxaa8W2Hm3WsKjezP3A+pMeHEa0At6LLgtdaJ/XNu+Hn6bHR5Q3CpAEL
L2D6eeIZU4YPDWm27DyF5aNOlCjeh9OImytjkyeOAPBM3BP/7YUWJ1GJBpqq18uh
QOVEiHY4OcmDXloZ0IdeZR2lUqiwgDyeVNZNYZVV13pRJ9Crez3cSoWwMSZx+tTG
sslriFpmr9QoD5q13GNBqWoDvwZmpESOGnn/owLdEeTSD2dLq3upSR2ynqupwPUA
JFJDhBfHTGT+Vcz+0G8ZqzxyJyBYM27+w1vmjJnedYnhN8Bylgnhq77OQBPMrmbA
pDUyrCB9JqJu5rh78bRwe0hykRcamsiDfQ6lLkrpuPqMA8jazMialDg0pA5gwUcV
zCeShHp8vp/CvSldazY0cWNua/8WUkGiX1k0qzOZ5vPW6m7pzATMOqKGWR0pZupB
emAMWiG1JLRopoARsJLaSJCp9TAGbg2hsKhJ8kow86qMJF6Y8DKBSGtC/0rXIyQo
n6rHOZaqBxwn7jq9E7KnLtHzJUAn5ndaycN/BxBrOoCEahfpJAPYVOOQVYnG1HFe
JQUczOEry5GMa5lXJCJmrJbtNgpZ0BrYLNbRbD/rofZPXlE8vDD7iyQIJ/9e89qf
EMCuupQvhA4+q2oeLkqY18v+lgQ64jFwDmXsJ6UL6s/L9cCta9GjYihcFwSBjhdZ
vxFil51fsU5iRyNhhmDNfJIXncEPh0azb3jsmHdp6V351f9tPPcT35nX5xoFL0BT
hmvXhKeiJZONRyUddDCvvMZR39yMi25r8eaYYMQwwcwHZWhdxBiykCoxhfvk1v6m
PhBhFLKeua7cjPHBjxkUYW9Tpk5P4p4Kagn+Cl9ZH9HSzenT4fUfeNFvgFdcxOGl
Yxxi/0CrAxUOA0v/5Ow82Cb6An+ZzhPdvTj130wBiq4RiCbjWkFTrxbRavHp6CPp
71tGSm1zEEDiFLpYQxW4khcVFOrafqjbCISoyifoIgebdoUULqjWbEIcIyY5mVB0
6OKHdiINOfd+oeCMBjSbVGWIszQlixICJhQk4Gl7fE6e05xFt7+weKDW04iR1sMu
PeO0wBT0ifUo1GoNOY43/xQsFPjBIGvx/f37r9RhDl4mXChN/eLUCszJ61Ih01QU
G8s5/lRz/YmeqTwYBE7a23p5e1OS4APrKENQdqBt0IBDcvA8B7zDzmL9ES6g5Un9
hPFFQwJekmCfB8Ce7mlnj5CPaWw1DjhlnY/uvqv8YIpLrR9tpS0hGk+7OjJV8ZbL
sJ9/FBWnaGCnofA/7g8X8q960DnboaVvfSogdvmSImoXKKSepErqW1O2OBwX/tsz
Fz20DXdiczHSmdDD/tSS0u7g+g1izFFZavLuilEwbc3vsJO+YIgX3sIkJA7E16sI
4MHJBptToYG4ik8PATYSiOLi52OaWLtDe9gVBdKLhRDPwwQMPxGZtHml+gUt44S8
4o7c6L+kuP6/HHBhWjc5Xy1A9VSjr3Wy14AJ+LpxXBB0+IB5Cmfqg2d/CVWb4BBm
T5LcnXDd2/p7qNarRghPbngolz3o4YPpMXxj47CYTO6eY0JSWsHMFeFUHOuI1JdP
Z+P2/8cX4jpt29kxRVL5vV3K8FpTBCp/JHpDUjdh4lBXurkiHWc5WsjTmkbsmjvi
vQnNhCB89RYTse/8KCU7vCKttyfgGpVioqUB92J6R+/kWVss0ZxXe7mwuBNH1Tqc
ECI3BIR1K9te/CcqD+FZN59K4NVozIHMalzydTPrCwiqXnMfbw5kP/A0bme55sgM
FJwd2LhojWkCPgL+2xlIllM6TcSbEnOh7RgVXz0uE0Bl9IembfqE7Up+IVuPrFAi
eQFVR0kYIq9NJ1qgUPP+V7PajHcHNCGmsIy/vEmFMpETUwfPJXHcct2Hx/Tg/Ekp
aWnmWzGkWxnvH+LidTwClS2lb5/18fd9GhOPfLrI3/vIXxRVcPiFnm31POCso9zK
HunUVvduBF/xa9GucuhOU4TzkxvDmSqlTo4Xk5DJgqEmnCEUmEOockM7Q2wRD35W
h23JcPYcvSUd5qyS1JnKbUIRYw1JF4O+irVUsiIOipOgd0xI5bZuK4D9odVYTI+g
mAYrGkltC+J+q7K0kMlC0ituEsr1w2ReqZ+/dQY77e6thBLMAWwA2PyQEIdo9p9g
QvOt5aw/DwbcD919kAMHQHcr0NwAu80ZzxVg7BsBb9d44x8gQ5LG1Qej6enPMUHg
3kTfcAojqWF4BndCnhGem00Qmz1dnc/Cf9bs3lkLbIYVwg/ZAkUklBq5sSUdifnp
HzTYJlT1dVublHe5S0bVaZUMT/gt2aD89+E2+QBATufg5G1CEzWiUAh8vE8AtRuP
9fSJgY58XJNEU5ZZ5W/VBGHDaZeNsLfO2R0YKG+QSyelmV19een/CrHzEskxdOq8
RLUlZt5H3yphVA02rR6Mhwfs2rosfc+VIR4HH2JQuEZhSTAGt9eFYfbFK5DrDkqt
3QS4+ydhgIDg4NZ1a4dTR6XZY1poZvpAowTsZ04OLEjIYw2jppAxY9U/N/Ci73IY
JuCP0lbs8OSFnRTfEHZomnXa895felsq/01EgnZtmO7+MJg5SYvl3rpAUO35IFs0
X7dsNjflre48Lm8e/2m8BCK+Z+2A6+8lFYTXWEGcgDvdIQEtfB90AGt1k9lB8ZsU
0ANkWr/THE0AzQ9//hh6oiieaEiLTJmzAeg8GH4ZLwIC4/+VCGj8YfXkz5wjKK1O
KPPiFFpAGndB4JX1vHpjJhjV26niHNk51wSOdMSUnDu/erryiDDSZHVrFQiMx9qD
tgX8gYsp27wdUsfWkwvhKeaz4LJ4Fd/P8Xw1D1k6iQ89u/Mn83yaF3YNP4o+p+Q8
7LrXZ3jAe0Bp5ddX4V2sL7msv7yTC2eBGANoczBS0yM7f6G1uSORxBbZdPynbSlk
UV3/k3KPNV6+xS6Um+82LA/tPWElsIh8dle5MRLlCwFHC/3065v8ffG52wLcYdQQ
RwGG7LkO2U8pHvzB2TtwMkyzxm9w/Sqzl7OF42CtbsQrX12waqVdbTq1Thc05C2m
k7IXbyIRE4TIyxObSQzzhjLiF9W/TTLpYPaBOijhqgwY0Jq7tFhjvH/pQbwSMAF7
72XCiOsKywp/Atd06MPMD8ka1sOH627rM3jPHHWu0U9aCtihnHhHEJPdyyMDtJbg
hZa4G20rMuVyJcArOMaXfgVBNrs9CsqsGCe7TJBP96n4m15Sz/inrmltwB3r6KtK
wEzDYtSFyPlHzPzHSd7p/Wp1amSQoOCHiRiAw0loCPjfATYB/TPLMNH5eL4GmQcE
D6ef93ojbOsVQinB7oKGJT0eZS2zg9xIZXHbR9KD5WvFq1OdBBeb5jyiEFqMaH7F
aljvO5RdsB3XvhJYDJkRw0iNAGpNeZq/GI3/+OnZGObedsxCJ8g6hU3avOivaf2h
Gsox+vNFgaRlObu+EbzDV37SqwsRPbeRevrR5Fm4oVF5Tyqq87cFsc5uQiOSX+GA
AykD1ER95Od5Q3KoMJdf0D+kxC+rEVkZksNEjQr89mjwMkDx5AEPtorWQFZB6mm7
qxZibmpS/Dnx/U2EXnfIupK6lwl25Kn8bPJT5Roa0Om6YtSXpr0In2J4RSJi2syI
wxoJSq/ozS5FMKhipK31mTTQT65g+hoXAD22ZIZGQ2F3jopEXJcLtG6iuhLPT4Mk
1F18iZuv01ajHUQr53mckFbDLVarQ2OTjHWQcrfYRLJkRfDTl5IbjPh74mLM0i3Z
b9PhAqmKmbW6XZFWIwv5u4mygXPuGxhLHFlzhnKSCMCkY9eZJYelV0KChS3l8B6v
5MiqCqouqY3zUav8EScZ9hvSrvJ0RzWAL5640n+sW7paYf2lvikMH61fZk6uH48k
hYWN6t5+H7DnGgxHXvvlie/3Lz4Q9DewjMlFl+KgDF5d82drRp3E2IUcX1DwZBeW
fu7jYYa8QpfYM40lVtWDjCpwQTCpitbn0OKgU6E4nZSVNi1FIAPj67Lsh0pYXFVB
e26PbEZxnBbHjUhiHJEdN0kAJ925vd8ZAibEqMVerg2Ntks8KZ/XFXWhrTRGiUBM
xrehP1+xSagBTpkoIRjsYXSPkfThqVdEf1iHmBeYNHATUPEwxOW7GinlnzRoP4nP
RGEK2RGnggq40uFMUGSAib2Z1bDg1lF0AzQTCfT6VL9nUZBiW3DP0pYFdj4CNMnC
Y2j6M+BqveVC9932OMOT+PHCB7okF1VoD62WLWURBdqkcttO8/3661P7PzOjPN1c
OJq/L8JnvuIV2Am0bdKjx1NS6R6f/ItxASzsusExY2wjJD2IlMEl2aIBF8KcSk1u
l+WSYJKU7E9k+KwVBMwpGh4OZpIrtLi2zkNPWS2uUUiTlFhIZbbpe46evC7gpJMS
K8hL7l4pYOmHZwVllY/U8ibqu6JBkod3dDPVSAvVr32S/ISGT0VRqtKeYSIqGRwu
/lfOAI0Xd2kdAT0QOhnHMpObtF7nNv9zPbkYmW2q1lR4UAXigD9Z5d8OXx2XLzjm
McgndDyavSTjhdcJszR6EsWXlMDTto0zw1QzEgh1xRVaTq6CMreEz4qbpJ7txl2X
Vr1ISB2lHztxG2zV00YpXpwpjRwj64w4lwt4eY5KU/QXkDX8WVWuBHsnx0r2wU8d
c6uvfzmm0fnLNj8WylWCJ+jZNtlgftLPMrpoa+wQcy6gkqFnp4/tjNYtpiaiFFIe
Hy1IGvcwTalz6dhPTo7EfIZO8UleAsAnxK8sm8T5BmIYpbVNoNiGYSpcoHQJyKFh
hf2AG8Hp69nqgjlyb9i9c4aHN1KAhAw/tsT8AysMmFz/32kb2W9KxJ1brbWhnshc
FQNJgg6OigM1H6P0MkG2I3cIu+xuVqgEEuSZU0a1BoINR9pn9C8CVQ5nsOlU2I7G
aoVmCIesTueDh5rdgN121TvQU8yldb0D/zgrrDjSKefMGb0TEBgpssUdGpHLXE1u
Uztcra+vxUO+KQb+Xcl2moj5EMX7Yt5SNliRteG50WXRDEJ3Wsl8tYzun4A9/rlP
7kxP54ccV3/+EIOQm4vmjkC8psXXlx9oEhSpT44DjktnRRKoGcLeKUZ/GNtlJdh1
Z8LEHzO5eRdm0iCl4GRSUWBGR14RT2OZzD5LDtgIiBYRbNaoEuy5wnu15AbOt+zm
cbGzXyeNglWHnK543F/EruZ4akG7ENFtHIPcnchv2AbqIt18nHLaMd8L1+xh9IyX
w5nlLkbxIhs/b/2Wl5/fgHpfGGtD95P0khzQKPwezhg6tbYfUN1Agg1BT9v6J1qB
Pw96qJS6SMIBcHJ34WXf8ISaByHAM00GZ++JahV9b361a2xoV3CCeep4+lHD4Hdo
sK14H0XqAGnuBne86wtTxt84xCKLHSl5iijfitD7T4/c93a/hp7Z3O5peXMxlPvH
UxNeikHCgdWLyBFegIrsGd1ENI1/rbXfY3ooXu5N2QErjbtAqlaWUjEUMUippxrQ
xa+itM9hofTzCcYcVeh6BBCBVAi9qFUMYAvELmH79tvI2Py9pnmn1i+eOLfS4ZtT
IdgP3pRqwS+CYeDxry4+WHhVwdi9DOHTa1UcAEaF9AFDIPBgSBQNXQrsX7i4r2jm
ms0RVanNHUK10603lbbKLxlqnAp63+374xpK8eHcXqY4YWJTAVFsw47ntTOdJFSK
3I/VomWCQ9Q4fYNZU279s0cBrJNedcji5t7qyW9wVPEjYoLxiFp2M7FrjshXX4EW
ozttenkaxIxDmSR+IUJK3VcOTZGEiumpXs4novMZbDaQObUuavCTIrUaKK0E7H7C
C6vtG5plYN3aZCIgN/18XLrAPK8Q89bw3sdvVi+OFJw3zR807Pb92MVq8Jw2PX/b
tYifoQ+KjlXdBp/eB56ywf2qttjmbKvTSqu9X8GZ0qDpiMhrjYS0C6gPKegfbj5A
fin3pGW7Y4OFehSn81uj+RO94ee2UN1Fbva+H7tqVl+/GMOKvVbIcqJBgmSCQdB/
6HZ3eH++JF1iY1YRy+JuQkgpdEXfDcNIXTdPeVknzLJHw20HJU+qqY8SMpcsdGEi
FelwEj5cQPUk0u/cWaTL69c6Fxktdi5JCdF0U8huYy9u0e8AJ0TyL0sr4W/DAn4S
0rj3miq34utfggoS4ODT5lSyvV6hIsHw8au0pW9OuadoMrhezWcrse7k7ufmfe3S
/5RpH1GyCwYq+tDPV7bFkLbtypGxbldmnhpTz6G3U5HlfojJ2s2vXtVI8sS/UBpM
BVAPIUNxdYs3S0yImjiKjgjwrkUeq0uW24/InNsDo+0G1l/iTAdXCpcxWrl7no8Y
yavCEy/ZkhQxZ9zCJGBWO9jgKyEBreUnzdUqjcV97XVywPbCoEgbQNdt/wpOvqeH
7Ek9kKLFN3IJG3cBe2+yO43quvyDfsrxHJB+EJG10nBNUVzGb2GpAPY6tjciTy0o
XgfTTNAYyW081LpQDN2g7WAUFD7aSfeapGEPKDzWjXbSnvs0C6O1AtJbabLHi9B3
qKQqA61e2BCLmnSTDgWPc6AH0+S7sLqfLBdplrGjljp4IVEbT7PUEqtIAbQT584K
7onYt77DDU6Kl8y7eUqjhwxAtc94QkGNsfLWy8IAyxYyFBpxjkmDoQ0sbrHZ9aXF
VCLu9qM3yhj+9hzrhH5OrpXOOfkJVy8I8pAYawB3yFLJfx9AghLp1oct9pLYQuUl
+kogtnFfHerJ7SZHNwX+0PRs01Gd1601O+PyYpbCcc1ZSS1VS9CStEGG3Emqa/ZX
GUSR+6KzWCAyg+Wskf6h6EF1+zbfTz7tqEhUEVHQ05OlwkE6v8PDcb9bMlg8MZ38
Iusp6JuMAT4lFsBxjkOoSiQn9f4Mf7INc8TA/rayTzoPssWyXiTjKmRnAqkQGCIh
8GYbJccJUSKOkQ50N8xrvigr5N3c6aYi/yhgsPlaqRR3W7ebqKfiaTusz2fOc/Av
d+PTZEezwYvyRANezSSRKnc19XxR9XIrZ49WuMbUFQ1/8lG2pMcp3CR7fqkDLn5G
JWJhT4kvYaDTJmyxIXb2Cm9jh4zs+Sly8iw0g66Ig5oeYaA6eTpaiwhqyEUzmwvy
LVSSpXZyI9lK6W9ZizqCA6xV7T7NiiXvuFOoljiX+mbdFg4LlYkuKyqfuvOnBnKP
LEOC02pKt3VaxfQdVIy3CpMF5NJkefrso1fPQ4Y9p49Pc1iAfF4Jtez5Ba8MQQcR
JRQNSDCGZAVbU3aedj1UXXJaRgmaXTV1ck6Z8iYGZ9DG5htr8FN499KMuRigEdSt
vQ2zddZtkDQ5bgF9x5ER5ex3lq+2zOOpRe58YBi/DmchvCck6RpmDB6x+6nNf9kH
gMa19eW/ylm7ltlfWGZ1hEUQ31B8ReR2VtRKInWQzcfVjAnqa9GTC97cXGQt/rGr
YETsW4KyhLtxrrcvkmDDPtKQ7FGlMZmpBZ1DIJp7v8c45vcmL/PchhGItG9q1cVy
qs9dChJbTlHRDXaTJFfpYtiGMeJOfydMJMw6J8MYFqv3h15z5yO68q8g3Jj0a+LG
tmYIuOgDIYTRi201noHf9+8PToLzXpotzwXBJNSxdsI+Wrg15SlgJKAdcHBCBEuP
CGUM3BF45P66yXMxjRcuwyCjLR1N8rh2LwIQ3IjR6LRumq4TWOOGyN6QMgXU8/FN
UHpwLOBViJHIWzH34ZOnPd9UyfhynuECUbr80klzs1biK5I6s0ay1KVlC4nvLaBJ
UYoAGDdkBfz0MAlXRK3+/01WjLXgKk95aU9V7fKyGXLCu1RgSyDjDpIiCjAZi4GX
wlgBC2WqnCUsVGe+lHrrt5kz5xV/Q4NH/I37XEgjqnx1LaYMlXyLHLT2i2d9UYaV
b/X6aitMZFegu0TfiV65dJCp3qMgmrZgGicB0Db3oyysaY28pu+uN+WkOdbmAIDt
dlaGJ3v59M1gemtIF6mQNc/imHn0BtTkk1/6/YJsoTDouD2LnwhFSQrXW95rocoS
p8t36Bxleao7vFlTdSKOc9A+nVroGDZNqefSLPOD0+Ow7N0/I362u0JrWYkEfmVQ
B4KwLFbKKPoOWVMkX4mbJOpFKDHuoZFJ7RVa/J7YyMlDpZ4SMQNKrTJB5wc6opGj
2Cf87zrgI/yB6kM6RxVDS6HXDEec9ISon7dq1Q31U6/U1gY6nY0gyEncRMvQ9J1V
cHXSKvoPDNU6aMeDlxmEpydy5T04LVuLU4unXABkbD5f52syH37ty5nGxmxvFhiF
yF9CoIOO0tG0l6gDyX7k+TgoWs3Ve/tfD41HRFKwaZ69+AArtO2cv63xNaNWMwW9
Elzme4r8LfRUps5wL7CpAMPKl2wzfupsCSpcLUKsBAm7R4vXXeJh1keaev3uVU6i
ok8ElUi+kWq+qd1OnbqdjsXfZl3QgunKnRgB8xpo9R7drJhXNAKer1RUZP+PlLbg
6uB5P0CtBfZhZOac0eMeGuiWLIefnKtXMapDF41/IopGoqBzma8G+HXpGx7JmE44
EGOt3D+rCiqgX+VqnfYrGQJAYHAq4UwwLclgABtacTgfltifyyBaE+5i9DSa6JIa
615u8XhltrAr20+tvXzr9g3qikD7AzBzYTgZAlv4ZKL0ItM/g2JxbFk0BbIs8ycP
wmC1UW3PsBIRheZOeqwvLw3lzCaGdB5BFc0YZsF2QDhENFf97njvKKNdiHKBCnlG
y/bv0yMwub7wr2jIsnJVzZR5iZMqJHWIKdEzgRSQ/679b71QeQBQt1JdultiOzg+
+djlfsW8NGLr+3+KJpuAQOMf47g4LXo7VIeFvCOP+dpEbbBOo8/tGaba+ndBqyer
Z1iu+kgl37E2g1AD5kWVHqZCMPpxbs9NUTv4Qjkzf75R2pV+bMBxVsvk8LnQlzuL
0BGrQlNAE121N0TEPeJMmLDryjzmpHCqFp5PmNiCys600gv7XBHzdLXKRBpDGTQS
FFbz8NFg92OUZ+y5O05kkVXWhrjWS1asjtDPb8+DEXuqYiX6spSCUkw9k331G+o8
uXp4H5rsHTD1m+ScNE7PaXwlilMaWTbP4yIyuKyYznEzecYuLiQNOMNBk92KguSW
99nlrOZe+t6/vwjsHf1d2ypTRY0/tvEEEdJFwb9eeqS6Bo/hwp1NYFVTUFG98pkT
dtjZQYnsQAi9oXZ54DJpcoRZt3xBCsuZcw5vst9GDkG16v1yqrgPJ/S3WKBQG0E6
OhTiAzeI04ht4ywjhGhX18TQopcFvm0ra8h912q5jA3I5agV+TFoGER0GCW1/5lv
GtxTsZIz9Yi2Q1lJHdz43/X3OqIpYRetwY81wzWcd7UvgMOo9R9ajDCSMuwtTRbx
qrHlYaZGt0CEdmwugSprXgIWOwIoijqEb6guRlM/jdCgzEuw89jMdF0IO0sXtx40
n6x54XvrXkrgWVi3XUuroFVDB5L8QWr1NZySabym87z29LY4zMfLjdPS382Zj1GI
IuTLOiguUGgVBqGOQYlXpHgPWkoL+hVxnghQFTPUnJ5Bl+h9vZ2KIwiXuebTvZix
azi8hE9xwJfzrQawXXygtphj9Lx/xy9y6fIQ9PfOk1m8kZP3t7VYsNlj2zKU5GGp
4yRK8ELU8/3cPVpnMpkc7k28SEpzO1HWaMtN1aoAtwY4LsvX0rDSCaBf4gAZBho7
n3MXqnPAn7xdPpjiBUslEBUhp5+LlbW2U2WGdNsabFcQOUndKhqr/NBO6sF1vLA0
UOlxY40iJU6bSrCeKyyrwK7OTCg7kh/Sx7pGNMVUK4gwt1QylxhwSz4pJKw8S0xw
lDybyA7sTvWzN2Kzu+oxwz+TWTxM5SNOF95vpbENWOEWaC9h0Q6vn7dudryRLI22
2WmTiUU4xjw1iWRv61iJhh0jjK/4neUVwr1/5QMACsM6IyuX4wfU/vOQ1yqeFXFU
8or1Cc5Rt0yta0Iz3LX1Wob6THUCm2ACR070SyK6E7EtClV1qM6iStaKKkOkftaw
vXwxBLTtqZ4dGS/VTDmaQyJ+Wx6pd3i22BykQIU3rlN0oVTDq5geOibxn/DQwqk7
JocLH/bSNEYrUnCooHbLQ+7U3vGTvEjT9hRp8Leh49VKiXeZ1Ie6ifxBVgGnmp0z
2RyoEl6H+jeMs1F+E0kElLbgXq8/gM3u8y4+nXT3QVY/+7pnLdyCzOVY5BJpbPE0
PdntJpLLCgJJsH1FRlLC2PC+sGVoxaVx4ZbOsOu1TLSLPRjD3ZClsdUNodyPTMCk
PZjMvlF++1R6yYwcTXCcT9qAlkdQAJ2iaqZLLqgEaTcUtlciTntL1CTnQoWIwAeO
CtcpDs2mjH2NMifNHtIsUb6Y7apClGdLvP70XBSdwjx59BDx6ArmAJDi49LQ4Y6Q
/pehix2dztvKq0srMe56tidHmEIbo/7CFNofGdat3PfgaNVvIGWAZidditgOsj7+
CYyfODYiqJtZQQRVnteSEofY/FmzN2dVPwM1ZhgwWP3gOicW2GkO6iaXhltTAnbu
6nIZznBxN96T8+pYa++kKpTYoedXKeikCexG0fAS676fiv02xa4phUDzGsH98RzD
5p/eLC6I40ac99OgEEHayJ5DoI4/2PUOrq5YSVNhB7o6pbzBmzq4EgPf+rVRobxC
XbeVYJ0AeanFPTAeiEiTUYsOFs/o0kvZVVP1E+cfN+BLzKSDkwn+Q9MDoXDYCViB
ySKHFDJdWdKFCt8u+L9GSldh2khsLf3Q8L/S/bVOp+/wdP/WQrp91scBQzs1w39h
lqYYAx6+BEU+AjvataHtezwnwyX4w7KcEIku5o03eYkSw/g9m3wWTeIUxc5hlbhu
xxSDb+Tv3KUBRIdU3LV/WIv9HzZVkvyYX4N952mrZAEhiY62PZMM9wjlole+8MxT
ZgU/GbEO1HVDb6pE3uqnRtvYQgv0p3G/ZdGfO1FQUQgZbJ8gybr6c9V/U040ybdO
eye8ZR+Pi30aVrCzpmgcnINW3qPqCKGS4TZx7TYnmYB1g76VDmrUtfRC3GgXudEr
WWdV7bKJnWef+hvQh2mWB62Rcz4TKMA2/MJyMlv185ReRlbQdAAoe+GOz5f8P+Qq
MovZOBtd0szGKkwkwjahs1qmypL3AhrOO2Qhwujj9kgXqr9Fr2CWiqRBd6qizU0O
2KWN0vcAjIdcykGxXsp06nF4SI0cRUkKFsMfOub4ELd4zg7DDcOU5d8Q04KkmAUB
H2Fx8Ru837uEug4vpGu8Pz1MQ3Tv6Zv0lFiz4GL7ycsRz5YKeP0k1HvVCMxaDdBS
67K0WkCknz5s5+R4nYZaDxt4hqmoX7hH3QC7IsLWw5dSWdk1MFj0+v7lJR1OjxlF
uS9kM829/m4cjYXnotY2EMkJ0kE3csrSq8vydiwAcyih4frGQYqLzDg5qMcVvlyK
aalDna2pb5wAnFYRTt/KiHS6wYaGVScr6C9+b69wofoYahW03X+lfzIpD2xK8Qr8
XdxxBQ6fH/MKSbQCI+5x6RgrVrY5FmQVbB/gUXbuaUv2ss1qy+QuhRMN5z8eXCAs
45OemkcRnVx7uky9pail2KStTmPYKt2g1bkTafKVM6tuG3xUvc3yw079Fw8SazTF
VmgvcejAIRg+rLtb0S0amoNFG1UGH3RjchfkU/mDt3IsAD1+EY4PKGhp7gzxWCwZ
gFanNOn0qgz8EdIsL4lcbpJrCO2WY9u8eacy/WM4POcguD0ZFgsdVX0R63KsyYiN
JnyThZW9SOwx3VVH2hNafl4gljfKaRMfqHMuQOp4wBIwucl5LMiE6GTYLulk0Xet
amykZmUB7hanP3BIrlP8iy99Y6Fp9VCjslpcAdhS1ZrTSitLXok3IYPbutiy+GC3
DwWEsLMvvwWybojsg97KTcbM6kfpcmUuKarCIsYk3ccJRYULwisw1UI+cXewjBfx
NS9ZDfxIA0x9AnJNu+G/+jJLhnc4YI5w5aQbgvc6XuvF+7K/QeBHUI4lvoC4lo/5
8UNUxj1an0tQ2e/e573YTpxHWH0JZJQETb/Tg+ll0hTur8jzm0518vd+FVAkmiJx
3TGyYFxN3K0tQtT7LobKQRKs+n/vNpftnrAy6ddPCMn8ZRb4pUyPZTGDTvoNhiI+
2UPGK/hWGV8C53O7irFMDwv1A+iil4SCaaXgtaj2kO2GzFlbL/yCFgufrZlxHI0x
/OLiPzKaX5RLyzGPo3+ibNm9bKyPXXzAtpOLgR98OeNTrIqLkrPqtKEF+hvRoNHx
JsPYNNbE14NOc2bgkRn9GOVSt53Kao40ZvZ+DBIofvFKyB4dg41o0uVw/jyLDrOy
dahMszaCHcZ9WAhhFoft41kecKL67ZIVaUsD8NLRvsOFs9jsTi2EUUMbex67EtLz
E8g+RZm36MI/dXEDUYWvM4qOjlFnW+FPuiwO4vcT/lt7KizPJ/nVKBAzZED8KAsJ
Cx7wGt5OnS7aglQCfMd1uLV/U8xlreG1LOCyY8eTU8IPp+vOfslJxhsAJXKGzvvM
uVmpcIv7b4ZthiJZ4+YRXTWOYXSeiJ+APyZhgF54iSlssAuNqk3PUCEw+ItKrkKI
y/DsrZdG4p7Q0i4fWnJZlVyugRJhngorfJCfPiXxsrWb/YpTzBqy5VdTR8+UNbFF
k2vyHNPi909FZTBtf6TkLPB57iPYr9WjvfZVMGhp3PSrIF7upV4L+9F5MsTsrPxz
oBH+DLOOWmHPllrZ7XUgugeycqH32W/oGJiLaqCos5ZRhp1YdmuNbizLoZrws8nX
mGpVuVK0bQPIe5unXfpbhk+B0YvmfmzF5FjTceQclCh+VzahGzM75o+710gViqga
s5qWa3HM6932Vl3Dy3DM0hUY0iUxFjPcOzI/Lt9ofC8nkn0yOQlCHPkSmnxEgK9y
bu1T0+GA2V3c31J4dFuE1CEoV07bQmlhYM8r5BQ0kwQgx7t82b6cyCD30oMzZE6E
GNcmRmQ38ewi2uyiF1yoaI0gaiYL6Az9VApYCSkZ3CAQEcU0BggxNMrpZJZ7UpYL
50zeTxkTBjXcUlEPIpdjvXqEUWygMXbN2pyr9obw1mcFxjS2VIysLUnf5aHqkaVN
MJnJlj76roBXMmdqfL/ls7W/VzN2+dfixfqr5bmvSFQi/c/dn6kQPj1GF1RSn7nj
btqRPSvevk8GHrbXiRR0zVBOPgmcDjRAaFr+y2uA+Xf+QRpwEJWN8cXuEqo9s8Di
64QoXsEZx+Jr22ktvR0jAq2X6KFtt+xUPIUYULbfdI0T51OcxWQsmNgvQPsound8
neRZ8+Q5Dek8eyb+rMK597atTYcbeKe0ianOWgqb9wjd2OhQzqvjQeR/TPTAHg8t
CGAbiU5RIhNL3U6qAUjNGcgC/HDRtbeUBB+YFDGMFpV68vx3ohJJaZjRKSW4Vx8w
GWZ7mwM27iuMbhsXkEYMuG3n7nRRxrImZfn473xvMqwhSByp6fyajUzavjhPj1i2
17nfkbZquutNgPWDDZ7y5eqMaEi01vH1lq7Q1yBXwIynqtTbInbIJNylaJ6Vd8US
8WTD9r2Fwb4Sq9xou/yoPA1HlX0AMuKGCrGDouJzfteuZ3VPaGcI1HpUh8s27J62
ahjbqiRoFZOhs7HYGa+fvXPDTOltBzXFAoyyqTpNdHo0gArXpl++HtnlRccTfJt/
a3TeRj6KHmZbhR4+LF0XarBv60j1E1zzBDHuHnDzMuScRN0arVfHR+XbwgHrgg0J
L123oY8YZhocTCAXtLeP35gGWpG6exbYKNc2bAJkchlTbag6SR+Jiq42Mj1SrRUX
qNgl3pSOind6ICsC/Cz5ei9SsBnc11k9kpm3mPZ5nq6CDj+iYgfsX/UezOLNVTOG
lcXfB8O3BEfAc69scX/zK86fzxyR7uzO4FppleW31+ZAXZNxypQ15ZptKBBKsbFZ
9HF5DQzB9H/PfdUD9R2sirgAYnZ8o2LxsoMcpOjPiBPfl9byQDKaj362ikZXCe12
LrzdPB6oAOV8MunolsWUrsMyOT5L3nMEf2/hUnNh4YGBI5djyJXCTAFoqCJM1iHK
c2zpnydpDQoL0OjELP8Ixqm93J+tSRW3Hr7+xVXQeqYvRpXFExQlKH1huqkv8Qm6
2TizQ40xWeufjQd8FEqOXtOcBMaszVJpXkBp8Q/AR8Sw9ckgwNaAX7shZx0fqs6r
wwUAtJVLm0wTzktzGv49Zi9Rq2NjDV89WfmrIMLBB9MVqm7vuwbadPN5fJjH3HxS
FVgGnmsfPrLDXmUmchTd9msWSSwnB9AF76IIBp35D3C+fedDVDt0+qXZtZdoC7oW
wKCJmFZ4SFdUojK5vFxOK+so4oGmCixRxGR9jBTOfLJXl166jbh/BPA8iqHudBSH
XRJc+ZV3VZA24pUGaXzx577i1mbzqtFx1fDjUiTCCgxzHFQr1dv+W9K6Gy3JxB9R
WGnWlsrI9dSBZtZiUvvDNqRHjN69LO1L4F7VVj7hrfXzHas/4cUNoOEZl5IEThOZ
ddR4pJD4ar2ZvIkrLsJQM4LtS6D712SWKwOAQ+l8cDWQjS6AlV41aKCAJFDr85ks
Xo5V4cuzdDruyjRiEPkqEnChMU1exRSV5EW5fpBSdvjxOAva5hNjeQr8BYWpwQFI
0l7Xen1ntGEWzg5A83E+c0wFbEz1K7lnsoqGiUkYL43IEInJHvOrocsoQ43chemS
4L8SKLZ5Ztmb+zW17DtKi6ArWpQQhCkq/+Sto9CMzvyJ/Yeu44EhCpOUXl7sXp7U
hWCvgwAe2rwemSlkjwWjSRwzmCxgejhn2kBsIr1EBw0WxqgsOdoAyAaDJlNI/ISu
tp5xnA0ZU+ZSMDJ5x4n+jLw4mg4khd7SlveDQbk+RrrMIq76Zt2ekNVzt3B9cYte
FxLiTk4QF+2O3zjxSGLBOZNcwt4y4ZgF7YEk/XN+uJwWb3wuJoA1d47S9fvBHQVo
B64eHINeylOV/gKRd678snO/MD6bPl/1rAAvEtR24HeBetP0YH8vsWBx/EDNHmMe
JOKxmifPI54j/AvMclYVxndGSx8M2QD91BFFeAOLww3/LAp+GzDszkMJ7E2sXDHv
doEht9YiQVCvgCHbS7wPEmUdbstO/QguC1E8FDX/OrSXR/4Xy2VVTgyumFXYhlU1
4ghM9qAHIbQsji0ZxCKh/XUPtGXKK2PjZ0cH5xzkwzVolnQ9HyFzcSJNSBTp1qco
+L+D0oELLpWH/l05gEesLL8XLhnG3zfSDQPrfQuJnptVdtzxmif5Nga7iLhyyQTx
zAAAbR3PzQ/5a+u3p99p4QTxfErREA9Yc9bGBF6sEVstNvz9yAaPU44zq6wh8Kod
CSLm+vYNFUyfB83Cnvy3DvMechXopVLCNrtMOZJ2rFulEOlMTomTG4bEyQAgdkN9
/FSNZbeRJM2hTDLZoGohCrJ3rddSs+U1CeIcR1euWdYXDuwm/InB83+oBiM8hBww
qIkQGZXUYpFRhLp9gZS3UX+sU/m0WuLWVrauRqCWS4JIvUE4WwvJHUZcd0xiWV6c
x+Cgcm0opj2ewKDveKo1iO+HgU3zpOo84GFkF44OJXU7t2cOzdyKy79sPjtFdZ96
IyBynM2RU9oSAtyXs9j+yXCNh9aeuZx/gSnvboe7g7HRwqwqz1HZ/7bN4h2oH9Ju
TX1tC1DVNlx/2NfOaYca6JkGKeivQ2robaVDihzFN1+dGXyhKR4JiaDXx4o15S+R
PbbR+v/mSg8OK7zTO3UDajE5mOIK3IKKR+N2hLnIvnsRAGWXz/BgsnrkU1GGdWEJ
Zy6SkJ+9Pzt9nd9glC05IKmHISgj8AXYM9/fff6TARzBtKIG78YxYgJnZzGoEJfw
KVbbfpimIeJb8NCetHW1SZ0irz29x2i8czOQ5bSFrkeeCLSeR2Tug5MWCvWy5Yzb
wRqwEvnZ+aZB+qlEMFVKs8GybLCQMjh8fb7yzyQp5SqVLHWzipGjOezoHTkuv6PP
JC/sUzwCW8p5LoFlYH/2GpXwZ9Gqn0fXetcMRszRnkK0Vu1AIyjdP0u8C23NQ1gG
jHfcTP1kBwQHGHTIkjXjhk4BNSxI1Q1ncFdRjwTccAYkaI0vRqGsKPaLYUVnf+ER
8ZNUUauqcz1STvaXcK11OJiGHef35JdjeOJl32q7KfJXc+NoMBYlZ5MYL9ZDmH3b
3xC8XAdkAeUZkxLXIVVerFF8bqUiWw5sJSsYskKswEsFfoBxoUCaSgrEi6QhoBX7
YRkP/0dmdIdiP3NHmOb58i9W+buDivnIyfX/aTdNuSVKuWu/dX4+TLngfoe4Tbey
7MOX+UbyybJcpvGc546cSpuGBLJnFvXNz5NMwq02H5uBfptDW3CS/8J/zBp6+4xM
xJ6NGzA7txsruFlCuRl4ZxyxmSegJcM35MwaMsoD0O62AU/kGUX/Gl2vqYtmaaUf
1LDzItVV9/FIknRQZ1EgPjU6CUsPrUz/yb6LUFgvlWZeB6hoENbg77iL1yQrqU6y
wR5HNJvukLCekk9IpgRBidQKoWTAnTRc1/K1wAiR3wsIVdWsQmyulV1cYgMGJRRX
J+lAX6MhE4oNhOzX3RFI7vEMcdtXkcCiJKS1+6fkM6W5Wz/hWpr4OggyLmiC5oDd
p1FTWNaViQ1OnEh5et6bdRFHprOc28mzls6yxK7qUVfPOE+UCBgZpblhtgqqNDs0
Td8VchpwlTsyhfwylMLmilN1ew5G5ChaQ9kfS/Dx1pGzyNilprF/5R88TgTZgtmx
OhVdZIzezPTHnl3e6gjvqNeI1Z24Vao8EX7IqZqTfpi99ROj31G+sRLjdMXPOP+P
8NEBaMxCZD0/DDCC5EwuQOTyxIg+G4WTEkaPl/O29oM8fs/TaFKx06Ctcz5O01mH
OQVqFFeQJftK4UaDjj0lciL0IyTdyhJ2tXtcNiZbuDb9bR7Ztn0EvIUEmqLPQHY7
oosyyvphEB1HRh6NZIK7RgHjJMnZCaSlaE1yoWN2HfPpK0NggRSuWiVBPTDYegHd
lOlmbEaQDgPxeTOPiDv9QBhhQBXaRUpQBzpyBOpWEJsCydnPjIsFtf21W7J2p5qq
ohWLIp2mKfA5c3S4FbW3474kKIH5z3cmMlgwFXyYsd+Em/mK4p08j2mb1aq+8+xR
BQYObGDKWEg5OkWTAknEvv2PHiP0NMFCFypULmrIs3icKeZGsgeUJSzC8ChY8P+x
NL4/fTiIl8drf53/kABIPrCPY2l+hz+bUXf7b0MD4SUQYqumVE5cABZ8bee4mGwW
Qpft3HPr+PczgHOUaHbnaP/UuNCKKp12W0BjH1ZsvdRcmaLvoTAetqn3LhZuKl4T
S+QRC958WlT8lB6/4rr6dM3k+SNdbgqEtQc8dDwhCYed6cHK0exf3SKajtSvktBA
nhhgKgOrTKOnDGn+QMCRruB5e2Lx9SfOO66Ab7ZiRMm0yjykskhD0NTykMC759gC
K984IkKOBLSivyKD2KtC6NSsDsoJpFjiM0SgOg3wfEr5B9obh00CY7fV1jUE65J1
S0TA9G7Ie1ED9lA4yN07CH8XR8Zf6M1DZA9nAhBSn2I96hxdLlAvrNaawDc+mSky
k1rSx1S/1ANB5ef3vMGXYvyuU403KudK6XL2DULyfzS64mTbzBt45eaHZhmtcXz9
dYXAE2kj7VBsK0fwkod5Y1Pk6GGZuFJV1i15bhaE5HYWm2Hsq4fSgclDMbjMz/W7
Y7qWUjB4Z+htNwWWoW26uwZt00qI3tbgCwRNlYD1lRia33+jvmgL8NY7N4lrxoMK
xA5qtI7iX3UzC/elEguI/Ddv/ZxkRftPb3Hhe28yebD70sQ4Obz980r+SCREEdxs
nzjjaXfcehDhwtL7Ostg6uAGkL60AwM1rNN58gIcO9LMSDA/em4vIYx2iyw6vgoj
veOYnOqQ/4hdaFCSbNVea3expllP/SDHlfrmg4419/eoDoeFwkjE/9kcr4tcA2ly
VwOyd6Bk/ZlpXoGls1PiBylo2HDjR+2ZdBdhWy+Re91hhV8tzlT7hiD6b6wR4m2R
hExLBu0I1An+NhITA6hPLHMwtSOIyDLynOzlr7wMjbbRlQ4cIzBQiF3yon9os7I3
MwItvFVEyQ2kTfJ/310LbHk3vz8MiV+XRoE2EJ3xDQ9gz5FlkoRlak1yY08wRxD4
EO68GdxGNFcEXSU/KUK21PwZYfE5SthFgfW26WOtPRGykddH36gVtKwO6cFMf5q/
1WZUh7EnFqNwBxeanagOnYNSrKr2PopxZGKDCXoTG/r07LC0anqhzvyZRJXR35d1
Ky19CfyR5ljH2KnPcOEVTTg405ryULGvSQsbNt05B5zoXH/YZd1g1XtRfMzVWmx0
sTKzPWirKJe/c7NgTFtq43Pwdvxa3pMPLyn7VgtYKv0kMPGj6wH+HhyTAg7EATBe
iRiXNAQKrFRkcK6650Qtt6i2+O147SUskGy87u9YoLDLlmL01TO2iVDyBXeWIJT/
FVMFmGKFWCAXGLecOQFCPEtxowaAlGbpV8S1MMuSJ2FFxSjkp4W/Q9B30B4RmLGu
ZcD5v9ZedeIEg5AjjnAroaBeIA0ZuDxn611zo94npFmkybnsFoBnXl6E/NjXNVY1
ADAsn3A5TQClpX1C7tniDgEHRougx4rhD00dA7Tv+q9wBdQONvgFjWDrR8jmjvIK
JYAIHTwAcuAAxC6Fy7j6lV5zUtB8+olmFfDODE/5lUcJLYkJq/QFci4G4dUr2cPC
z3Djy06RbD0KuuDePR2gdRwoSKzXnbS+vNwwE2AK1kKQOYtxx2wU4sCAL9U6Vj/H
h86msmKmwJ/+e/bj7lya1fV9Z9VoKG4l57XWmppY2QyFkfFkg32+iV+aG3KwKQ1q
aljSHbJY5XMNCvZtD8udr2iZ+bRJi5pN1N+aT5Aag3tZ0tJJiKfHgySeoSRB3Iun
k9LTLvRkk0M6xZnarkHDf+y5m903sV4LWT8obgmYNdBHee4VAfzadtm9q/qM6Jd0
bVCkOg71c2wrSjBJYEX4eX/2bg+hMHBtDmZ+fL9SJuMQrpDLx3v7boER3YorrnuA
9cNI8bERAKJ7SrKaefvQfLiEFXOkknZPdTz/ouDcbHdiQGDRZnPWvsM/LIhyrY7D
5DQdms02683oBnXqYU8LOJC0v6GqZr6vLcVR71/AKFdOoRtIYxWckMNHffL8az2/
IkAmH0HOp4mQomkJAsBgn25zr0cAC3tq38E0qzXsM98+Ni5Y22ntOTpGHN+UlA0C
qtJjMG4o7i1+iKzIgmLGI355yO6SdA2DwjDB6CPsWCX04vsCqF/jqgzPU4/iPU2C
DDBQuFcAjrxSsPDWQF76YfJDp+gQd6vuThgLL+Kn4WMaNVNb+oVqe9X80rPSGtmF
kDlfQxFWguKkGujfO3ZKnSLZeygOphuQLVZZw3ZYZC1jGrTDmeDOZJBwXKjxOz18
iWohkrYrjQsK0N1w440IU1Ch4I+R30yYpBPsOWdlJ3QOWCJ/9ZbXX9NkevY5APP2
XudiyceuVT/A8As2e7k/9i80Nsi6v/BzKqw8KXw60kjh6ifq67slrqIouCnEF+Fw
awkh+YJqhih+Ct5IK+nAM0veXa/cS3+8l4yzjO0uWagwcQ8ztxiHSbqilfIuEESi
I6WhVfcwy69DSByH3sIxM0Na7KInOo1+QJbITqp0IGHJS2aaqCnM+FSlb3otViY+
QvIlZayn+2vEZvErOWEAvqAHQH8qrzIlC7Wh254EPGsbEBmSFrog83TjOjEb23dN
ww82unXXoo5VGmISLuc4HMohAOpeYi+EUKq00cpZfTYYsxztlfwYu0W6icGmp9Vi
fjtwhip+/uyfQYzRkeAP7vDA3Hr7WIxXWR0+RjyOgslWcuV/jN/g5bgncAchoBPe
mOUHPaYTBJUy02JmSXS7nI5S2MJPcTNdB8VOSgDY+6SZc6cVG06AZ1SoMdwpndqE
4yK7+vIifDX73AyMLrA2G0E/sGvpNQS77PaZ6C/Wc8lK1cL5ZMkG8+f6barQOLeI
ZV+ytDF44S/hpUbO5SCeHExpeBPXc6ac+L3tvTUC9n7ozHfD0TSwb/uTTvu+r/QP
Kr0tLjZxJi0bTrRbAara//Hp7mwRVTQhgUF7NwU7qgyFrbCI3IM2UPmJBKQ3sfkF
IBSt6Of/5SssBQZVQ97wqxEcBfKmtX2V7BfTnHaDwbABhr50hBM/6eeT+hcARA7o
VrKqJhQ2YCvOH2M8Q864/tco7yzIOjgcOwtuMmAI6ExSHkWFABDIiD5j91gK36ik
ZnGZDcd0e0OvhUI1JYNn2jUuYvizmW/zOI7Wq4VIgpeQsghDq6d0Fg1sXw9JTSRO
cFdYAGQOr28BuF4CL4lr9+VbdejELLueNvBgBBmaoWPKW5NaZeCZ6N+329FsN6pc
vX8Kv0P1HdQ4iuGiDM8NGiEWjom+mOTK6FC7suim60ERboFJ5ubklsE0lfOXoOis
04IoPMzDdR+unCFv6+1izp2nmji2W68P0GJauHc+SM53WvVFw3MSFkDWTwLbEnet
KuJXLduK9rlgJpXiRfEtavGE4YKl+SBDuqXohjdJL7PE3EUxWIfiOgVuNQ4ZpkMy
/g9r1nF01JonMq0cc1tZq05nVvUdVxQxT3RQAbz/pjA7pjdMJEMP8B00h2AErOUm
Dlm/uULSZVkR87PjI5Lbv2pStKGfDAtFmPv8pkE3I9gvbx10NN6d2EH5fVFF9/vM
cCgWOQ7A7x/BROuZ1kBmWuITZEOlg9VeGa4M7otEjQGc2C8erVt3SGmYaK4vYatS
dJYx3F1RqbTsNh+Ug0h/5voBKNHOFdhaafk/kLErbHZU8+QvIgFHG7LZdnAv1ddC
st0EFfknP2h8oX5TKoNEfI/O8WcJBs6Q2a8ccj2suNQtg9RqNGEbMjVt120u7gzL
EdLbyaD9baXSKCKx+SmGMTIyZPQTjyR4i+T/QYXQpf6Pki5UVFwP2hNgW9u2TilW
yRaAEaRHx1cZJE9rARUAIpDqNJR45EQ+05ZtmN9iqt277nUWIyxcBaQntCljs6wK
Q05UT6ks2d/xoZSfWAOl/pf8dkoMBAIJd4KoFSZI9D2YY2GWXx35EuL1f/vZPLu6
ct+64GdXJ9WpFWSuNw2tKHQLcm5as5Xj9Fi7yDbdheIlw2vd5Dh6FUn2zlCgsWV5
2NbYnw2c4yKeHa+ixELttNoHQlR0bM9lW+6zSQOhMlVnotfFGHH5eObD1YJTM//x
msg2uc2QoMwk2P9ZNe7eTZnQuACKnGXA8b7ZHPDwSJr2VDNLOTBB7y7pM7ZiOIVm
u+RfgK14+cz/e40sO5PnuUWD3SeC3VOGM7jTUPXh6QRghT2ENTteMPNIRYPhV6b2
s6F/uIZGTGPPdJKwi9wAqY1nH4tMzd6I4PKcXVtuflq1NVnybltpzTJr7jJIhYSX
ysZKnYGyi6AccAl92T1j1FPh9sCeRGRki5vkreaefW1Idd5vM2J9d1aRBxDVJxD9
4+eAUSrftgniJ2z0kqqJEKsdY3UgtfsAM2rVQK7iEpefcn8ETQMScowrDZHi/jAv
mYABW6DeZl6rkOidwBh+ZPFlYdU7+Fbyhhe4o43dGuORY7YmPCHFY8bjmJei/i5k
vxr/ygS6948SV6eS1puSaXPjKNWwGo2bGvZQEvOS1FVUpRqZp/ZDpEZgNN5MrycC
YjyUglu14g0Ja3ZT+Uth3UcCrLK9Zbq+mYB29c5OQs86/OHka/arxj0TV3JN/qzo
7Uy0Io7QYpyTVJ/9asbUMU5v7lQd0s9veCzXiFyXfcE8sdPnUuWgc03idqbI94Ow
3/A9KtXhgTelsChtHeE7zj5B/ts6qZieFpJGvVEAFZz6wSziB2zFdrdm5Qjg86JA
KdqrlIQ7b7KwHvMn4TlHvvaCfa5gYSoOglMdkNtU5EqfT+77psxIXnp/HnRhRsqj
/VXhADAzUdoy8BmAd/nNfeLjAP2hRiObf77Ez+LCukaQvuf59yXDMWRPCteNNuCp
bYbqvz+zvf0xNQyTFQgcwkzLVXSy80E6b+At6P3jRjQIZ7iXl/Z2eFaFasolIMXM
/C1duSu8B1gusblVueLPirEtCiXGOxcE1oUqcCNkkfCY3/bKJVMuQxjTDFsdz+qg
7axPDS4lxsveqNDkSoO9xdM9jVte8GLL1P+/yultsYg/6wxdVInslk54AGqPG0Gt
Y3xwwAnyuDFC4fFLpknBFGL+5zN5Tr5M1CRjBnJTsH2aWFWo1I08hk4JiyqmlaBN
5hWnJ2Z7ykwH6pqnAJG7ZMokYalVlXmE1WBg9LgMqsO4gsenop6MsAflY3oPIGrb
m5Ax6AeGlHanN1ZO6qBDBEGZpitKM28HCJ6JEjtJCi7ai3pUeOyIC/CA52D9JZuc
dZTR+9LC6wa4uocydXmKqvh45Z/WZA6dtQ3z5WYofWRuCi4rZzvxzm8ByC414NUZ
jxPNMgbq7xlj+IHXlSi+p1btAUQhtCY7tyF/xfGWkN7TfR0VObrF8zwN7pceBNfj
yc2aINCotyXbRKtJ5oTNzK7hXdGW2GmmEmZs5G0XeTvHel+qLlIDAy3jnc05Fu5P
qEL9GOksqEfE2geuMIr6vbKroRopvKT2WuAlezSkHbjQqyjW66xwa9rlxWgqNEmY
etRH8Z/1+K3dU2RygW3cQ8LuaUZVZwhgrRhGNU42IKaShX03CAtq8whT4c2xVAxR
E1Hy5Pv1IpBLgK2x8bxGdjVuMLu4E8qwvSPujDc6nFnz7QyKbSnt0SMDWf5Jd9im
f7uhlroBI9AsuOKLQGUm4S82TLWoaXUDH8w1xnKJJNbShM3Homy+EiHO7yuokC/z
yjSO6TVjE09ekVKQZL4l180zHytPRT1pBaYKkvUUWED+7ZXv77kU7MSs6AH61GJe
jsDt+KLy3hXLzpWaRCRkYf3263RgsX3+TSiPI4vav++KZjDIVFFx3hzuLZvc76q0
7XT7dBVIOu5Vn3BHnjKMelX7+l/0KFG80NSmm1/fkvj7rEOhKCrwN35rLOUkw1+L
FUBaD4VDPuSY16U0wXkYJ3XqwGcDTd8NS09Dz4bEw4SALUZzsGz2qpAPcSF7GpZj
2gfqyEpYS0+B07wyd7GBiDsFslh8NjoEejt0RyzwhpXrtkre2BlY2aquQimun87z
WlL3EunsDvVqbI3IQ4Sl5J2z0sCBQ2foTR3YBatQNpsO0JglxBuFv/R2SgvSKVOL
U7l3kJ1uLblrQwiOSrTDHk0uQSDpL7Gjd9UCrQvvjDmg7yhFXJCP1FpjnEuUGSfm
WZfme2YLfJkG3yfXwVYlegKsz3AfAD0LjRQuRc6nJyT5kDYTtXj4/TEQAJLB/ByM
2+5UhspfEC0QJveSGVH+V4Pp9OQNpl4pb6gsja9v1/57r8cPiMIDKS3GjgYgUn5w
9voybsTtbsFEno9AY2G5MVmh/1SXHJMa5BOL8ieztkWgJfNtQBOFnBYFPIfFrFAP
1a+BmQyPgqcLADb6SpK0+Ru1sUT4UUnZMgRnCFQpI04/+UOxio2PeZlikP7yvSdT
uw4xlMJZCawjpRQubU1FyJZTUZJm+6+Wje5Wdw06XJ/scTXleRyUIqaG390QTTex
63f8YHu145r4uErLXvY7Jy4CcaNsxYWd8xGg/tkzE4Mv0MqaL27lthCH+vuuhVzD
kZQrf0TtNWRYHwRll3sV3bNs4wbNtu/giv63Nw3gangPxi90zjMlnLR06/QO8ZkM
iPSW3GF0VmmDUgkmUl7S1qHtLo9vKqK3Lzxyw6opbmz6EMz8Yu2FXb5t5KpsI0zd
1pw9S/+6SPzQNDECnssEhVyM+iKk9HCirCuPIqAfl7m/oW/gx/vXGtHZYTy7cxza
l8jVbbVv+WYdogtoIu+trbPJBIEtpneFWH7cVXiJ06teE176LPgxpTQ8ZhW38dl+
HhaGvYQqpisw8QAinWobUFFfvQb5GOdM1dBSeECBJA758yvRU9VhiCbB8Zag7Q+x
TeyHsOb40bxGpGOidB2Mo9jo7L66oqm5wEu/aG0qX4EM+Bx2baUbqNj52WngY+tV
LSX394ajHjY87K6XwwlZ6Xq100+w6eUYH/w7A2owcpSmLpaFCYzKh9KTT/ocYaAD
86CqFy2m3hsYOLZ3zwTL+zhYx3EEteBvTpqAU2gl4vF5lDWxpE3AKtUwrGQut8h1
CWMScKoLGn+YuDz0nzKnOOei88XoL8+7WDBSVXaSnMkVUhOXz3cWdADEvtNrTk7f
jU6IP9/sEpKzsZDjvAcO2WfMO/OM17kse+3v/IyhvWleWRvVhpR/xvYCcBZYYUSu
NL6Qq6btCnP0aKON3R0v52krQhyO6UcCBrMjS4TeqZIUnSDsF2NqCNPYeRKDHJiW
UPClo6jzpRNE9yDFOwnAZZAP/fU9zes5QdcK8GmOHPxP3PwU5pnWFbrAYv4+6g7v
CbclGNlef2LiUr2ItMpGY7cUIROVeJMlWRI3wswptBaCgYslMzFe8JGF4ascrqVz
RRyngk4ARM07ZVhBsGbSUg+hlBiLvtSE5A2eSEgL93TMrXpbBSsUWs7lbrkMS9G7
oYE/BFa8O1XmIEOWI2TKrSnnqMzJrGXssILqguLdWcKfmwwL+SHXO/wvllHFpPwO
KQGzaEKcyfenW8DU0Jl6wa5sqL7ZVCY6jdeMI+lcvZYntmcx5WYSvysdJHp09ZYr
WteBGKaINC/aS0O1+7A0//z7acNx95NXv2t1snRUTDvtm1in8HUkIiOkt0SkQlgA
fcqheTeDNHvLw5iwNzk4V0Ex9rkhuY9iVGKaKH7t/OWTdFZghXmqquPBDVVZNebn
0cd+FhDhkQPMVuqyOZL3pOJNr57onBpCefBim0JcpKWtseOoD37IA/D2T9x9mEOj
tIWscdJiHO949miM93Zf7INnFLqqpPaRqSXk9yry6c6DDhgnTgdBwbnlQDnQjz64
UHncVQhtU63yUnEvK1ZhrK+fpJDJcvspNA8EitUeERVjQSGvD6EH1B4atjlDNExr
ZPT3S0mYGWjjUihi92CD26qBXGuTx2b+cBRYa4GkhqPa2jFddJOoHmiXywdxDJCa
SuuDi51DtEcHsaoZ078+fTo1VrBT91U+GbGaoGAC0Mc6yvnQCEfqXA8Tr/2sNmiR
4B6+dzM+0x8XHsJfEikl4Hk+jxZBAiBrNXvOrj22DCU4EvzMKgrrTkz22SOK3b+p
JpU3LfgATJHIx4IoGBeZkn74wq7953zdwlqn+S51VDUtdT+Palazr1Dwr4pDGobH
qOkTJG+Nja63uOjKXFuuEfzk7C8qxotLWbnGyGyeznGHMhgl1Wfzmkhwqbk78Tlk
W3d1F1a+al/Hqd3XpYD5jXdbLi9OaDCyO0zDT56YcDvdT4yrpln7s45MsZPFsRhV
Z3e5L1Px9Y78JUjHKucGTjHDYFQ6mIbDovVXxUtxPPbbncId/lxKhGnLFovhn2Uf
2OGtNbFRQdZrNGa8tkQHohmqyzNzO+FO8ZkjFHeRc0o8dooKVgUElQf5gbyM2HzB
7Gr8IAUKioQltFYlZYNiqYdxcydQ02REUTzpcf6GDKWtO+EQO7CEtliAxDiL+AQ8
CVTPXZxiHB4IzpzczNNrsI+kxUzig60qhhPFRJFWkdmWUOT5Az6EvZarb4NP/czQ
SGw7EQhuGOVrOHXRKn8TVLQI/GQlcBLcvUrKxD/Cndf1TwvSMN+LZMLkE7A7zq4v
RkU4f/1DD+ybBSqNWD458TPBvWW18E/JYnZOGLbeOIsqroAm2aNoCOjFkPf3VrLr
TF0s5AChkKyyfpSjyPcxWxhaQfqXtCrdAcI+6oE3l7Cd9LNllNaa6CZ524zjivm/
VDsZB6Xbxo7qRIM0tqaKNN7UjjaSo8DaNIYKkDtoKTVurlv95MvgWvmkd+ehMzAI
VmGtasUqB/l0AS/1PPYX9Q7JjYHPwGhjAsD/6xBRcskZep07Las25O0/RHvyRmpe
GGtYPSDnbGXyiTPvF4FX08+65QIeT5htWlpFWdXKZE+h97CmG1abHvfXa4UGlVPv
rJH3thOZIbvvEVeE5Gs6Am986Ohd9A/OZu6TfLpYqeE+irqM9hOaspwkRJ7JWTJz
6xPQ94kL3HIDz3tK+w6A7aqtSzDEVV1Of/jju0yEJmOJAdY7SVDxWGModL9QWbKL
/MrEvqUfkEeXFXmIAnIyS+hbYkZhRQpZL3/hQGuPhIA49q7Vt5gA9hYuUgQhPOFS
Bz65aIIKLbGuIoLHiPHKhACs6AcYbiHMrEDutXjdymW11tCopeWvau7WzvRQLT2S
5x2VQdd1tKe0C9YND7wlZsxJy98rn+M2lT1YovLJuLo0RXK7zbw4B8K1X4wFR0tP
c9/f0VCkr5Pdwak63SwSojGCiafA+EXF5HGUsWTsr33W1XvM5jsforqVTA4dBoxB
WsOsbfFvMFRYWGSYhrJzu+3KzJXnd6R2IVrmkql0Q278I7gAPn7euHcrzv4swRAJ
Nhz/p3XQo4aubx9nFjNIYVGpS2wo3LD5qxnVeHoZt9hrDYozZixzM0abYuJubsBr
L0Dvo7KK/NElRUrTgomRJZjvsPRRbcLwEGz/AlqRR8TE8ZKXTFt9dj2XfjVHVULi
Mlzl+vqfx2i1037kMCb/khrp8HPcW8XAKY4tqH4jpUEs3DQ56raItctYMz0QJv6W
XSCYVfRirz3VTL0LOr+V9NicXxJqm4suFQG4ugPo6VUkMZ57bCGMwI1d1kW90hDi
vp231FqRP7ccbTUzQyK9F6/Pgqh9WUO+PVY54u4evmXFRQ5iiSCmmcbiJWqvY6OE
3JIULx+qWQnFQzZ8rnq6nn5aveeAE8p0psDzEXUl826+XqsDw9UBfSQmyFGwodPJ
S5LuQeCFQ9Mr66jybHhRYTTx0wq/Svoo6QZPpf4Vco7Cl5rQa64hjpGtrU4ZbKT6
fjQQIw2HXNdmI2FUyu+Rniyjy+qn3Es3FAhQHHfqsrMN3iwCgYcWkjB+fvCseJB9
7DHun3670xyGOFE/BqrOzOThE3iFN4v7a+CKVoLW/NpVyy7QptJw6LSICdLIUZLh
wO78EY1dtV1ZM5zU3Z/wiPtTjbr712SRPyD/RP47uKLcrse4sTBeslSdAqO7WyxZ
p1OLmMKLYbQPg9K7LeQW6pk7/UJtFvvJuaOFb/9Lu+fKeGQ18KRB2PA7nZE5gqwM
3/xjLPRGrOQywYD6oWSCv1Ggtk6HQLX44tqI/WbDw9SHGkNKe/NmLv9f0NTq/SqI
szmiuzN5EnoOaCnEvEIMBtiF+C0sE93f1NNhAhAjvqz/XNIFPv4aL1lKQfAlkmyd
JrtWegLS2mkJVZEnkd2GydHJvLDVwLiZjBNiU+mVgLLPOtqcF0KFvvH+E88Tkljb
3tunm8+yN5xClPjDO9Ahop7MOSKD3XTeWKV/q2dd4X/zSVI2eK1whvGEZG3rO+cR
/lYOM+GNUyRkjruQQUY+ZQVKoBkDRqOYFbk0ki+e4ztSzW+77ocf9mR3Dtv2/KwM
kHns34YWecJuEgjTX0M/RKCZxG+UP0JzkYOVXuHp1aRuAcHeuTM3H0hjmEmpbeYz
EKjLjYAYJkikxCefGZympsx6U3R/lqEZotusHn6zIHgwnWx0jCc/zhlWfb0nu8gz
1rCKhrff6/vOJ2RR7oICou+miTGu76ug28DF5n8f5mvJNoLtrb4O5KOqbEJoNKvf
2It73P0CCJbUKV8G9241AXfMg5SUEoyTkCfD+z6uUrTUzmarmsGe7rjiT43n29gV
I9v9z5ZVRSL4V4mpUHh8UdYgJ6VNo84CFE5PUAgnFfe5LWBw+i9vDrxapeDiTku5
buFf2UOg43eULVTSqA82TgIKhdWCL67vLk1flGPJRcKe07BT9EVLsT0h52iIDfbQ
EThPTNoEcltXvkYAP8FRpHs8/cOisJJXZcCzzzh4cZ6PMtAvL4LdnsbkYhgEer/Z
O2EtmOheDExYqvTYtHFyBDVIezUH71W1Z9PNrydb+eE+UEJ5/bfIWkibsebc4vNY
lMvxZqq9AtGA/1Kq8qZw5Eqd5Qdglp8Xuse7GWEbylpf0R0Mg1FIoY0cgL3E3I62
D+i5fgAdhcYgGP0t/TWjgo3P2nD3i1Mj59JMErfTHX05wEvQY85ZRGDHHSyB19RX
G6vvaZxXXrYLialdm51d/KnS2CNSPpGqETM2elpqi2udwlPc8CT025M9IfS4eXVi
6nhokLoKWfCDf4ojVtH0TAcF2dX3ptA+C6EtWr3ZBxUPT52fXW3iBgjkGS+NzKrz
2mggXtwZ2/tVagsjffrjLmgB/YYT+IzgfKZ0VJ4T7VYaZBGFHMD/FIMSXRjC9q6Q
2QjK0TYIBZEVTdWHFHPY6UhURAMDxw4Jf2Sod3g1zcdZsBQmGemfaw3ojg5Ojv+7
6dCLePmAqvYjN9UsjbKjdTIBJeWX1iUuvPpB9dKonznYzTJ1pcOdbgOQQjErp7Vn
eT1LQ5buyHe2aEBemz9rFckAMqIJmB4yYmzj7rv66UCXOGUVMgyPNEs+pP8/FFIe
meHyfFxaW/ll7upYWVsiNFWsrCk6AWCg+KQ8vHPJBCF731ZkEtiMzkKZNqVS4Z+6
fbBhxIG3PssZIdO3+quPwn1wnyW1A4ehK9HrcDE3ojIFN0uwrDpMeGCTAvodSxsl
YQ3KdLKknV4HZdIahfj5TVl6oBfK9NX2H0HtwrJHnGcdM+Yx8reo2KEgRSCUw7/P
Dc1fBYvLzPqFyFUpU3nhsxjEMd7/cX6vyqiB6cmVLTGtaT/1Er9/xpBFWj56lSeW
XikDBHPz1I7uJJmbt1Ab2pLF57PQerek5Y1QgTKc+V45hh5bcZYTdE4rwQ3hZEKN
D2Mp88LYznWhuTH+OvT762AOGBqYIRDrPBqycSueexC0DXnEKN2VjZ/QHd0/2eWT
F69RiT+/FeM2z9MuWrbjDFdlBNtcWP1m+Xz9YL02L8JzvJzM9qHqs6cqtiS2ZYVb
Oq92AUgtTbHvo4yM8BhOMC5Q4H4TI8lkM70m2Yj+PSGlv7GTJhBXbWGbK1+vEC4h
kvmDfAOmf2zePdtrGK2O3vagGXLaWDzuZxAqBRnT7t5pC5frpjik9L7WptPm4whA
3GeScMga0IOemihnmdQMr1jhlIrwStJGZ3JhidQh8RspwCKyIE+StX/J06uW14H9
YuxFJTqcovzquz43BjYx/eCDnnWnxDyzPhMCLAI7F7l90Pib+raw4agpoNFtcISe
53wnXKjGtZmmuy/3Bp29BA/ufAJ6cfwhDUr82bygUf72FlOcP178MIqmeFaRrsPR
VWLE3QF9NzmvQ3KoL4/ELW/Uz6NHmBaHhTW1KyEOPcg5c5nd9zhbNvFio0+LEuVq
8ueYNHpqT6Lizs2n5ZzYliUP/z4pxVDnq07+auzAn3AJNiKiKnaWifZwJ+RCYzFa
qM+V6xongpR2hOHfpOmM8AlHDdP8AK5yarm83oggi+VAEJc7IlIoFLVxYsxipv34
gu7XTKyp4v9rkU0F5CygLOPDaGqAo8/5ec/ThLd2Z/qvxfqri+DvcyUSGrmVWh9g
G++zMTKc9SN4nBmWFhDerpV0dgRlURp6gOTwJciCc9qC26mvlLKzWYJb/xnXocmA
GW9RlXZlh3qsNYsaGcdJtFn7gCnweeiT5XWji0nY/4846+74kk9WGUdNTxwiubRW
mcjrC4+CaZZMfBylogV/Ejipfpdny1EV532zE2e8S6WlHJSpZEyEM9Q/YHnjQ0cH
bxMbA7q40JAIqyEpRFlKfyKXEafCjCD1Qr8Bu2fl7VA5ig9RbIu2/8J6hybxo/lV
DsqFVbp+ZE+9578fcaTbOSp698zIhFu3h0/oOIwoFmYnAOnfPxc8m2YuGspjLG7b
j4TPAapyDYWaqr7UkYoQRZlfOVshLiE5G5CtyWTJwFJFHc3uGU4ojmQ+hy2CewFS
A0BgoNjWKeomgNXze+YJZB1/bOvSW/kiMzrpKA5BTS6rei7TpdCEwt8wiAuaN4Vq
Z864DL8wY/nBFVbN7ogvYF1vR7vFx2wrYcOW/VKB3+Td/IHUpFfBTn2bO7n8DJvo
83hU9sA0NOGyO/AWZU6e/vOLOTI00waTNI2aURdWhk/mQ/CGzmRnraxtbbofHNmb
6/LoZfH3xUVY9armq8SXzeOhzpjriqB2q0ZJHTP73yHzWUnNJ/Df4ZH4dzrDxYI0
cxDLYW9xFnFRckh8gsKWz4YcEOTVePY4FGwzO4ICnv6wQ3k151boJ/3F9Q1pPL/h
tpf/dGX4LcROf121tvX4ZwnkKAJoEl7lENADhLS56On+WrEjtIocIHGV2En1wsl7
H35CA4jMn3Le98n2BEqzjsfFH8OTgGLCSSPfhq2+oDYZzo5E1XiqCMzJzAbT293l
nq4QfOd6TF6Ow8liSTMSgwWmJbR9QI2+JN+YK1bfpeAs4dsVvC7E7YsmIQNS2aXx
Bz+mirjXkIuGioUddvXAzyJ/2v41bB2FN1U+SbV6kms2WFOMOCeuBO0X/xOHFNZS
M/PiX4wKNqxAF6Tgw7Z8gyR5JdXZbAWO3b01HP2FhSBZkodOP0bepR3jEhkruf8E
QjYP5VoMfAG56KUiySR0Z38mNW0wPxGcl1Zb699fo7gLtYa3HyGoC/kWXdywKMOa
s3+//RHa2KmiPkh+VVPbpGj64xzkMqYwMULhyIB2amfmni4QbuaVBwTpHeg05wQb
VpgmSVauPi5NY4m1vSsAbnRCl0zQlNjjaJ2LHYyqmLxuVnYMxX4YQx1rwlJIiYrP
5tAEhHcpURyNEuxh4pdJrP3R/2u56cQtJ2gztSYaS+ui2U9fEi5YE8uxqq+qbCDZ
2+Tbb3sP6GNwNHjtNHHftzAvQ5soEPtjzNWORxsyGNBWOr7N7IGx+4i2BexMKX1X
BF7pQS884iQV7PkW8ddBXW5FpyOjzosAvhxXaVe3CJCP92f3TQlvLYvd1EF8pLNP
MR+Mab47768pTrgqoRjTpsv6trGcK7VAAv5v1c+oR1OdQHtr/shDW1n3PE9MiMAn
izdiO8f3gSP/rnMAPbI52pDp2G2wvxxAUOdxVo3SXeeWD6QyJLk5xiPD9UJh/8qU
HYS/+AOPDvUhu0hCMXy6b2FqA660/EbncIrUxbzN9Sk2ETaWrLAjrCFG1g1nnM/P
gjTaq60iittT842nroWrFP0irY1hhT3mW7eYlBqP0mtwLVXmF+xbkh6j5EIcZNlu
juqKIVooG/IS8O3GIWg/n8Yh8hb6YtqRYxxswUN/Zqq/tKey0sqNtZ83uVoLbcO/
6di96O56gPGRvvkp4w9fUaV42QnmwA9FLLL6QlCICUISmJoGpMWWtrXrTuqPlxkQ
qtpQSQ1SRKZ24tKgerD6HW1OHoHqOqfZBNzJmPQBod1AfpbXG8vIcORbFbUUSUNf
qizST2QdDfyfZ7b+Lsm6Ci1o5Oc06em+LONzbvpW2U9SI6ByRVDf9jF561F55Lek
OD+E4lFjEEGrlZoGF0uNG5l1e9Zh0sTjJ4zODkm63FgivKCvF4LaU0SYieHvTvl+
5eDCgd6q3Q8pKftQKXvYHpl6EiezeD8/oJruYJwTdvK38rIf4ltZazLX98icjmXC
pwghg6OmwJUQUSFrLGsYWMHAX00HV1pR+pgvAysiG67/T/Hn9Ywhqh9ef14WDQgU
c3YNxVY0NodqknvqP4F9ufUZZJdizE7kD8DWUejpTHkcaNR1TKnigZAdE8/kq8IY
xad3S3kG0b00c0sx0U/ZVQFQK5oqrKrreoz+Sil6DRGLaeYbRY8w7CaV3R/34+o1
wgz50XnT+wIQR9hRHvQ4LhNdzxnd+FotsgG4E4QUl6mtwthfIZyi5k1UVYv1LG1J
KAY8OfUUooHzBaDcVuR/Q5sBISglubuqZVzt5EyC55FkMHjH3byeVCKlWTiuj6T8
e1nZ+aZJWKb+gEpUANvvLT8CGDLIsInK++RRdE+pGJZmE9Wzvz3dC1U+D4w2bo9m
4x2ZNN7qc+NV8nvvAHgwirllfOqw3A/lW3ZZ7OSh9lJ14UHSOGpFgnESxi0OAXKS
p1FOLrF7KUtX/IOZZEwc68Ih9TN8Pu+3nVIa3jhxtzJkQkObOqHH4BJaGNg1iZ8/
B76Na9LA9XnLgi6LVCPLg9gcwDXFvakKzSRKsG5dbV4Fl1SW7CxCAoVr2Nr0Oh/f
EVwe2x5mcDfbuIf1HqTq8Hd5v3rJzXmLOsKAuy4S5pohzFfliXgSL+dxMHF+ea4k
DUxQqdlfTYhupUFkwrMKTdMx9vFOLi+xQbU/FHtIxjij8RmU80eVGHpnWxhpDxb+
zafSDvPeYtt2sbHQNgEYLFYWsqXs+/Gr4hiRXPfanTbV+6RKifSsk/3qeQMqdisj
jTWcl5J+zBnemP+t3yTEKcbSnv++WueprlvBBFqHFqBzTkeZ8/4lbsi1lOG2dzuU
tpd8K/Vu2qafAh2+4MBJ/PWzlmiokxGEDaaKyg6Gry6R4nOpx4lTkr2ZGyk/OYff
RO43XEjaotVJVKghfHGlHP+L1wGyDj8oRZ2Y6VCc55sHJn2A/LTDbBDjFEngtTKP
ON1ImDXXngcNiSQy7T1DX8oSkComQmdD/1Mqc8qxrF0P0VoQcXYLiVfUcTyUBY30
+I+5mOyA+PmZ1ot+MhDsARUUV9662erHHI7owVLiT8qMosA3y9oFdQe9hVAI9Wxf
hWSWmx6sF6RN1j4/XL9R0s9RNl7GPiY53HluwB0PsLpVjtIYpyhq7ucPt/BR35yJ
MGnNF0bxz1dZJfWf8eyepEb8sWSRLjVvB+Qy5idA6Ug4N9YxH1YXUTh4wEgIOod5
lLmUyi3FiHj1ej7F5iiDwLlnpqarsvXlZEpKG7DKn8j2iRIfCF35cp1Qv7TcUitF
SghgLmS4eNrIuehgjBGuS3StCa2rigrvMgW4wGbtpIPst3qhN0eBoXrv1FVPdyvE
feHXvpms+nvCmgRqpInDv7AEg0B9WQ+A2yU2VH4DDY6QZ6HFv8B0P+Hk/9M2SQYw
11EsmcxNL6gvFJaH8hfz7LRw+TD5m3i0NHZpc31hEtXHmEtKzqX6jwO73cuUqdeL
od8v82X2h/IaczTRYi1jcapNcWimY0nfmZyOiVHOYJL7yE/rV1t615LN/Lh8gVv0
WRbpKslZjMe1eOpx2ReA7mr2+LgHNaHqq6Op5rWZomL6gz+3kznGUQygKkDEaTL8
m8duKWvOhxthdbW1sSmGzxsqBru2WXP0OQLaiKa/xWC10zM6X2vTxZhEXbum/YE0
LVj17Ftdnhkb+bPQV4FOHaqMbM7V4V4pXmtf+z/6BnNjp1eONor9euc5/1Uj8Tcy
4szTOD65tkB875A42jHtYXc+t+AI51RG+5+GII+SAP6EG7z4RMF4arqM3VhosmAv
mrkt2+iUIaR0oq4ExMARkXj49nuTCksoreWRvjeOrbLd4elPKcdApvf/CdaGh9Ml
iMvtfGqZl3hJhYruYckmnUN0rU72tOOBDDwlJYdP2D7eEUwE4yovLDp2nZMb2YHh
PcyzncXOZPOv0cAH9LmS4+JXAuG9lwO4DvGA1LdQyJoeTK3RKEf6y7Or3PA1mZDM
j53Hpdh1zNaUhWkYGxpBow==
`protect END_PROTECTED
