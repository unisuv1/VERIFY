`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
OP3BSL2SSGdFc+/mjjA+uNX4s3/ensVgMX9JCLbQ+/KmtHjEpohGvXC+JhHmX7Xz
Kq37bwTugTyj/xxg8TqOpGS/1epuR7KmQsJ7F0vPgD2QQhI8kg7GVCwTLZTfX2Yb
7EWVC1j0tEsqPVyfKqUpwfxB7sCBs088UzF8gb9ffMBKhcT01xMz/6ZKs3sf4w0p
P+/eKtjxYpQjs5ipPALKgT/aZxM4AbSD5OEllv+vnBlG2rOYPTrFaxizUBOVcRdZ
cSF66zz0BAe7Czd+N0k81fsTjDdBtArPMjRe5bN9cDO0onQ048l1lkKOy96w/x3A
iGRs+xOOF96p+WF6E2SjWq0yt8mzZ7qt6IDlDU5YsxYn/ysIJ/GT6hbBqacpgS9x
oL+GBSNOuJfkQ1m8yuQiIVKnj48nyapZv+DSooFwNarqBpCCkDIu8RnBco2io9v5
OYUB/JPbpg7bpJCPMADAoUJg6FuKxFNff3AmEulOro0nUEuSDg5TNdzclSd3WuTE
L02DWJb7e0HrMTLbJyRsthGzq48ldu4gMyvQOnfRYkBQcw3k2jJXz+H37bKAStmp
0Z3ImKigCIW/6/qT+4A4Re/Lecftrp6/v2Iqm0CQjPCNZdPXWCHHagAyGM8P/oWO
8ZFq+R+Q4NrZRa+KyUhCkGPPFp65619oq36fy2aKnzP3dLbvZCK9uACPMAPTkDiV
j877KtWESkRF3VowExZIeWUl5HFz+TxMNx1j7VBqMD4vcUq0OtPZ4uIIIX8lZ/lD
gAa5dVFJQ2QOr8gYaQpQ3MrFmyuEj7iKm5tfU1QJix+/i73ss0ouOr5Cjn0BN/T0
6+XTJ0a6+ijtjtm7KsP4wcom2V9AYcM/D0/bInA6nRPmN49mM8u6t2Yb+BBOlJNe
Qy3q3JiKuROi7hj713/M/y71dA+oiH9GH/PP8ZvMG8m3a1AdouXvsKu9nRwfke79
fHs1v24fkzepj5dv2CszdX7Kfooy30Yl00BaUoOrdJeLVXgnJfDfuxJ/odiXqSNF
/BoUanbb6fDadDie4/tF3x3Cd1JQ1A1ZoTpGQfvJZXIkIKa95iQPCKvR0tNxIH6q
UuYDlsuZHjpfEWQ0Ikrfyvas/Q9w2pxCRG2kh0Ok/2rahDHO+hpB+LdFPBcdjoPo
yGfmeaKcACUjBCdShaKDTMX8ozJOfCY+RoLKeY+0Lp9avO544s+unL1akLM/JNsv
WaJ6fpAmYx5NdU5lJmwrYvo5zhMNZnMfe84Syq+mo7K3QOmedq2T5p6r4I+Jokln
QisBZVgA+zT9RbIWODpiRhcvY3IkI31ioBbwRpBB0mPJMpEFngNL04SLp8pfn73+
u+UoxsCUtEPnb3fNjbKFcz4JUIqdKvMLhGZi4BrCXT8vCo2UZ8pQ+mb/blcqXDx0
TvIylmpbD1+vuo2f7v4eyJGfnB1PvjcGN3pRB4FjQpqUtfv/PFdO7yWiFAk2hJYb
s2RSNzu1QniZ63gaSTflppM4hR7yx9229sQ4w0aJ0B0Dk1lN0I6enoopBmZhPOiZ
6jJBGkSf/GKP9KMLqwpHPQ0XG5wCIUq3SHk8RgPy33tPrPtwJ0m5ybSJLVBsqg0R
v+iGykVupRGw8xHJgEL+Xh8bRKozdUbqzpEO3YMJ7ujXj+rwJK9Q+VGqNo8luI6q
PJtK1OoFVGJEIOj2RapW4RwhrCuQbzfE8XW/7Ipoas/ctidRDIIOEYR3UlW6OKT0
+GggWyUZtYJT5GOhw0SyF5PaTQy4dkqcZdIoEbaoVwZtykGjvlPLWy1+ZC/IEC3z
ZJYFqv7kchaQOjr/CnLC06V7hsRHumcPqzi4+PaGerVJd/WGqekIax0qQzJjvutl
I62nXXCLaXGvyCwaZbic9CB/pMhmv6yVHscBie5BMOfy6OLczz1SafIH5QmhCGDE
snnoaKaOBnmRLuviuP3Ns1V9FumQmP0Wjy/CgGQ4Fw5b2lH6fXsreNfHQettyD7S
L8C40X3O4+c7O8r+SGbL9ZJiwfWEAEhZCDVgjWb0t+/3Vqhawcdnv29iVgMyUzJe
xUOxE12vaZnuMLCnHzJD+dNythvE69QVrwLkIrUT7FhrvU42BQMLbD/6Z2bP2H+5
5zlCtPe6sgCEBuvgwPim9/cGP56pUUnxcaX/mkdLe7mQcAWW+z3TLdd/r3bJFI1J
tDo/DB6HtYNVj07x/7DJ80cCoC/zpfQP0ZHd36/gZQgVPctwvbpu7t/mAI1jN0kJ
Xx89IUjJ2I4H51x9vpJJzh0cQs23kYVvieWltf9F1mLzeiVhTIBYZjdqUxyqteD/
U6JbSIaMBWd39JzyFQu1klwCfZz/Keeij0d5YKKTsI1E1KczvMBJhsxcxVT9v5gn
PPCZ+Bz3Ijk3r0r0NZFPuTIbu+S24JnphKNo/wuWajQIP/z0xRGRFw0a4WJZtZY5
b+qPp1bQYhfc5HVmfiLYa1w+YlaVnqW67b+7j1uEiJ1nwbFqvyXiwJHoKwqRpP34
3F3uJdUzB6lQRwESzzRKINPjVnRjsJHxOc8wkiO7x2r9mAK6C3gMATUpSQGV/hmZ
M1Fl2yYOEoRPPOa6O/+EIeb/hIQkfxYmFGDJmRQXNeGjT1k1cLukneL1O4/5R7rZ
8pJ/qXFVmD3Z7/DrBzriP+zTZXG23iSvUn2xYbPrHuMwgfw87FZeAp1PGjIKO5cS
GNw1N3u6DU2lIfi146EP4XqwNiXeOdju49VNUTK3H1C7xPmfgZj6bPQppXvzcPgz
YGGtnvGCvfPh4MqYk4wJZ32g8Tn537Cqt7Hs/zTomb90bEpa747ttqeV7xetlpmr
W6Q5tousFU8XhAAPqdIaMbLtsZi4rO2HEdGZN37uNB+kaaQBsh8R844c87A16E7s
O81Gz5AA/DyU4HKuTNLfas1e3q7KK1R4pX0CD+vKcX5N7q35kwko+HIDlgil4osF
EwuOcHZbP9bjKWajyCqoK1DQ/pVpbbG+rVMQm+f55iwfbmi9bM023QKJLj43rHz4
JL80UFgZfmodSdZ5gCVZHfG7VWx2RDxJki+ISUijtlmAwLtHNUbIFJBWwkZC2DEx
Rcxh1EKGeiNyIj947z5DfEGB8QZy+KJCeZMUMVNxHS43GsVC2nQfoXNv7leTp0A5
hkSKLqCe3if6uLE5MNhs4KMRd5PcRJwJbolcLBSlzyh4QRUg5MrYZgSF9aBgyGvp
025E2WUrbCvroZn/yUu4jQVT21Jcgi3Q3bcZVZeAYJpAr8Rr1vGi/EV7mt/j2ISY
7VPqd9B0tl4ys8U6fEJmocZjgmeZNepkKyfruljEQ6FI1XdSHPXtTz6pGk+UNc9m
8pt7LGm4JKU2yFOHnxR4mep6PbXUKNYozlbpKE27iXZ6Z1sQ+4oD+tbChHjEbW+d
S9JqUQPtANCVnray0j3KRelFbbAjdgSrLfL0amSw6lkl1MFegbU5ML/YUgCogOoB
FCxlkkzVdmehKq9b0APJISOKle/wbU+SrGGmcDYg7YfYZXOLA25MVZVTziTocu48
vi7RfyVNHj3hgsSbJaOKoA8rHISniO91mh38X5ssl+k58+cLbr+PG3jt9IWrj/xi
bUnkFJVl77yOhS7RnslDiRrHslk8glsgO7NczfJl03i9BtFoZANuWMgkPumYjAr4
7I+yAa7K4nVwNIJPVZqHMw==
`protect END_PROTECTED
