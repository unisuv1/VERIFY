LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

entity XCoorSystem is
	port 
	(
		Encoder_A	: in std_logic;
		Encoder_B	: in std_logic;
		
		filter_delay_time_encoder	: in std_logic_vector(15 downto 0);
		filter_delay_encoder_en		: in std_logic;
		multiplication					: in std_logic_vector(7 downto 0);			--- -*-
		gen_en_encoder					: in std_logic;
		
		nRESET      : in std_logic;
		clk_sys		: in std_logic;
		
		X_Raw_A_Filted_port	: out std_logic;
		X_Raw_B_Filted_port	: out std_logic;
		pass_dir			: out    std_logic;										---�˶�����

		X_Coor_Raw	: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)		---����
	);
end entity;

architecture rtl of XCoorSystem is

signal X_Raw_A_Filted		: STD_LOGIC;
signal X_Raw_B_Filted 		: STD_LOGIC;
signal X_Raw_A_Full			: STD_LOGIC;
signal X_Raw_B_Full 			: STD_LOGIC;
signal X_Raw_Filter_Lock 	: STD_LOGIC;
signal X_Feedback_A_Smooth_720: STD_LOGIC;
signal X_Feedback_B_Smooth_720: STD_LOGIC;
signal X_Feedback_A_Filted: STD_LOGIC;
signal X_Feedback_B_Filted: STD_LOGIC;

component EncoderNoiseFilter is
	port 
	(
		Encoder_A					: in std_logic;
		Encoder_B					: in std_logic;
		
		filter_delay_time			: in std_logic_vector(15 downto 0);
		filter_delay_encoder_en		: in std_logic;
		
		nRESET          			: in std_logic;
		clk_sys						: in std_logic;

		Encoder_A_Filted 			: out STD_LOGIC;
		Encoder_B_Filted 			: out STD_LOGIC;

		Locked						: out std_logic
	);
end component;
--
--	component QEIFilter is
--	port(
--		Clk 		: in  std_logic; 	--100MHz
--		QEA		: in  std_logic; 	
--		QEB		: in  std_logic; 	
--		QEA_Filted	: out  std_logic;
--		QEB_Filted	: out  std_logic
--		);
--	end component QEIFilter;

component QEI_X is
	port 
	(
		Encoder_A		: in std_logic;
		Encoder_B		: in std_logic;

		nReset			: in std_logic;
		enable			: in std_logic;
		pass_dir			: out    std_logic;
		clk_sys			: in std_logic;

		Coor_out			: OUT STD_LOGIC_VECTOR (63 DOWNTO 0)
	);
end component;


component Encoder_full
	port 
	(
		Encoder_A					: in     std_logic;						  ---
		Encoder_B					: in     std_logic;						  ---

		nRESET                  : in     std_logic;						  --- nreset by power on
		enable			: in     std_logic;						  ---
		clk_sys					: in std_logic;   --- for A+, it is 133Mhz
		
		fire_multiplication					: in STD_LOGIC_VECTOR (15 DOWNTO 0);
--		measure_sample_num : in STD_LOGIC_VECTOR (15 DOWNTO 0);
--		multiplication_num	: out STD_LOGIC_VECTOR (31 DOWNTO 0);			

		synchronization_en 	: out STD_LOGIC;
		Encoder_A_Smooth_720 : out STD_LOGIC;
		Encoder_B_Smooth_720 : out STD_LOGIC
--- 		Encoder_A_Smooth_1440 : out STD_LOGIC;
---			Encoder_B_Smooth_1440 : out STD_LOGIC;

---			Locked_1440			: out     std_logic;
---			Smoothed_1440		: out     std_logic
	);	
end component;

signal X_Coor_Raw_internal	: STD_LOGIC_VECTOR (63 DOWNTO 0); 
signal X_Coor_Raw_full		: STD_LOGIC_VECTOR (63 DOWNTO 0); 
signal pass_Raw_internal 	: STD_LOGIC;
signal pass_Raw_full 	: STD_LOGIC;
	
begin

	
	EncoderNoiseFilter_X_Raw : EncoderNoiseFilter
		port map 
		(
			Encoder_A	=> Encoder_A,
			Encoder_B 	=> Encoder_B,
	
			filter_delay_time	=> filter_delay_time_encoder,
			filter_delay_encoder_en => filter_delay_encoder_en,
			
			nRESET  	=> nRESET,
			clk_sys		=> clk_sys,
	
			Encoder_A_Filted => X_Raw_A_Filted,
			Encoder_B_Filted => X_Raw_B_Filted,
	
			Locked 		=> X_Raw_Filter_Lock
		);
--		
--	X_Feedback_Filter : QEIFilter 
--	port map(
--		Clk 		=> clk_sys, 			--100MHz
--		QEA		=> Encoder_A, 	
--		QEB		=> Encoder_B,	
--		QEA_Filted	=> X_Feedback_A_Filted,
--		QEB_Filted	=> X_Feedback_B_Filted
--	);
		
	Encoder_full_inst : Encoder_full
	port map 
	(
		Encoder_A	=>	X_Raw_A_Filted,						  ---
		Encoder_B	=>	X_Raw_B_Filted,						  ---

		nRESET      =>  nRESET,	--- nreset by power on
		enable		=>	X_Raw_Filter_Lock,						  ---
		clk_sys		=>	clk_sys,   --- for A+, it is 133Mhz
		
		fire_multiplication => X"00"&multiplication,
		
		--synchronization_en => synchronization_en,		


		Encoder_A_Smooth_720 => X_Raw_A_Full,
		Encoder_B_Smooth_720 => X_Raw_B_Full
--- 		Encoder_A_Smooth_1440 : out STD_LOGIC;
---			Encoder_B_Smooth_1440 : out STD_LOGIC;

---			Locked_1440			: out     std_logic;
---			Smoothed_1440		: out     std_logic
	);		

	QEI_X_Inst : QEI_X
		port map 
		(
			Encoder_A	=> X_Raw_A_Filted,
			Encoder_B 	=> X_Raw_B_Filted,
	
			nRESET  	=> nRESET,
			enable		=> X_Raw_Filter_Lock,
			pass_dir		=> pass_Raw_internal,
			clk_sys		=> clk_sys,
			Coor_out 	=> X_Coor_Raw_internal
		);
		
	QEI_X_full : QEI_X
		port map 
		(
			Encoder_A	=> X_Raw_A_full,
			Encoder_B 	=> X_Raw_B_full,
	
			nRESET  	=> nRESET,
			enable		=> X_Raw_Filter_Lock,
			pass_dir		=> pass_Raw_full,
			clk_sys		=> clk_sys,
			Coor_out 	=> X_Coor_Raw_full
		);
	process(gen_en_encoder,multiplication,X_Coor_Raw_internal,X_Coor_Raw_full,X_Raw_A_Filted,X_Raw_B_Filted,X_Raw_A_full,X_Raw_B_full,pass_Raw_internal,pass_Raw_full)
	begin
		if(gen_en_encoder = '1' or multiplication = X"00" or multiplication = X"01") then
			X_Coor_Raw	<= X_Coor_Raw_internal;	
			X_Raw_A_Filted_port	<= X_Raw_A_Filted;
			X_Raw_B_Filted_port	<= X_Raw_B_Filted;
			pass_dir	<= pass_Raw_internal;	
		else
			X_Coor_Raw	<= X_Coor_Raw_full;	
			X_Raw_A_Filted_port	<= X_Raw_A_full;
			X_Raw_B_Filted_port	<= X_Raw_B_full;
			pass_dir	<= pass_Raw_full;	
		end if;
	end process;
end rtl;