`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mkizW+Npzxep1aK76PwZPncnyKhEU4v7BBThD+zByXmoVwI0h5FNED6wL4P9YTNj
vBL7FF++IqRI6eREgHPMwix9kig30L4fH2iBPjEZ+5LyJDeqW0s4+mjT9W79oGcB
gFY6uxwPR7ZCnCSQj7U2r5BZgywEWgEFzYa+/D6FDLis3AmmSKcQZbTfNip05hHj
wIapdJBQRowjwmDco6NT0wYTXe3LqfgeKsGNa0RuUDbCqB5X3zCT2MrMwP3Q8d6C
BTIMpMu4cJX9qoVSoLd1cQu4BlR2pzz8440aRwuM4HVQX9FJUBKLDJ1g9t0uOmiF
53or/KwUrsjoj5utwh+ZDst9mh/KxzetwRP4t4TO7qc85QniBt93DGYsqbaSRSN+
iV/2dUPGQD+23epZhqnKMvTKIA9JwE7WcBcxmLQ1L1b2imJd3AiZvkxLIukiZrTL
MKnJF6GMqQs8eG5IhHUQ3P4oTyzIRBnWEwLtCTkR4CPjdzj6VGIaDxFcRNSvwy8j
ZrnD0scVyDy6G5VxTGG9wwV9IGaTKmMbOGQVEMbHBCmt6ZtPrfgMBBFJsLzY3YOO
5efvA7sIDXeE/VavLk/ESIS6mcDbDZla1OQg/3hbFx/pfRr8Q6SUpUaB/gZ8O+cz
NwycdAvPILf2UfVms1RtiQQ/sM7lEXp6ahkinFlkC47VZJG8GOMsfxLmPFEKxhyU
/Zvb2wgLX9cAFPBKLzFVwt6l6gZm+dZTllbuGyGOmh13fujb+Ut1AqrfnH7tUmM/
OhhIA4elp0jFmgpux14A8rHkcTosrDefFMyysMcG2p/GpEDMZ4ck0c9Xt9Q3wYgb
hbn9pVFWUrXMiIbmi4PoyCCwOgtpSML9F2GNQTF+AHGm23VBresN2+7bOTfZBxPR
99ocDwLaj3u/GcNHahIktheAMGVdSHTJ/yJBHmDdRaWZBad8cl2TWpWnakk+Ned1
4MbNDhMJaryhZciNOkNSH079zEu7CSVLy+nwN2KTes8PtgrTORjUCjWkTkTMYCfA
bFSf4JDmSoCUAdQxHmYKJvkJ+ON7rWvIzosQlHlfhuKzy7KS/hWxe2DwjqCejc1I
iGyChlZjRcytpbt9kZda91z9Fhj+AsNm5oHl2tCsHtOSZiXU3+2oVy3/INXPaq6K
Fl/qSO3PAcrsLFpmxVdQVwJGhJsPunPVcQihjTA39+N9gEsuNV337G+En4qJUxBm
gyWS9bKEp1UnjEZkSQ4X2K3zwoJbzR81yXjeIxvKhzoCXlXoMgbmqHAhbImcoqYc
j2dTN+WUJxlFn/0q8d3ZhsnQfDO0vNSay/LeXFUnBxNvMt5t7u9SxDFyphyRZ2uF
nR1c++wf8Y8hOkXasw1AbGXouk61f5b2sW+WKL/RFtucOmWAUJrHtVow+IGvfN8V
13Li/ENMJrIbN1WKz3CuZAwKkbKOCzI9yOQJd6/L2PlgtFnVniOPkem6U5XphUHs
UXCA6C4J8RYqkL0+I0jZQvc5mPxEXePJto5FfoORfPyqhw8j87asyHZyIeeH60D0
mF+E1l/9RLRU2cCRylFphvQvqlifjNrH7+YmF1qqR05JVQJF6FZM2UgzFq2qQovl
Nm44Zz1aslEryHwCvUQZWrNKcj+VpVnX1Q6lyBH6Q1Q7MNvHlRynSmI+C0bDraX1
cV153Eb934DLwQPUpytXd3pjXvFQoMXX2Zx+aZ0Id8pcM/AXymuuncSsKlNVlXCT
H362CEOhfLbRBLcryfP7IN7istU8aTNmd8pSB7BDVQJ8erTGcjiAWBcyeMQezErc
Mac1ubstTKPw4s1Ezo0nWm8eOgKwmYlZg24WmssHfLInIdIXJ4L0ZaS8IMspYOBo
BXkwK1Du7PTeRwTJXub/Gca0BQ036ENmu1sLPsjozevEmVo6Jk8ydzyJ5vcqvKop
XkOkxy7peeGyspyypb6ACPDqa7AOXLfKqX0ko0X9AddtQNPzbnVc08HkPQBkMYOB
RCo8gR+PWM3EBjFEow35wp6xZsvu1SLrjLCAZN7yNC+jqV9JR8nK/X8IFBTP/9qG
af41NY9g1URh0OqGbs6KnKQSoeAgOOJ1BJnqN3ON+bqwldjYB8tORnPhm58zuCMB
u4GS2/3VKkRI4OSxvZENo7aX+RsWWivp7FbMw9MED6U8XSu4oQmPF4ocQ9c3WhKK
HY6Ax4/wN+LGWAV8vqz6PQQjo2IEP8cGb6SAjm2jyr/WpDxtTjuigVCRQ2egY3oq
Zoz7OL/mNEeWc1vBDlIL341c2lA7xtl4ZJ1Q2LNwzdLGXxF2iEgh0XqTmXSCwodE
b/jzt0ML4kXtzHvskJieSMG7aEeI5rVa7S368MDDVo9mlxEoBjirCamu0aokalxl
4crmRO3orQGdiQpNYhkCu9kmTcHZnaJidX3e0EHXVvTDKI0H92FUNT25Alnu4IFS
nHge5bTbIxp8nJccf+eO0WZhhXusiF9mE76gE4/sThcpq8HUSVT0ly1iagpStoDF
MiJptuUWypXAzu28E4ET/7mcskoTy0zK97YdSFae/9JmeLP5pRIx2b2tYRns7EV8
82QEYhhCa/cq94FUxtMbElqAZml9G5iH9J0HL+EbYTadabHs//l3f1UxK40XQKIa
TK0yTH3rJqW/STHjMqUJU2znCuWoHzHtaE9sVRkRgaCQbVIwrNPRnSM9eUGb84Os
SaOwcg6Qb/zPQjtJo3+UUGCj1x1pfv2nbH0J5kpMazf2+PgKO5czW/meEGY95Puv
EZ5tfuEe9BwmFeFftf/51y7YqNEQGR3fk2QzwT7YX3Fn8bouXkfHIgQQh3dUbW2b
vEW8wKVq1MbVDyp3Y5ABE8TH5jy4XAzgj/orUb9750bPewqXyYDPgEu2/aIPShuo
lnyOMI5qciFokqfLErmYGSpah7oCsgegHzwaYpNOX29KT7CP22h++TC/ktIFSw9d
xHbWSSnKXtvDpKoDJAwNrwXZl6IoCdqqtcNrY4XoIByJdWm9Ca94FUNNiX78qdln
rlkMMOxySkzr+kyluHWgdcTdgMMwW75fwSaCf5mdHOaLSRhey5OR41xpK8axoO38
bHxNvgjryhcNi6FGtLF2UZGL+DkWrxsiWokhVvvhgfGie5ZI0ZHT6Py8rVySOTpX
/QUrSJIpcF4R+gttbO2s/fq+y6vdu8KkIJ/r20Wj7MvppNivmvU03EfD8Qfyn71H
Bx8v6QlZdqtg6NOqUwNU1kq9al37Oceoe6H4XJtPvYkDrKOVgtLIyDcWdc3Svshv
wtDUt+CoBbL5UQY4RqZf8MQf1uXqe19JJREU2jFmyCAQw6SAYPxguXpl5oZBaEJ8
RMi2qoEEk+d2nXalgXETwsGwCngles/js1l2fRAMtnijtJywO3sQ3S8KoYRGDAGk
ZCgyFIRkdtWbsFJdL8PtxnTkKLyztIC15k3aDnab7zKYPg0E/eRMlWN1eDJ9BWBe
BP4jlHqA/s38LMhMmJlCV24crmVn+fNtf7/lbjtHBzlnNHMcO4KYQA+WzVTjZtV5
Ani6+S6QS9OQyuCyXMXDe0C/poUjS+nyr8yAxQm+nzL2hnTTwyFy1D2tGGuhgnB3
ejTKhErg+JvMRL9Ci9NYZ5LL5lg8fBa1z11rxfvScKtpPSTZvcXaGfuEIeQkVt09
Amb84FV3527RMbf5LFqhsh5D8bQT7K1+8u5creY8yQ5vOnQ0aSN+9qG7Yf+xw2v3
TGE00Qs8lPpQmPhVZpBxZ/+/rM7bYWEXVXgvSbAgsGcnq6ro4Ymq8wSSWoMrZYn2
YkWDLnjTzhe6FYm/vc6col0WIhYmJ/mYPohcL2d/Rw2LnIDGEagQIZNeGQEqMJRx
sG9xfZy5TO0UpGgXaH1hj+wHxGaAtLroXbZnVnf/+Xi9XeRNw1ue1dtoZWRW9G23
pOGeiAo98eU7Vjw6kLtgJ7TkFDcXtBE3jJNUG1iu0tC3mTaTForQfcqyWv4NzlVu
MxvKmNQ8LOouvbwNhtFVJ0D7meKw14psxqmEBOpuzkTxZEiSimr0zXhKr1ERWfDa
b9eHjR/djvV6NRozU99Agloduzl+3XhONhdymg5LH/9sQ/pY7zXjTij5VbMlvDjO
7LvXOsZLRbnfYRLaeSsPECjx324/9Hj621b0bGjG9TWMeQdXe1T0fzDVXofIcFoJ
R+p7CpFI4A9NxR3BI6aXA8aHldh+/wSDU2dEqWfTmEm82gWAJ7Zh98n54hIWIrlU
fEd0n14Zr9oOE8wDB1OM0w4A11APdIiCNNeke4M9egBXdREbYEhlLCDNU6JwpzEz
0zy7LSHwuI/3445O/38yelRF/DeUxXfXOqNSw1q95B36yCS9wH/QGkGqSAJ03irE
S/VAv8gS//30RDh4S1EU3LEGoVgtzxj6uxPF+nx0jz67DDf1QxN1Fs8AzZvIzUlU
rCKdKprsr7g3ny54xTkI5czop+WkGiC/O4tIqZ/ad9QtCIByqNLLO8Gcaa8EJaM4
tkEb7Mf332T9vheXb6mwiFUK9yQsCfEVQeuKoFSpLXnDluhhs+note7ISL1o27Mi
iAtayrZ6W2ZeEDuf0rGbFer6BfyoR9s2JQJmQLf1nBHygQYbuqW5qQk6YhAi2IYe
1IT01DZWY2JJrt6yEZjYz21/DIOdUSDWunNxx7QJe/S8/EZum/oevBgxoMCNI9nn
/9PJxIoOMRXaMssob1esKv+psZJp+wlgBSIGdUa5e9rx4wCZ7ZsG0uvXQ1tlztdD
sLO4/CAtGZorzBl0gblR4Ty8f5NP8Dun6o3iJF/QL9qiKcpBc72dWLN3BAJsCjwI
f0NSUKGUKT95pQTwqrXMjgcj6arBSqPeO3vQuxmMt+360vpDYyaneUB7N9AC1jJ9
jV4iKHoxIcMZ2S/WNFmjgAX2nvMTFMnXDjmILyfP2Ey74B31ILq06ydtCX6ustpu
dclnJEc+pYOGq+kQFYtYq/yE4+tpp2XZYSNIY1O0OWOuGLrq7sMqt78Kdwh+MTYJ
Hz+CMESQ5uiqRmgyiSQaH0ot1/XIrVaFlQMYTVuG8+T2t5bWCQAWpTPOt7lpx23f
XPACtuWicd8v7j70nvKxGTR4pjkUbSl8prmoW273SoTnW96KrMM2nXnu17YkhWmk
BTj8opOgfXuEeXVw2woAQLjXMc8Q7oU0ncvd4K3VplVRKnZ04IDJG5camxV4h4sZ
+/yVfDMiexUjjnFs6fW6WSaw80+WqXYxnstX39SwVtxk3Bs5LEBuQoV2PPLx/5im
s5A11MKoX+XjndlqlSOiBWJDbOpHgzKwMW/XkhKsdhH4HJJmDmh/o/cEKj5gSvIA
ib91ZCwEA8o4szn6u7whUzPXDL4/gGj5+cIFU6LZueqqYk7sTCmJCI1SQuKMWPPQ
RAruzxpNwy92ncSAxYJNvdPd3GbcrFTH90l/VinkwkHSCcMmbCH2qpDPKrh9sQm7
n6QxNpdtvos48oY2IrbL4D7OIcPZ2cy3pNKqmrU6sVRyVerX/bijDhjIM+JEhOLP
UxEE5B1jVg0aR1YI4/BLGCp48PNKUKALRJz2Aly3c2eJmgfHsdgYHg8c+nl6hCzm
33bqKS1Ph5gtrv/+O6BITKGf08aVziYZ3FLtNujHjKkYyJhkD1Emp41iLW/oWQmn
Km1vnAK4qpsmEkhr0CTcydxCZHpAd2QLrcXCA2lqqU7oarW92IgNMegTjpflxOb9
2e0bsWMvQisutYzZrwFflKd5sv9kMeJQPPc1woAFz4oCQb33vamOB6XUwjtpRSqP
OUAgj9L7aP7aWGEv7lwP3BVCmxBpHetLAawZ47OMexvLZ27PlD7/F2Hf/icHvz3e
A8sEpiTXwBTAjFZ3NXTwbxUxUC7waJU4dlAurA5RsMbWrucgf2j0qtR+ofk3W69U
SeGebBFpmMT5cO2hb7eCdkWfzYfvvlQJEzg49Sh9+tYIHGRiEKnOXd7HSXcr9+yU
bjHHCtodnkx+4wWxo3lrKOsslqKvw236x7a3uPauFOuw3iXVO/OrpyBIHr3o8Cwr
RLJpXmN5aefIV+k8KR9etE1SOBherz7HxnrvJyvqwbAWyuDhUHXzz0HsGnxqMlb6
txeWnE01A3gBVqHcAewnph/YCBDg/l3stZTXE1uuOEr+xO7E/mz5SwLPpaZkbGfM
5EVg1Hbx343nM+9Dxl8rYP2j7YZFnhJEhdoOuU1oLQBhydicYlerPODabg/D1DXe
e9vx2F1nRwizFR3sv3beNoCqqnxk0bAciSXguu3jIa/qL2+Y6Zv9zyDf7hJD+pbz
gkIKzzHJcxdgo/LtAPEBbPxjMeUUEvSM8MsJEJo08fd40p73eNcCKLVw1ABqNQ/q
cT4fuSlQAwDupBNWJ/ituGsukiBhFIQLN3LJX4d/+0JG3u9XbTTlGAe4wS0eeRfS
c3b09afoQc9u9fk80rX6tNmTWPaf1qJLWZaSkqvEMzBPclWZ8aBV75x8ACUTDKTX
iAzVdEI8uJE1ooKMVTFAs9ocSboXdzZmy9LLvEslTR4lDR0CPQJRhx2mAdjxSHjb
q2Bx73wQZ9p8tlhPLt9ckRDD0p7hdpl9Ld8YQ+iXKp0xI0xDPIsASzewg7sJAmTo
KIbqdULAN+GSUD6mx7QUMUkSHVP93lTYlOVFRtlR7bwdLQ7CVfGKfwr+o4s5ivsR
cs6Ynbwxxr2pOWHbhhIB4tzcYCTHLkY+1lkEc7Q7bkiOV9RHb0fuCJDqizmke4gf
WY5HMRxD69X6OYBeAnczLHI9REtgWV4d4DzjYzSnSm9ZVW/p0bmF3Ufo47BGOTml
dE3NVdfPVgZ0F3IxTmSvLbjrabatnyHxb4EqXUW21gI4XvsZgh3qec+aKzJxG67b
ZUkBiRX6ExCtI3CRCbU9Q9X+hA2v5qB40HE95dLawM8Qy7HBZPnx3SxI/lpgsUEj
RiWS2oZk5eRzXJcZxpC2Ox4ALN3qW1twooa19pvVaHqbv4D3iTIUcN8AvoItdx1X
bnKgFpdJYz8H6a0/RGtzd8r8RTu0Yt0stV6Hkm5LKQRTqzZZVYARc4P0tTR5hzvh
uj8fMoAnTQL3Is5xPiiixfp3XH2lU9uIDTWYA47uuXEit6GLQaWUjqkZxZz1DwJU
T7KPHcsCMyi/sjB45J/txLeTTmr8iUvM56VLw0GAgan7GlzOQPi+fgIgG7PuVILp
LC3i+txByG1yFti1qRiQhttC5OFqphi30lfgOaFFey5vpKEACOWK9yrmF8CAqjoG
V7gnu7OV4H6huvu3FJZH/DE5a1IEX7D2w7g1JdYeJqXeNLbBxscZOAuey9dDFuKZ
KNG6KxfUAXg0vP5iOsg4jXnMDSIVU/sSvgnMZN6ONDtXFb6RX6tFyOOSNfu9Qtd/
bpvpFzcoQHLW7zA4Bakvrm84+Arp5/TpnCqfWMlSanJ/jP1iJuVy+hOhkxz7+rio
2vESD/IqIbmdIPWW5yPaYqx7ZgEZJQypytvx5zbO0H3PY2Rzbx4v58lRWbtAgklX
d9j8+1umDVxysihLHo9TUi/BDYtsuxie+DDYmSdzKy5E1Oqwcto32FJgF+rP89IA
S2vAvrTiOlj+a3x+7rMoFefFjG1r78zqZf4rGfHFTLEHNpaKNsxun1N4jZVWK80G
wKyr80B1CTqvONuu+sn/oN/tPf8FtUUp9BD3C1P7z9K1uWirrJFg0yinf+i/JOqZ
Hm8BDi22r1uWDX6QPUAYOXHw05L0D0L3tMkJ+GM06B92zL7RoCswyMClc5lrWpJ0
K7/FMP3c24dZ6IBm5GTbfCVPUEicLyvhHTsvhvvePpkU+GFcOKyKBqyVV5hfWQmj
YhDhBEJP87n7rhuGk5G2L278AuH7BWUB1oBfvXZntSLkXMmbILPHLWOoDXaee0J1
Cthjc095/GFt01tCrdvXRxmvdj2JRuK/KFYap6xDF0VxFnZSDuQJ5LfJS8pz/Yg0
PSkdVh5pzMUCtjWDlt3Glf0LPd746xgRoCMFYTcwctSPOsRyrkhullIeCFiEFti/
Iyh134KK2hAN8FdIBDsr7/D+W2jJwlnxpsaNzmmMlKNQRBemVn3/TSQRyHK2Y4GV
TH+C7DulaveunwVwj5UhHE7Hemw5jozdA/4tzyfiZwdmRDGIdgznYATfZG2KOZ0G
BxjKNtH9ImBiK9RE2nPA6/UZJORMeDe4r2Tw7BGU6KwWGi66X/fuI+T6NlU2q2AA
8SL3oM+C3C2iZfkPIH2OluoEa+MqvLqCdAAPNV8OH56rhO88xgfEY/gOJrTiL06y
XGC6qoxzQC42Nxu4Z90vw3o/MkX86/Fd1YX8uhnhzSYAQ5EdPP3lUzMFiGUnJFYi
9clYsp/kAs10fs8kOvqrXY3kkW6Zo7A0lqisau9FaTABwICnj6XuRryRkpdnfCmp
3uA0WizmfO9nr2kDH6pB2M1a4HFywDpBaFfE5VYILU71IRA0YfsRUJ8lkOmIZp8h
zsa7rt1sjofwEedoaawANsGHWCEbuYSkCWJQrXFT7UkBpwZaGd8XwrqEvbxWCEtJ
e+CZOaA6y1pegk6oxfVg+c4/rjCbzdcYejdi9o+0peHLjdZbt16RYCIw+YjrAsiZ
c7jrkRcbNhImLL2zNMgKuXKEycwHEgkQJcqMjvP6PRSIji93EQ15DXNRXqDsy+lk
HH6rdtZKbRYoal2oRNpDMR/blpVRAJDgKNyVs8G4pMR7/CiPPX2z2XTU2Ab+G+VO
Z0leO9s6gPa+wvrRTlm1AkmKdv8DKf3R+/tTdn0uLOp4kW0RPN8wc+3HJEqvPjNj
sZbsLsIJZsAdVizcTwmQ1IXCsKnQ+aT98K2ORYNu2Mn39dKvksSzU9DWGGEq47Z+
YoTOCoax0KB3aLRyM7kAycdHpWxdHY80ldslfygWbJ0F+CrRE+BVJ4i9jOok7ena
ewwxLz1SetdGE18AsExIqskBwxlX4FCqG6m3w8D2/2viAEBSLFcLaaicn8Ov6YJx
6MqZoDhfache05BiRlo7D3Y1p4H7yWxQGW8+UDbhlgHP9Iw3KhRsdasehkEZ9RV0
Sf7TaY70eXIuxtf7L4/5Acb5cU0pCeW14fcxMA5zAKpNzHR9llD4gcaCs2RZZ8ls
PMQSFLZiFMqSckh81LPgXzoSsa70QRUkRHH9sMvWU9w/968EEjTe0Ku2P/zpOjhQ
TYspk6Moa8esizjhnMK7yPT4vvAOQLd6AOjKZBzDIc0PWPMinngMKMLqJObTv/Eg
k2K0mENez6Za2sEmioYRTgCEydZdIehwjjxsdyWtS2ZN8BnqpKE/voYf9od1PUMR
lpoKeoLVJ0c/Yw0STvSamkwH8u+Dw7bOXRFnWNdf2hFPXNUDFpsMk78ipghZUVb4
jUppmvhxyTGprOWbcxkQVs12IdxN+T6BWfbSCxE/zcruMvGnHdcP7eN826dzFDEq
evDDfdQV/Yuf2ConszoGwmRevddO98cfRhNFJeuMTQMmO6DGxDfQSRN68uwrTKka
UR92ErNCRSMzLWYiS9Gqiq54QHQaQCeEfeGtUGYLy+0DcLzmfg+Ht3FYgssO/gbF
AEbZoH7V6NLT7J4t1PO4qfNnP5nn7om+SMRlmeOfj5rwsNLIzL5g77neN1nGzBc9
Mz4ubyoBCIZsk+2n5dtNHcXRMDVrY6sklsA0iM75xls49z706qowUheVqfDgiaG+
9vSUKRRGPhegINf8j4shdxPA2O6v0yQ19+0BcZ8+qeDyeiL8+G5Jkm6yKvSAkozl
HIaNgfOx71dKQS9IUNY8nskIi287byhnde2YU2rJ8ytIOSivMMFHEFiSfgnV3bOK
CRpLycbix270ULxI3b4eT9EVs0IhNtyBw7HK9ngn+888PORlu7fHa/1J1uZsK+0L
pkNxiScoN2lLKtMU7mqL6/EoXoOW7+pEXBidabQ0VCxQmP9UV8xXZXk52ccWtfNe
WeNolhgYBh/COo3K47+ccNPJ8DPpRI6AkrlFlV+x3iyDIXj5xPobmZrVZodKufre
ro8ixMjjcj6N1E0stPz0jYO1evI37an3NPbqrFDV80YoIZWusTWZ0IX19TAKnRsx
Ycc+7O3+RuOOjGcO+m9TCTuq8Ir0FVu8rULZVfXyAqUphuVWbCf9JJTcyIJUHK5U
sx7K41hMtgTER9byYa+htSmI2VcArM+x0pJttyOJxE71/upaE8V4fa9Q3RHBOQmn
LwCRb8/FlBX8pzcrvntGQGQ9qWK/hQN79wwEFixcOF7SI7ym8Cb9Xuz0yiHPj/fP
tvnc1AZgie3QrADZu1n+3+xHcItw3wZogWlN5lc/McQMe/QTCB8EBmrTfX5haTij
LFWd5h+BDLzdsxjXr3aXexjLfS5fhOWntY+QkpF2yjqdl6UX2Wcgk69H+ZaSJxIG
rHlLSWaLeC1zy828vDLPL22SjQ6rVokRiimJVDYRvABiFGBoonNN7wVfBMgYkBYO
JUg4m4ap9XXfY8X1AzJfs/5eAftvSSlTdFPnVgEQ2vqWkP4jZ7jN0x130X9cld7W
Zd1mPjzYysOyiQBBinueZ0LGv7zUp0t8nFOTUKDUKxYGBHE8i2iVYHhfwAkSPHaC
5xlEMp5qXpA22Oeg0xUUttFZ2ncWZF3s4mSOR3mbej4WplQ5yKTxhVFogNJYh9+w
MCwghzixzgnj7QYehVujpP7w+qAWqMJtES182focUkhozMwXSIGYW9eRRaX5SdkR
I0FVvrYkT6u37mpuM7lugiG7cC6hXwT643I628sQBOOzKArcND3jTS7218KQu+kr
xBFJXxzNl1TO/5SlBFXlQAJNwc75pQSHNXcKLHEYW/DNGXd0zMdx+JQVtQ5VyI+M
IXzbDEaAl97RK2kzQe/IQzzc7HjBFYfOwKwqs/ua1fuiX2UdDI50dACTD9hHdg02
AM0NfVt6d7/9QGEAzKO069/BPU/Bw5ENLUXQza8Bb2a4hG7iSa0Vbp1k/C4oJZGx
CUOQ+o9SBVilR1S3NsuFHpsrpzOhRq3iLdCedn1gKRVDAx8WicgG8X5KJelTiTmw
rFCLi6pbdfV6Y2s6qwc7vFpDMv0nYzbk8Iu5/4ItcH5w5GEDxOsHZg4q5NvIrt1J
gbO4PWp0c5J37bPwnvEOtJlgT3hdhrUIjOtkY+mqYBGaZ0P42TJA0/TnFafCJQDT
QAXVq8Y8ZACTYcb+OQagJOJkKowe6MkZD03lus/hdvzk11Ck0T9qbmrCIgOkow+x
VnxS9h8HbwMD+ADzfc1Oy4OK9R4Du3X0RvEQIRhOyQaNeu/PjTL4thYLi9di1KiS
tlF1b62jyn4P5JYylMZ16zL+Twb+YeCBy6vYrKhCaRr0xsbMMJOC+jg379leYWq0
JYobq1eOlWjBDvgoQXA+eGh6FG82spCstqdnkrCxAajdBVmOTjIaZmQvHAfhOylD
YnHIZKWAkrJyGHuI4Vy4mm64oyRh19woZ0JzcQUmRPaOBPW90lKR2Oa62uGX/p6k
8lIoVzLarGDMuHxCAhE69ajld41eARwqrDZt8ag+oNQ4sNV8XWvyqx4Vz9a2IAd0
h4XOHe2UECjb88XXm3vYhp+Oa6RDcIh4DIDkuPvxfKde3nau5U/RgjnenaFfKXG2
86R0yVNoXXd2lj1Opd6vj7nAdyMvfOOPgBswFRsCO9p3/iv4Ckpojg6zema7jnUe
9KSJTWa2i3t3RahlYZFOfbEQhX01i/GDt3uR4knKlIbo/kN22pjFavZsQRUy6Yqh
o8w6aLpqLI+meNcfSJMRx5D6TZQWXSoPLG/gCx5Ikk5gSULm4nE2e6pE0ORbk7bf
/sFR/+8ahGpqGonT9GrBU+foS+L+Y6o+10DNkccLT/O4jqJ91kXA/Wd0Wl9FlIMl
IYkTB8bTVr+nfh1CmI7VlB9exN02Io4cuRw7E4GYEfzefuAG9gxRAVPk/JMGEId4
JB3aboZ6DxAJbmym/Pc6NEVFdgdOFDciwZ0EX4Vz34dgYtV2HuQv5600pekFsec9
pGgszKJiEkZfsMoWpvytLlJbnu/DUTat0FT2tDXv/hG5qTT1c2qIDrL4ShQOySpP
Pvak0esmdEUvC7a/fCwue+ZteeT/xGZyAhx76YLECE84iCBZkyFO8D/L1p7lsgmI
9e+NLrZ7edd8e5LdVeNN6Gs+Xc0MMQQHZACtycuBYqqiMjjY9eRPOnFdgaM+KcGt
UlKwMgFbHBFGHCYOfQ1Tl7rYfC07LjN7xWIoofiq1AZ+Ype+TUlg2jnrsW5W5Won
uyLCT3oBVfUJceZZRzF8ITV5PULik7B4EvdsM0s9Zl9+0MmPdnFHbB52FL3AqxAc
+cLWZgsGrNrr+dTnARETfziJYo1YCBKuEpKeThVCZ02M6jyq33CPjhuC1jDllX5W
jBoA+TKZ3AoQ9015Rus9tDRADfJ+epPrx6AuxaHi9ootKJyORhxJv6BgQ8ffwbX7
YIJDMZqGl2mdw+mRDPnKjKsQ/z+llSjdOO9tLBKfAObTze0Mtw8pYqmI5WYwpqKL
68DwsVZiaujQYYLFZ7PScuyu3NEgD9Fwi0Q/nHLiluwewLQwcKaP9cUMddsVL3/y
q5SjlaYYSWey0vYYNfzrMofh6RSHEgLFkOfqScbNrskxjBgyjFlxYv7YUtb7U4CK
caqC2ldfsrbj3+9AvaFhhljvybGtc5nvTgjXYqaXnnpIMzktk0MMJqxTFROVrKsM
HBGh4rN47RbrYR2d9lULZqSsiTk5fWtOjlTLkvUuA2q/ZnxxkJmdcaC4nk9JBEEi
k/zbpddJEjf6bHxg+XHBKj19A19KvNIwnz//hAK0LU60qv4s46Bb4+CQjEBpC1+K
rfyPOmbvcLYHDwvVV6E8+N3wu6HL7jGawtMFQ3sCe/ov2xXfggmJpYEtCjXLKLot
y1kx/YjDlKqI/4GWalyRw5pRURhTxemfKNoyhTg668R+L7B1LlSNYufIUCYj9YlR
O0ToxquIEhlc8vfgEsCoffNHCUAYapf8cmHuXIXbxtiWIiXlDlFBiOOfjq824Sak
/AQxHlK4Qjjy2Pwf8i4SPwlkjGzeyhromYmFaROIs4oH77y94l4fhA0gL01+9tSo
r/0DXi2bEiG520i+6joctPj50hygeDps0dkPQWtahl6aS3M9ewaQyX6Hbo/3OZgL
hy8Hza9rky7LihYbvx6QpHuDBzLwqGQ4Lk14iugDWtgM6/OHiPtWvGVzmz6yDm1A
a8QndK6Apk9FxW8Rw6MBlo+nShBpy4czaU29bhx2Lxj8LdqmF71BX7houfdEKwOf
yypU3yBe7Pv3AqCULpP3GEMEX76E503Yl/Ao69pNirIy7HWPoR/Y9x4K/lm+0baV
+lmvWs6CXxZQ1bZ2ibDGnLIKxDrlvpTWp7tlhsBy3i89IJ70AVxykZbaiaicOBFc
AOYZwQAHoT/QDxIRtF1LsjDR3bpKI7eOt3YbAi6HcK3LG862deH6UnVp6zKpRYqa
exw3AedJPyaarcn+Sdr9OUAMzZ5XafwuozSxtLPXg8kNKCpTMRl6Tmc86TyaB+q6
CErb4TRlwSBa+Z3SsLOy1POCz81ypHLafGv5UXn3lTdHBIFZmQvOwEOkW5PXGGnl
hGBUJLU6uMW7hmcck8Bcg6bPzC9NXc3oao6TxobW4go54nD0y+n3Wl0um2cFUAT2
Hx6SC0wIxYlV11HLk/iv4sLpnxM/WmFsVnZbBT3nmbuV6FLqTR/nq4kiDzPZTY43
fx7vqRUgVZZvKMFkp1xFlAcKlRDVM/ORKSoifRF2yjOeo28PX46oMHLc1OaYiZba
xh5jE4sGfLZyeH+Dg4mn0lrs6UqtHJ+P26TG6iljm/ws+Fbaxh5ARzjESNLG+EQh
dnha6k3mFByl6RUUEifgbLfVyISDKhmtxe2fKIMmuvtj+/dgjgDgrj+WJI6En/xf
bXNfQyzhcaHlsX2KnBA1fITVKlSWQHBQrCC3CRQJUkA+yAsRxtBBopjriqgH30eS
lcuYHD/RZgo747SVE1jpRPjywYFTGlLPlGRNktzNIWX/yd+sx8gRm3Xu2At8mkZD
S+ORMgUVxw5O3OZnUH0bBdqk+k7yH12Lpc+wmBh8gtakn+s65xE5WYgXhVUXd8aT
hlRuk9NfWsjoGgYt5tDrw4psEdPW4zbp2lJ8fkHLdYXY4NfshXASI0hMLhisBoAb
QLPo8Flq5DFMboqHz623ietAGvTGdGHinWQu0NYHsYMTiRyScJsH0ehqL8u3sO5r
j6TCIAqbvOHnrBWn7T0M9HK40dd2xyndK0WXbLttHG3SroFmBYNo9XsvTiFYqY3e
kQ9gFMm6gYjBBGOY+PBHBDSzgjqR85rvAw9JjABcYwCISPL1NL8XvaFgzb6DgyUh
YjbRyuiFO4ewSTB+pXUBvElrXs8oZMvNoGoXS8Os/tDJ3VxbiBRRjk/TBhXcTrNC
ZanVCm/JWJSu8SYp3pQ9No0mi9NtUQAAdOPoMPtxc88t1C4x3FQaUyPTag2CV7aK
vTqR09UymAKlG9pAMeMOlT9YtWT0itClhTTP2ijD1moU9n/K0OFb+Jeiw3SoI1lJ
hD16IK1IR7jT51gEQUFTzL8BHUBAYNXpgiZtqaC7OvpuYMwudpc+20RO6lcNCKDH
+IkaAh8gCwjqLnu3QCekn9qZOUatAMNem8OXyb/98rr37OatdACldW3TM+f51enL
D+dY2rPqO8B9qh+JDTmk0HfnlXMTMar17egcDfN6kXfK7SFc71ftdFEsWpt92teS
AP27+5WmxVUtqreNjVUvvFJ/k35sCFTEeW+H5IMzDERvDhMfMyuigGcn8Y73wZBi
4rRrbqsTQ9jCDmbBH2SVagSWDTFmqWaQeMOu2e3cRco4r1pBEkv0IFuWQuwKpqvm
LH26ETT/KXmS6ygKdbQJtwuPjnB1OxK9ROeJ6j4Q2yrmageyVkgb/rA8XrbwUKIL
bVEtGhe81KZ0Au+OG446AmvYlPLDEqIXubULKRZqnkyuMVH3Ltqo0XFVbcB9dDww
ntQO/mSyZnE2RZRKBi+UczDPn4djKRJ/UidPxEV1ecGVbq2lhMtA/PvF3cEn5XnO
1VVSrifrfEyDcIJ5ZpGWmeZDnRmSqNgMrNOWqWCeinvDimNKFlsYOOCm4FD7bfM1
xld0g7no69jar9H92eyv3c51P10Ik9vS7gTEqMxW+pNt0x04TE+3d7ANq/B9DNln
eWFJG6CWskqNbNavKbumv+X1IWU90A8MYZCcFhcCoecuiHOLrZ+fLpcpv4Bblr/j
Mgm9akSVk0R1Y/6jCIiCdDtW2witdDqQYJ6YqOn126jd9NXgH7pcUUwGma1N7AOp
SODyvy08CGJULW+8MOxXDpWEgmGQekBxlbSXbgMpNaXP8Oo4cMtjB8ECA8fcZEZh
wV3p+bvoqYDBA/ItqflRJ8TY4hmZ1ZIW6GQbPO5i8NtUBHqoFPiwbooegmpjOj4O
XzHu7HPK4d7Lqq8vkz9dAUpp+irNJuuTl+hs6ZrziJM6cXIngyG1ABUmUdMOd5LV
c/qJ8Ttc3Kp4ZvlE/rh7cFR5Mv/yT0lZi4hahNtpnpznjSc1ZlPkzSfk4P8cDzr9
pXGnnVqdcxyW1Y1snL/xblnH2pOOTKaoOEfcrT7G63JCoDEKe7CjbntQYRb16zFW
60WDP3RMcD0b8vLX3BHZq/9D9diKWc0tvoq6MGO1zebzroBJ2ZA0cF5zSjvav+Aj
ZoiylSo46LmjM2JbMPosAZERC3PVx4yUUe8yLwaXsnspLrewdYfwT43EUeaelIhe
OA0C9v4ciQhbcJKi86k3SgNIJgJRgNds491IKBR4nM5kPIlgBkp6bbXa20ATriOV
b9fpsS/ZFBHWaVhkFk+JVyC2j2XTMy4PzWTYq+CGXdZDiYmjdyD7zUuITqnVW9TO
UL83EstLtZrmK+cAAdPUDeQiRoPzVVtcyRxE+yo8Zb9JGjBVl/xMQPy+f/XyQ8Es
yl+ArG9CyY3kmuNbo3wpfJ0jM7qUrxXx1kfaYk3xFSg7Cp+gIOfUnca8qEGD1r2b
QdeMkFd0Qlo0rEWcpNsc1kPlTA99in9ghSVHJu3oKBxAwb/PPfVNxUDdIGaMgGvV
ZH5IghdYt5Aqvzlfxfo1X7OtJoUns+vto63GuxbAfhzGVF16COXV9GWkhwhg8PSR
Q1ZvUOPvo0lWLfhly0QsHJ9nsD2tFpeq3CH5TDGS8vlIaCcqeJ0SPZTBt3dihywT
Ide3U5rCCH0PIDGdMnKN6YZ0/QDzClvX6jwaLr5KYEvm2Q3WMPj1XgJt/J6XpXm8
50q3iE7Ey84xdcEeUCJHakcOwSiN5lZMQE4p8JQWhF7AuqrHIOH5bIcjmEbXUOHD
0Of54K3AohlKvE9dL/cpNALyi3zmHD5i3/ul49SA2oPQHa2HWg5iDzAWHnqDadB2
tzQZ2jl0XsegPKKIjXgSm/2PSJaNoysaYOLCodHrY+sYa+lP8w8AkWCBSJN9PTKs
zfH2pDvJ5flTnLDIaNbM7KskelfPkSAMNcZdCXJ+JCJ6zEErMuRFO3JqCttiIw7G
NSV/HX5IXzrvpe9d2osuvMXVVYoEjjb9LSD94few879IS9wp0Vm1NtEWZFtqSKGI
KpBMjnx9duUx8i+xF6UoQ3lB/7A6Ew4ds5GCseHyLM/twDtQSCrcPpX7ib6C18cL
+2caIQR/pBwaynt4IWRb+PvKlsSAJd0Rg1qyCJJ2JdwGH0Ov7peZJ/I8nNFSvlFU
uMWXMR2yebcO3xMmfZt4LUfkLdi8oqjp//wfI/wCP/s0PQL33Oqvs4a4FQ7AKdna
vaJeICwAOkGTGvht/R1dL79jzTYthKmTjR+rvkSVUxj5loF+Rtv+OVBw470WvEJ1
UfLeifeqW6FSMO9/DgxKRGO2yVOdeYvQBaU0qQuO7tx5izsmiGe9uNs4REGx4Qvv
LHRrgiviY3D5Y3+kDbngFyBjayC/l6kObU7uODYeGFLpyA3F/w+L8s74PA1+qfwc
7BBa9Gu/kMjIz4s/SvGui7khIahplZKP14AIejt2DHvgaUQzprzaeBMZ8TMICAiX
004gcoRSgaEaZDisknBAfORyJ4MzOB89jD1idxutLY+S7hA4OGJZrDPJWVZ4LsoB
xcjjgUFMLP3qmhKzT5LLMY2V8qB4s8fwRIwKzTYEXp2PDd6k7Sjm93kKYtA5e36/
yrJedxjYVyC2Y4Fq2408f+Bq3g40w73KZvwWQeKfzwEU0s22BLRowmIk2ZosPTqv
GmrwOlEESILS4bhqmgW1W+mpk1ZsYI/8mduAVPks5+h/aYn7GRkn0lXV0aoRakx1
t6ZyQ/mNCUxGnUjywCfZyihguTLuzlz4T0q0OgUL4tcfkTAt0x6f5PnVg/8Ur4bm
0IAaKobRrVwf4yz3VjS8iWXvXqMVc80x3N6sfn+Xvvo9aqK3cPIY1s5qvrdieZD4
Qs3Toy78WaRcVAT46hQBudwsY00ik+rWoWZ6yyl9ZkfpYtt2czNIDyyzakxRB2Gm
M1xnR/iK3raiMvsa5wrUgke4V12iAAbc0xMonO96+hFN42YLd5LSshIfF9GJ59yk
TpJtHQeFvcFmthniDMW5sQSe2GFWl6pjaZVldbxv9crUvMWexXBAnMezYB4nDvsO
VLcSsyoK2U47n7qJTi8ySa91Cnzo1Kq8eFiLI3t8Aa+KpMwyZ4O6Rh9ofGbmpX1f
SuV3D7i8Fj2+ab1H6UY8ivVNLAFxMn45hN6bVNWP+X0PrZnyFLsAmU30FOAJUQf5
26FFBNKxMl/CznKC2XqWkaJ57BNetIeUXG8NkI1+W8KyWk8JgedHC/cXHVo6slYV
jyZUE0yIxMVylBLPuGwNKY56AUGP+4uNsWnmGKOEgm0NMz0nsPaosCKY8YU3nUcS
gAD5LTm7Ecb/uR5Cq8eGza5FHOGGLXyOvuLCUdlbOKkTkLErwnpPWookryR1PSQh
3uMy9BOLBbZhlSl5/WvcLurD+tqFkSN52HCnHXXEmb2Rvb647pagaT5mmUPLCL2g
fSr0M//eU4R35dkek8VRMvoqSAi2JPwTZ+EDwlOmH7R9QfkvviUsIU3cSPZoNZ+d
gQY8ZRNYOVTOpPeb4hrQKPn+mBNr2xBpGkNj3n0b0aJnQCMr1BnFpZKJLvE8OapN
67zWZSZw+bbC2Ptpby6+5c+KJXaV2NCOzrkO6JHW8SDKl208LB/v44LYoVME7TPi
zTmMk7FhyLDzWDHmMIK4Mbm4uVz0cGvZCotQYjrIEiiX3wYU1L7zulToOP31CRjs
CxZFo3U6pMeyIzTUxU5MtDI1dMF9FKEz79Tuz39RFyx3Yueq0V8akVSqn5NBRepC
a6Hsb9nalRJ7B0E4F3lBwcdHjx7XO3hRxCpawIuhGzl3CBf1TDtokhKQEMFJ3LuK
eX3HLux3V1JbiMRvr0igSoprl84NoyqwfDBE+p8acEenW9MQbfJMr2KbeDEsDcFl
K/Jyd/nvN9GAc1qRiOv/lcBuSI2pvGgd9Jl05Mx2OfuNyFE9oaANWnYUxsagiceZ
zENyAy8xUQVoBIp00kdaPZLpy8FrprWk+xFAc6mQo+xgzQ4PpUF7icObVM3206nd
xtIFVyp7Cwo3S2DpM9hBVGeveBUZHaRlw17CzbY7tA4Yh5h6GWgyp6i1VqgH4gM9
mw6KyZx5UQwnIhHApOdcrt8/qc3LDqSRVyZ88qqHtfNwCcWtJgyaNWPkgWioAKMB
qhsJFIJnNh2mZsC2QYZ5MXkPWjtLB/yTulCr/vFUufkZgxhYlKyNkQN0Rx51QFUo
ZPZLE1LHHppOPVQyT0gssPywcT2ReBZuK/wg+LoSmlypFLWwpXcpUiKRus8fChEe
9dWfLaWBMe9GQ8OeCdiIUaflH3K3uyZAHDAMiwQmgcTCMagSdTbROnHW6ht3riP+
N7lNmdkLdRiAny6hwmHlsgPOkU2UxmHUBQx8Ok1Ml3ieJjwu4vgyKHGFjd2iTiC/
8lB3yC7tFTz1jbZIDC9v1BbX+yS0qpvvsXSpDS0Dh2nNjEFkgRGLzZ08oFzbB5hb
Al2ou2kz1ldJG9ivahqgmuX+ZuZp+b+uTPw+I0P9H3uA1WLAeyM0qOgw1QArVy75
TyXcpFQgEV73oGwH25na4HU2TD+ixwMbHeZ0VUF1umdnpIXW+LJVngzpiEfWGjmt
kz58ONvA0R6uawTBolbWhVmzF3IkzLgMPla+PqkMUiufTCeLmBtu9pC6hCx3ud5/
m2mH9S4Izv03+PZtt+/ZMv/wQOWuKuAmpVp04US1nOdWfYBdh30J1gDlK9F33p6a
cQSt+FF+EGRuMvKPEP9XdRuhCGuvEat4dkElQGDx/1v6pu+lLxKqwr8yBw1y1FIR
CBytmJr4Ijv8xmk1iEFBWb7x9QpT5SmzoViky8KswDVIgRJGwM13sNnwoGXDsQiO
HelzaIqGlneDVzw44V1Nfxgon6yo0o/St8JWCn1Ly+2kVDkPzS76kq2lgGMMcpso
lSZq5/0j7ZzJDLnUbf98OBfHkntbSjdt6jB4qwrESPuHz3eRcxZdPMo5WILNkyo1
KiJM2IZRJMRDt60zIgCYBtuRiykbWKMGnUkyGX0SKRwTzIAiZAdsrTWwc1QOBzZi
89dIXmHUuHWJM10R+4PFuydb/E8XylLvcQW/GYMEDQl61lLlaCAFXSHjkDsf9EhB
w9vS6+AuYPSTILR+XAK3bVAKJfknjnqbsLMK78GdzUUtx/ti3PvwHTVYGtuQKU29
V3VJuE9gnd+W5vYnNdpAZMI//e89AzwFcHqaHrx1W6R60KJCbS5bC4s6dTNjrEyd
YrXvILLC0WS/owHfbVxiHRbdKUXlQCD5R0kOU3kUjE4FsSJFbEchoXc9mvsZvziR
IE8uRVf1aE5lJ4i8PvfKy/QaHkAgtUlakF+4fUNcJ11RJwUcQSJSi2qI7k9/1tRo
gp3C18c+TYut1lWH82WOV1xHlMwMPh/uUyjClSZBsslVo59J9VQa7HT5rLXLeoJp
AUZhs6mNX0FPl+I1Zqo59P9h0C6BrjsSFiQ/3wuhHnFSp4Zji1knI7kkACzeZuZK
M3ZaASWwLaA+u0l6E1EAL3GlcfCCAqfPFlolX15X5TqlscD2Y+bHisLGlKU7V9H+
YmFiVZfbAwUp79FMGGJm9729uRyBnxFHBEQbmubaTEaqyVEYyFGtLdprCS0DK4u6
xnWkI7VmkZiA4E/VWo6ZpqU+ZvHwLQDaDqR9XjiIQ5ZAyf4HHAEn2PIGaiVOjdEf
saDVqxdFtiB1lCOAw8xg7W2GPnf9imWPJzVgy55CvUt7XI19dil0bZ7r/NQ1IOBg
jeMuzuNDFIQXzQbGP1039clU9+bV0YiUkdJCpuYbz8/1C4xXMrLuv4j6qghnOWof
ERdD+jOYFOGI2aTEvQiR89S923GF9O1WXXROtv49yJBVrAKM9ApMZSRq18l1tsAk
GUn5UW3rP+H+oFx68II7pV8SqNcpgzKleUnr9Eaow5U7A/Iqi+cW6oBzHmAXAat3
WuULi5kuvxfQ3+rvJ8g6cdQ7JfpwEUbimfksCqve6DQ+tFBXLnoc6LknsowpkB5b
a0NhmceMumS7cprYhG7DCAnqVRer84U+sgBWsOI+SYtyVbjXE3Lcy4Vg6/mpt1/r
tgV6vPzMs0oXAvw0vjE2GTFLpYAyyIz1d4m6xhGA6gCAZ1cqoCh7+qzscRbYS9FS
OURp6G7S9SU3h8dChs5AMULUI8v0UDbfMB2mx1yJq+HNg4V2Qr8iykZv1wKka+ul
s2fKAwuBDoiDFQXG/3s9GSyJAqFI5MjzR4pA0jjuN2WYqHKcO+TrsS8AYBX+z0Dr
0kdUNvy1JWvv9RUfI9YdXYSa50nan3XJ79qIVVZcMGZzXjU2YTkD9rnb8vQP3cb8
ZeeueJ1s2/g0FB2Kaj9iec66BlRt2qBb9+QZxiWoiXKxHQmv0KCn3TfVMaaYojzZ
2QNNSdZsAQzZwwxXm1Xf3JO6X2xLwckqYb8KjU8l63kAwNlrroi4xRnv4V0KnNs/
fa64BmC61vgujEDLsjdxJ05Mhs4wgV0vzl5ld0lWXTTP+ZqeXiZSEH4YKHAFF+3s
voWoid3SC3UCI74ANvDYoY0ndJcCpPy8eKxVPZyXpS/AoFrmytt9DrEebUz/3pBu
g88OATyQPWvtLpC3ray12aVF1IJmuqKD7+1vkNIOVMjnqfDchG96yJGONRlbfaK5
eoP38cn2qwAYXonKWsa6oeFj+kWzwv6Ed5qTFhPIsYcuvZYfuvNfwTwRoA9bjDTd
nAzr7JdJxaToZqLIGcqmAKkMXBaJ2Bn9CHV8MwSTYNsArHH61jvayEuECADqgo18
hjB8vY5WET58J31OrJvjnDClGm4li5FtvgD11kC189eIlYR+h1r+KjweEYqpseSI
Mo1O1aoT/afBA9T88iWPcInX/8bI5wSzqEeC4q17PBVsYB0PAk3KLz3ErX499KgQ
vkhb9IbgCi+0jA9ENw14ir8VfabIOmdKCx/QZrq49rJCYsOFjSpTNkllKvZ1BWiD
lcmpDZsVWVkAQ6vLJkQMODO2wmnuR/SPeLWbza4On4c6n+KjzxFbke/UxZjkPIMd
4jOUCIPaPmGT/sdx6jq6XmuTBc4a3k9SG+XmOh9Iz0xqGRFLVspvCcaSNc8B/fdz
zl7frBRDDdjIbfy83d4QLjTjx9xSbFX6HMqwfG6pQSK4wQ7+1Uod7BLVRenQxDPs
NKDgdQ/ph3MRR+ygQ0GrBugDGjfnlInP3JycdXX7jEElWyZyVJKbRJ5DnnFkH/YM
5yL+9dM16Gg9rGwcBgrTq66aajeTONy7vUvzObw27/JTxR+rOllwwooljG6Eoz6n
jc3QgtZyrLYsXsdxaC9VxggTEk1Ay3T21MU/m4ipv7jevLpgzhrYwx9BD/Owp7RI
GUAihSYUngdpm95Cp//+z2hct0ldu2qKNgVCuOjglNiID12Nu2s0OG3KAMBxATP5
3+Z7Is9uDbpM4JajnNLHdb1UTXRXuf8/EZHr7VqvhI/QL8qnery3sXWY62zc1S4A
Mv6VTfYJnG557pgWbRhPelOzfcJ668/WVwuREy3QnhQ8VCBt3LHE7BO17Ivmt/dA
6KIUyxQVJyQKW+8ft0uXOO4nK3TcPJZPkWxRuILyONjH31xfEDbCtL92nkSWl3Gb
cSXSU2lPmv2xPK/lMi221YErCcW2d6vdaMkJ3wULYYLG/40XYcIlUVxPippRkWx7
1rXLbdCGRR4KZdgKUQXa+s5f3goQUeYD6178KvKPguxAm7CzrMjMiYCelcl2Igci
BsMPyl0Grr7nYEuYglABfyNnjtFB1zT5Lt68l2W8AUgypcT0cmqGDESwwMyJ1+ED
TGQNYcZYwDxktxwTFm3dq9tqDkDHl2H6E7sy4blgXVjI60CzkQ6ChtpCnetCmebo
JnI52oa1Dp8gW6teuuqtHuOZcNVht/7bqnz0JT2Fhga4wGLLcyDjJld7GN4pBYLJ
cwDREu7Oz5ZzU3T26Pk9EHWIbxqLIcJeXzn29B9oOl/710XqjWpjO9sxkEbyC3RX
XJgZSoxWzqOJmwsgIzenMKbnilc9KYvBJ0SQxqS4TPxa2gB0pH40Ev7yjbAnH4tt
xKKt72It8cWgx77GpcsyoKINQJr28v1zTqxvjks7tnVl5T76f/Y/11DON9Nmavpt
CnWJxtXoG2Ynoy1t3vvaRxbT4abTBx4OlzFz4IS7QYB2zkeSWEEX4yLuGgXnlNPO
4QAQZiMEUGPLS3qDJW1MdjxFUZwdHNSYz9BlcjgPC/YnYjiL65uIoFSZasqjegaG
z/oQFzPB0NIv7g5kkCMBKUCDqaJI1kiDslmnoH9EYsMXOXSV/ENHAYDPDHbQ+Rv/
tFgSR1c7B1WdaQqv6rtU15uiaFKhN/EaXq8yZZbABG4HwnoPz1JjWWe3mpK10kNr
FQSPeTtkCqpTTXxwgbjX5t76G4FlikWJZoEgX3Qr92tHZKPyL++tGSWI+et0Wgat
B6tprVD+RUlzeCIFy/WYKrZoCUD2dvfmLKKUyMBWmf70mBlJUFU7JnoUSyuA6rwf
x8+xPDTr60dxOITfahNf3d3grhJgqWwEuXQBSiASRTAmmoZ3OTtXaQMfE/TUuuOC
+P+OObSJQr90Kx0lrnpWZqn9z+hjRZJu+0+n2z9Fjr4J3vxZSxotdVIj9K38nahJ
QgWF9Pe7f7IDNsfQiMXhRibWe8qJqYSmyQ4Ck3fMBtxmXlGEEMXWNP7bniNH+7P6
2UAn9icXIp7mhX0db1rY10XEq29xZ+K69i6sDNtT2RtgU/7b5cHESVWNYNsTT9l2
jnnzmgeX9wU1cRh/ba3e5wK6H3ik4ftlA8H9XdvfDD678okaFSE30TPRNI3XQYGh
Fe38Zb/TibaMTMyRFqZOCI/eFp4Bj7kvZvWzmO38ZuPBJ98Ta7xSObhnDB4CiLiC
MAIHi8Z8ZyaTdqMkmzSxSlaVNO+s2rAQ9ipjIlWqq8rk9onXqGfKltKGIbzNO56R
921o5Aix4Wm2PxOz9vr6a4VN0x4E8Q4/L7pGEHJEkddqPCsR535ZIr8dscWjyLuK
i1pwPkhcXk7O9emVUxhCy00qWtIJoBBlFswwWDTMObjqpWrXNTaXVPRBARb86AVO
GSCjHFOd/8sL9SkTZvUOATwk/sRuCiPB4MoWnBwcJ1GNOcgtRbeOraDB1T0lGyKR
GEmvnB+58E+VMiMuKDqDDsWn99lmrvZpeB+CDCpPk0mU0FzVyivxU+XnrT9zdHRt
XLI7vxlQpXcd8I654U+3iwbtCcQP8AzZ/p8T67knc7ee24LQkLlVVe8qkzD2qb0i
EJ0np6Y0TG6oWfuN2lrVzh8MkNxMfPKVU9AYRlf6MVs+Owey1OyVnROe7H695nHa
NwSCUzFme8EF9jCqr0LUhM7ylBX1ywQcCP5DyLN8tn0qhenJn4DzBQ1TfnajPSFW
saQ7Omz2m+cnJoi/F7LSfX1wHM8DJ3GD5aAHlB/LLBBZ3voR7URkPNmBeHfrGzyS
X3OrIxStf8Cdbw6jYpBJGcgLwxfXAp1wfQw2v01Rc3y6qUVAauoLEvK/DLlfKF7L
bwKGwDylQ3pqKcDuIk9w+qtq3BgB381CogP7DaPn+umcbvGbqx7Mna96rKgVMQiP
6J35GkZUyHJBeF0DOCMNW2o5JK/ctCz/theHM4JhFs6l8lN6pCyOJZy1Js1oW6rn
l/ovZt/0xmiKQ7YVs6S9LWB7KqCBXxvwY2q2mj3AkumPejzprN0GuGj2tOn9I6Pd
Hju+hqtWcgv3qObAwsstPFwgPcnqlsWddpecLMZO+Unkw4NL/xrYveLxMqKQBj2X
nt4Rj/kYwcl8DJ0cxEdu6hmZOUYxhEKctLl4oZZlrAcH1JPx2j51eM2B4DBm6bmT
zS4oxr6o47nF59BHgdXQaUZi4mxpXt3w9ia5ACvaHvkXS6IjtZErgjah52eE6PVQ
SgOybZ7qJWzbITm3fQXxezkA9GIpAFtuTddxuuVSXo7swWRBL+mt6m2hS4WKi6DV
bu8jP0KtViCKFzkYWbO47cb7ShHO/QR/SONaWE0Xc8Tl/WqNi7OVKhHhgNJETSYT
eZ7/n/0yteOvbBrqlSUQnAwFq1KaW60dvA2JsOTkiwHX/mvPtfRk5XUDGEBbX/pK
4HmidU0R1UUChm6X7nJNu/5HtzxmLrwK3YhSe7enhiLRwTbP+4rDVGvQbT3cE7Le
QEO5kfsQuS32sOxVuhSWJX99lDCAxnxSf+Jrjo6m6qO2tE/8ifItX5ipN5RC1j2l
CEKBmwLwhwjor7y9S8S8DN9HLc8vncdaIPDlPfiCgcVEYPBeKMvM6HYziao0zfEo
pbgYmR7w69mXTWEEW24M+TvhsZWaV7Lz0ptdIlERCppHNVdBGCElQBdrStUOc9fh
IBhRw1TySdktI4MYzP32LvWU1jcGtSmoOWc3sPUIFe2Br4J2GC3ypn0kwn6Kwsy0
aZTdHdE40lrRQgy9qZbxfVl53AUSMYYZi8fgHs0uzQeTlSApxoSHEC6cu6VCFvJq
cRe+3CZpFOKzc1EcFJcwOds6whHniqG1y+jP4sgEI7qdqLt4eL16YTclMRkpmlr4
M4jyWcKK6MGlVOaFxZJH/NBn00Dvur6JUh5U8WfGKxoD2c0YOKY9xLt7mjfImMmJ
kVEfNypsSx/ptqxIpQ4Nn6A/ZBv+RrpSd41nwfCfyFwKgncDHyrRvfcTsGvT4RLf
IP7ta3YJYlY46Q/hB29IIqLIeS4ilTollJuIhP9Y09/pHH95eQssG0jnPFNNAlV6
rr8jZ6LJZwFiOEqEgWWcBp13YRZFN7z3s2VaHgF7tF8oVrJJK1SpZa6IxV24RkwI
PwgeZsBe3nLmXy8gHGZk7qgblgDAxMx3C2XhrCW155tNJ5ip/e6OOQ3hC0bEFoh+
PkpiiefUObhcYLRFJOX6rEKehWj8TBQC9SJaTVU0HsptRy6GVtLsV7t+yES9qng9
f5uN6+/04233CaozpuCag8cflW/LP2oYc2XjeNzfdvdqCnJfB3ZhqIGVSlgYqrQT
5PqQfSEK/ftfkc+UTtdfupvhHtrpCC7/Qu2+1CAghHEmyOZWxC6XFQfuIBwqXT3W
4MzsZ21qFKqWNWegRVxR40kboSr/0GmwVCzOfPxCY5nmQF0TFg9m9DEBn80oFGpq
BZkFO2KcV0qL8i6AmYedAbIoozTH3blROnWaynYPg5w+dF0Gs1WrYhMTSMhhnhWK
DKZrlCl1plUiC9nUrtnprgkhec30W29hJKnMj8x/8h9iShbFtieO1bWNn8zBvGF0
y95x8j3QOVHrvVN2LMUOcu5DEoUs8YeFCig3CHrv9Ewhi+aXBfyR8KdcRHSJtO9L
dONjq/5xcLj0PidDvvdPbWdBQBRWL7P9JhDv0l+tLn8GEQD1Azhw1/cEKfYKJBRt
1HENGbQYSjl4YurqwASAjeNxgQGdPvvcT7jbd253hyBS8NQSANHRLiwt7FMEEUy+
5UJEOBokEEO5HZGqizBXrcpETLiLOSXT/NmeFN/FNWuTsDbW/Mw8fpCQrQGyDV6L
+sqoLxsezKPJVIQAwo0ObKZp5EFuv/0rGvzE453/xF5VZ+3MBL/4SrAcaI1fft5O
SrH8DaCzwA34iYA9hFvg0ToKk30/JMZH0opcrhhwL1+RfGHvIRXkir/SfTJbQ7Sl
Z46pPpHjZf145IzReUAswZvf/KzhbJvsTrywOypYbBA6J1CZub7XbLMlyJsq4yNB
S/tfjor8Ae/Fm55Ox5BQIRtucDh3tfK7J48Gmq9FxAP6jmGE45GcPQx+DuAIWha2
LjL+viEBv5FurqeSg3F5plkzdZppUjluLQUWiHJpE/43+shcDbnTMN1mxP+Aa1ey
DDwCS+gID7IR3xGfPUMgzS7ioXtYa3lMRyQKfCDcLwO5mKEdvWfXad7XDmajY1Qw
0cySpMKNtVFC1WoHRNXfwJOzRHV9cWJEm47P0FqiUFR9wXaco6JNcNKRVzosPyou
FbqtvjjzCXEC4Y7pqRee3WWqgSzKK/5DEfbOzondnRhLEdtjgTjjVUtCfhwC76km
N/1URqjbxw64z9fqWQ6nzvNu6l02ScIhXmWyOrV1oHzkpo1DbHUqnJM4n9AQjVl1
R3prBIyO0zTm6b+wtuNBUc0aGF+KT7D8AHEsoSIloHXF0IpAmpMtV715PXInyz5l
q55XbHr57FKiorvh8dn+KwSSuqb0RrbEXWZ269+8q1zqgbE3luEEzhdJOgLzZQcT
KUonycGYQQLIw+ZCnOXaDSf03wTtezBgalxMMvU2sHFjp/AJC4hw6pwjgWtiE68e
C5PDEARBzjqrDvTS620f9bQlKbZBF8wG1lBGe/xoXQFgJsiQsokyub8MwnbUGTZ0
WGXxoJhHgwqY3tpDv3ZNixiq2mib8xsKnj55WGjFr0iiVZKg/ZYE3d9GieZPr9wj
tDqJJxQCn6s7lKFaTFFrbM8cd5pPWYQuaOSMnxOTcCeUTRkEbNcgMUCEOYGGIM9I
J0OP3a/Rm5za4QdpzcChneY11JXz6aWG3FYXss20rXZXX1ILTgXI5+0Zg2ovBqMr
/gdSvl0ytHY46cIJvwpl9X3+ERL2nyeubcdC9gwWXlZC+U5ZxZ8mvJH9sKCQWwRG
CvHYaxPY8O8otKEbeQ1x/f3MqI/YSFplq/1rsqqrAa8gjtZY7NihpqB92pSt4r0Y
TyPYmYfIPED7h1OOgGEGka5PtBxceYFQGfw96STYkw+MgUhl6a/kkORz5QUbzDjH
lj7AYRJP8/qPEF+xsbUekyhjexIaEu3kON8LU/YMRGlR9X3dOvApjyZZ99AMxd+O
Idx/po+xDI1QwyrqGzsplfG/E+sAB5e4H8IdHP9xSc3Ln5wQTxM1hZ008RXwoHrv
dxZqBmd2s9l/zpZIeTXiYtBDxFbo6ama/15zyKwdQ9tPqblXMV3ZsnPu7WA8KWpi
VCNnxDsplE80kVXgS1ZJwOzWHmibjG01QIkLdREm4BNwv+WnUVWpj1mjnKqU0L4Q
FeFZL1MQBARF3hlB+nJSJhpDq+sU3SFtw9bxfSlVvwl1JnMyAo4IHFiaoNzSa0ai
mgnldPy7XNAAZPTOPwoT4sE1fk6MzfHqP/FzlZlMGibIv39jcZwHVcGPkENOsF/d
l79xd+6zGspBQTETebDIhgSF/mFHAciB+VkayyEcRgi73kyN9zM2OFYWejsWZErB
D89afZ3Ak1e27vIrGeQeW/QDPuucLWgXumPwvD3x7kNaFpfReZA5KoyTV3OZbtKD
9jK5MKhFpd41ePChH76rmFHBYQUMom1F+6Wi5IDqVt6mInI5sL50jRGQJS6et3uE
2oQdZgfuQ7hluFpv4c8MyFyJN0xDuq65viFpFpi0PamD9YNNYoh/+8t94QWCusTF
q95woThNhC3TVMnsOXw1Nzo+XE35Anw6k3wnttP2zX9tWHmJmCUlOB5wozmNg9QD
Kxeu2uk6fAX4+8+sAQF/YZAm7gUFOkVsB7cje8plzGO08GJyfFVaSJb9Rm8PkreU
qMyenk6wPBDI8kDXRhsxALEY8ftdrpme9TGk2WgymPhUcfy1zna9pHHHG6uSZRAU
keu9VcbEJXjsWfOqDQYUEWCQZyz+vIb/qZM8LcSNG3q5dtXiZihs27oUvrqCvRIS
ZPNFRD5JrZkjcxc3U6E4LRe18JZaIAQR48qnAAUZGNAJyBGeC86STWROwSAj1joo
ff/AQ/SH3xTP1PF0sP4MbSAvsITYCsjECOIcyqgvnNWfODTb0MMCTl+M23/j9oLE
i7q7gXr/7ZkH/rxosqEkzaFOT5ksretpl3Jhspn6aUfnQaPvghPzyZhWP4x9u5EZ
wUejknsxpOfqU2P2QrDEZqL4B0h/lenHPnj0E10o7yyPUm/7pV6agwS2KoGOIBzI
cZXo0e/SgRvN5kyVyCgn7w2hLCEhnCgJ+3rWfHWrmI0nIUZXYRjT83CVm2MuQuUz
aUY01ccYVS3GGG2pphI89q++R1kFEIDkjxoEp+CwbYxq0ZHz8gB0z93KJmE+DOGc
Cx6qqKOZT2hGPDQ//lCnwOOu4411KNnABUPtAd7kK2niecPuQ8QqOjgivWOu6569
ff3bcEuVr4h7SDEVRuyK5ZI+zm+gBwYXNmQsW6+rvIfPNhutnO3zryLmpGUcQ09t
8UJ3skPxmv+5anDWHQz5zK9E+nZW9yCQptG1hsIeQ4c2WVVO9g9ljxrs0IYDhE65
YeceouHYdbi8N497Rqd2NKiDGMSjr1JexaNdMYvlAXwa6cytVveH+h5J3VZ9MVpJ
ZAGWBIsUh19qPfR0CEMjcMEI0HapiX6Z60FWK9eDlBqDmWsYsI3exwqh6NitYn68
6DuaA8hlE103hKSmZnapVNzO9fR9Ax9QQFtLb6/XQ+aTJ2aS9YIQREqY6cQvvEWG
9hTnHOIOUPHiEgZUKnNu5A2oE9oS+GWTTk1IaawUlfiQn+wxu6Sg3r4SCE88+cLl
QstjXrjN33ZMVBXAHN0F/Glvmee/jKPHGNpxGYANXMS1sY5sY6/IgJPCgugFzb21
6BByhhy2JE2IK7TUBsvoQ9l6lenUvnqiwN8mVUn1XLKIofqm/ZykwSg5gaUp0t7h
YrXITqws4sXsBcZxJTOZN+yQMpN8bcVUuilXJGmYYqde8HqZY1EkU9hjeVlGQkzC
4TgujWUwSqtVz8ChEQMpdl0NAmD6Voi3IyfMVHwd2BcGhvpvUd+5jxYQque9/gr2
kkHP8rUeeBAVTSP0az1ezJM3D4JGaZBR5E/6eAU2BIF8nJIuyqJ915Th6Dr1QCSO
jiHrxm3DaQcXxCYIVcktbRFfiDGAFJRMJ8Wa5OCcLCIW0McNh+ehH5rSHMvBQ3iE
O8QXrFhVTSWZjarvGnBPU7SR6Z8fo1G0AMMFj37NlhiJ1k88jlYB9d0SwHccXu96
xCw7WqqQ0BQPPRKFSVjtaTQ9c8TCWFETkZx3s3MKMqi2Dld8X9e4fCR0mGzgTte9
WU2bIMQoZe9BhGr1RuAdjUC4ezxcAhPIkCToFcIUjKsDB5nwX21VzeQYmxFinxpL
e44PCf0sI5bj4WpUIXqBkbLklJwtC/KCd7cdKk8hMMZ5amrgnk6r2lbpG8DLmOEw
blIE0SDQ43FVlCtWUfb77peRv3O09xhaGMDtR7ua9nATipjlMpRWX/oa/RoVYMPN
dMTR8cGpcDRCIY9LSpLTqQ9nCIJ9lKcPyHjmX8KFpIemXMsDiHfivoQrAgA7iWzE
LsldwVvFPL48KyuYtynCzXtYljVl8OYDiOcUhCKsAxCyu2d0vTL1LRZcVyJDdFL/
+ZRToHM0g2F/3OnMZq3Aq439gih+GdZR8EKIKNFPHxZAWQebtCaFRki13ylg/pIa
ei2GqsDpdEOEpznQzX+eENbkJcM3Py0y325a+6OLoVjz8tLGvP5ql5Yft7gj9SBo
TxK5ud10gsyZDeW5lOirZRvE8QDBUH3FU1kpNQo2skkt/ivM94yhas8kakN1BXGd
JeXv/DvVY6ZE87iXao1IgCIcTSRZAlH22JEy4kAv6OFPJF6YWPeuyq2/evP2McIz
qmvzn8XScgXIqqgEhYSQCHwJmzJRM6SilRFxfPjqTASH66lX37656nW+WtBR+5kO
ZCPbw4DTVJYd4QeChiqhEF4v1Xc3t6LSQZzCRdTEXbVRV7PkBBY+x8WKzAVDtj1P
QIAkGy2aW8ZQ1XVuIBybXOHrjeKefebr0oFbZbdmju1C2whhzVYIsUbG6MxidZlD
GCUtM6vFrAPJdktc2pP6TiaNfk8pABN6h0zQweJXK49uGXjRlp7GkH1L7vXq3Wo9
LSgnRiWm43JGl6NKuct8e9zZgB5xqIREz4D/Ocw+3Zdr+fTmgB3F2zyL4ddbbYSa
5hF1vSybkRn5Wxpc2RLxGygwS6MzQwny+d18q19U55kCkyFocU5+3MMLntbqyNKu
phBxEk2NbFE4jWlx3ckXsaIN+zbhDPoJi5ujc0ylqNU7LUhxaT3ELsfjOlXIGTdP
2KbKHZQj+e+BZVmt5Kb98mv7Vn5PNRyB2yaU3FDlPtu0QiaZUBMVALCcg6p/5dl3
oDM781sOaKqzzVDyT8cbxnPFE277QYcqN1ujUZfMhySt1SXWp7cyhXYmLMi+ysVO
+Rz3sSQ/FPNMlM7WvnSANXMS4N4DMZ4Y5T7dShf7x5Ck+FMZ5SVZWa5UtN8e3sqV
ogbp2MBB2YkJzCqaUaNP7fo5eM0eEG16yiOC6Wxo/DrBT8XFJizuG13NywxOWuLl
WBL2N5XTaCxhzYXpWX0w5rWJsGNMELuxh+p/Az1mVh2HB18gtfaOABGB3B/eX/Qu
moMPSXsvQn4c9oWZzqLy7MIc9jwGbHL4EhNRKv6pc7UyJUx7v+2RvpR/ufQo/W6N
gTYWybCNbihrw9VutsjlIIdIgKKuepjeYLS8vQ2gcJCj/nUddBs5yCmwKxqH5hi+
WafPCYK3AZSIkIe16SYHJxtqDuJh8ZvTC2WdQ9LAonZXLFiSNboIaSav+Fx4pc76
w+4yDUWMl0IOKGEWqu0CZQUl91sQNn/G3n1vRAv51257PMRqPzqhMBMbRnC/IIiS
JRMSMiN7dBMLRFcEPWMSEMeMwh0bxlIKB4+cAi7Z9O+EVZ0qGEqqG252ZGdED9LU
XUlwVY1R1T2cNaRLWoja3uZB9H86ZbL06Gh/WoxNK//KCGA2mJzn6YZu8stwBPpP
C2iPQHgGrOAcCYQZxsLsueO8acRsZucD9iJ277n3oTa8XWdN548QznNKUnDiFdqt
DhPJ/f1CD0cbZI6nF17+4ND5j+Vs0RwteIWyUvg4sONXTJN7hil9bnkC3bMRv12O
l7ZDSV68naW8QjrOtH1SLXAlSBb582se6L+aXUMgyYQKJIy+VQ0prQ4OKcCcOyEU
3vnM7N+l+2SC52A/iM9ZIakVkR5FjlRjvOwZTRkpgCoM6xgDfJOCkgnUeT+j5Le6
1FYCCnrqBoorDL6lNRd+Lg30dcoT3xIo8+OP04LzRK84GtrUk1XpZB4LYx5fnoCV
jextrA46MpW3FyuNO3q8qh5HCUppxb4WXSljW8pHFVMa1frvdUEAO2dcs0YQCakJ
Aoos3v+QPpZZjVzshn6P1zI3CxNQS59w3OskxZ4l9CxGo6znpe7wtJ5TG6Ia890O
y9nqBQfMxDJ5Y6e+nsJb1s1ZhuMVIdPDffOoWGnId1yhQstG8ZLLq+mgRjFDJjiM
/Nd86W5TEqxHu3nhd2VTDoZvP9Wmomh1uC1AcIVxZ8iJnEjix8diSv30oEdh2TxJ
OrXlLMBCIPpTVndg3TMVbOrGiM6TGOIvMLiUU55jHnvZtFCTujnYtzqw8nwyP5fo
7R0cDV1ka/+DElMOjRO+oJN/5KsOJaW/U5WNkeASUabOhCxAXlceLPoERsrApXBf
LsSkG+FUosRWmXa3fCwMklV3haWXp1L3q2DXEkJ9kerSp39pVisonxmXJpPdEhRp
DkWMPgyATqaU8ujrn1leiwuKf9Zs/Yh+bcCU9+4mRp9hB2qWU1o2f1heGvY/+X3J
VpbfrBrAiqH6mWWlJyyqvnLoMMa+fUf7eNVIIR7k2J1JQGGfv7iqQ+jE6Uf+BNlx
A2WmqYZuERkPif5+9GvqtEIym2JNHJe66VGREVG54lTeX9gjjD4jpEVdisgZmeY5
Wkp+Hfj0/9gZWm0qCEQYlXikwmkJcecBIsKNFcwH9D6FAqwXcNms+b2cSZFXZfwo
SlO+51cp0+2Dc6Ts7jP+bPNwYNg2fhggDkcYCWxqksrqMPKD2XtfTiEA+nV+kJvc
lpclQwCEPCRA7YSvOT8fBS6W6Um7oJIJt/4T92AsaUNpijOpz8FRq/PBSLBFrAhA
ChQuf9eWBJ46fyT595k0Voa9m9mVsjTuLFG2CiH1/fQqzsCxf2Sx+ZETIz2U9WUb
AQieyoHWEHWlkuqfn4J/5l7kXhUnM7Y/qzvRTHUknB7LGefZZSlDTBP1ltr86YQC
NtkAqB70yJlThK2SBWCXn1JfhW1E4BpqUVU6H1hyZovZbdQ9Vw/ferqtrvEGlBA+
EL59A7E3wOu1EOtE+O43C55M+oRXbiu2FrSeRRPROp5JP9upnJqsjkfWJjpkuiij
HfTMHBEIW/jRxUCt7iPrpqOSBqjGDNqgSNyrjWskFkcAWB3vzmB9N/4+XZddSFH1
Kpyj9TFrhXz+IHFKLweT2gGtEIOIOwdOVavGC/W6P0v0+V6AQu3K47A6N/LKvjAW
NZgExwz7CoaqXOtsp1+UDkDssze+Ftj9KL3qb8aCeyzyEpEUTusB4MqrheXArdQm
cdu3uoVbvqEWrdUe2M0REJK2GzwgMZP4V/AhO2VhWHx76mrROXBb8qKcjulEFb8m
pM01pbVujmptfnZCYuc0G9jP9tfcZCXZEkqnJlPg4tlKJxoOXDWhxnkMo9mtyGdp
NGhlVYLwrMZc8EFPBRL4vXT7oIQtyVVcV6mxyet9Ep6koZTIPDnqonM+PH/ONjgc
jLM8SvxVneKfXLV5fucXtnuLzk6C00CCjzjic8Cg1ihTDKBpckY9eh/0SuR+0QZD
RIBPwpd9CIQkz9JhIY0Ix7TWFauHT7WWgyp1qSTlUOMVbk/O17nJCOT26ER3samx
1N5BzdL//P8WmJqP0q00Ud3TyIgCxMSQyGtdQXdL7gJRCPS9Ut8t2rJ5waSIA7zr
ZhnpAOLui21yKdMwE+fSalXu6BZVj9EbUH+O9f7WqoctENfYEsTsxJBtAan1+X7a
ThNZwGS423BtCpmya2wJhWbh6W/kbXmgrIYk+c1KcJ8wZwLC8nsdzSbcKDKt0Z98
r1f5TMqDOm23vo6Cefq1SZVOEJzGjR+rGwKdtW8c5575bI2J5TlCao/Y0+O74hll
HZV+cFlKxLyPDGN3l4hTeLGffRIPFK/PmignE0XGknXi5QFHMzk4STx0eZZPIXBT
+DW5QzkdYf70vMmMeUQ3KMfu9hDdfUz4xXuWxxKaQkyF6FL57ZdHfjtOSqrxnOGc
yDaehmnS7XhRlwFcTzmcLo85WKg3nKukbjdQZmLCTFKTuX/t1AaF0qQZkiFHhdkp
6BHSCpG6JvYPUx2vTfUSj4f4VmcfmSrV3wazjCqXNxexLNexBiRUh3OujVaPzRZd
Gz3nuIseXPq2g0V6whzkSSwR6LZoITSpSSFuHJs6dZQ+YuWZSB+eiHWTqlJ+7z5E
iOXxW9tlXEuYWKBWisn2Bw1ZLPmrkhFxJDJlyZT3pNbFsXIAHvMyr79v5nid4KMZ
msVgZAikB0AGRhvI5vN61Q+3oSXzwJ6150R0nxKzUiB/ZqOJDSCATC+wz474Ah/k
Ck14a187D59XAvIVVN1UTPu4ag6vr94CYOUPKiZnoFYjmOa0o6F54zq7bg81ZujF
FCLWUT0ixLukpAY2d/Kr5wyZiu7RVhNzqXt9wOpVTZqmYwa0AQnU++QsEjYF8IiZ
bndbvSblKbTYf9HUt8FBGYusVdDaOvE9vWG8tHsT+MiXOuRAlghjVqEFxM/CjXbt
bjGmTUNAEmksXRJDVpE85IhXAX/FjtwfEWzmx4jIi2L2L87W+TT6YHZ6UMHlTYxu
3uPnNugdVaDLUgvm0Q+W3t80JFTmyB8BZzZPmTvGhkTJ099BMws8VFQSadyOlUwG
rU42O/yzlR/Tplq2gkFs8lUL/5uCRaNYajF6ffB6SLf2vjHig0x5azQCFku0Rd/g
Ya4STWeLuiwkyWPdQTYhWSZom6emcuvTx8SrRuGYkAfAAuZcmpZMxXyoQHVzi4+N
hXSwiAlyh/6yRgDaWUO362UgZjnpsOC8i8N+0sbS3kecLNgyLfMME/1JzoDv54Di
gfnZF3C0bn37u48PyELPZNH3sswTbkZLFJy9GHpY2xmya73AytIjUM//KNGLioYk
A4YoumDEp9Ix2IPGs+Oey97+vPHuy1u9aUEJ6gIrUMwZ+p3U288h4X6wixxsvNUE
1Dz6WHH/B/WOKY5qVmgksc7tx3sOxuqjsXaBKr5U+0YJzqWgIOM1IUHwDJ96c/bC
z1xW83tleCBbRDNp4ErpPc1dNg4o84F9dSWxiGHK87kQ8AepebF5jwYWIVP4F/ZP
WNEOrOknjSIngVeTeK0/xePqcHv2PG2z4EA3WzKmlBzSixZsmA4x5qMkqaMDVSHq
LtPpWI1dUD12RZx4PbnJRTgEyh7pYFSiRD1GNUwMHaveRCIIUug1mMYTonrfKTnY
QdFCtcfqDBTonq46qJ0ezGlmLNXJbSyv7XzPzvg2AphmK0NHMgpPqrk20UgnRlbi
xvF6KCd5ITJg7N8zwebUx6+w0fUQV0Rf5Yv52l81xUfcp54r4eU4okr1Y3lFkSZH
s3qersK90RQTkQt5O1jigXW8hjDw9Lil5oh2dtR1zK2JPU0/GxpivZjjRgzrvypJ
jToq2e9u8PRFL8deXhVG7LTiWkPpSxQTdLJ9/q7kXvvs0LdnmvfB9IG5O9A7MeAX
PuNjrAj3e2tMbAYt1kBsi5YLi2Wc1972+903vvj6y//LponssLTsb5sCo/8WA3w0
/TXXFLeMrFx4YmnSOWia761PU5Ywzpqjz2EbFEEdexQS7izPhOBKDnIyF7hpiJVG
VN3ylRQA3sisgVX+UWvTzLTWGCDKr5KZUrwk9nM+7Yy86gDnzu3RacLKGmlwpI+t
JGLnAk5aeVrJN9YKDhbg+nwhyEww1xoLsSv9Y1FjpDI4rAJr7TBj6O8iYb4io2e6
YBT6WBitzjVfvwhUuu9a5UVLE0nr3gZtkMQwsaSrK/ATHxOklvgCw1CynayQFotL
cZv+/BclVG34EmAaSQtdGA6WW7UEUj3V0Nl9HCNCmlI9HorQ/18RBGZfKXNjFGik
m5MF0jI4oB+O+pGHplOZmpH+wA83rvlzfN5th532RpYQjNKUm20V4KQAAxvGRg/R
/v4Spl4+qcVxtrbY8SR3zt5udaX7iE1TH3sHrFNuRaIyFBCqOZ4r7cgJtr2F0w2H
CiGBtSvYruA5WnokGNoT0ia/hffc1M2/jYWHZTXWF2QciiCN6ZWrL+cj8/RKYK2f
wmdDNbJGwYXR14087pzamEwuUz0xBHp+C91vbiX8PFZLtqy5BePBeaiEbYlSVUGQ
MMrEIjgd4uBrnjWUTUnWlX7A1GOgQvIo4zhO+y9nDmEP/NkJUoxJItVcj4ppjMVw
5511vgzM3tXaqFNjG7ZwSsjz/q7mexyirdjf8PHDc1fR2v/gkj8Fp1KaFmZ+KsmN
1vOmxxt+0IlR44PVphMgyoQdgFoFlM3a29UpmAe5mufyofsfFEsF2hKWH/2Iw8vY
92uFmvw6sPluMDHNSv5vp5AI9bCVWOOxivKdE0mM4axGqvKnHKDeUaS7JJiTUcKZ
3MIhLncK6/G+WIvBarP9EbRtzWOLPbTxrt7F1n5oI9uYuCCx7odv3ZxJybRNdqIj
qjz06OWkMlJj9jT7HdLTTOlklKO8bxuXDLpvaKmaDU5RBrb2prNp1res5fABtG9S
HAB/zCEGHdxvLUynW2aQKPQrOq0bb1TlM7ZZtKpFdSnqc5c5o9QPefGRCGEp3B/e
YqhVxnoutlLmg0xR2MHATHPo2IHzGJyILEh0ra3wqxcmYM2mEnqKUl/iZmsLzEIW
YMTwRvyvOnPkohIBvAZ4ZXQEUcUWKGRUnYlBUwLCP85fL1Mp5x1qHpFmAtQeYWTV
2Xp+csWi0XeKKhQfJe6FXs35rxCELrlhs7kVvvTERLgXF2jkmO1lR7YkJ4nFWcjF
gIxAIFmvZjSTp67rFpQxer8AHkXxMmm5u4nPYBmCnO0ZzQO7ddRwIhIYC5M9Nj9T
fcvE43XvLEfr6YtduqrpT6J7uq3iMccVNyz1Etfnz2FTBjBk7TcF1CI4X/Y8kaAr
NfaMntQ/DqWLd03AKJmInGxxGtboK6g81Yb2jHLI3n4EVBGKy4CGKSH1n0oHi05S
KAO5azttLitAdle0b8SgrUob5vffFunvbW5MlPxgu7bzG/7I6id6nsohxhEnpWsh
Tk+BUkCarhObmIjpJRQbxlVKugTcI80C7dSjUEVj/LwwbrpZhmeBt1qs8Xfrr+hW
9mTCNTVMpUPuGMQ7Islll1cFCheKdByryoCjGHk5vdUqx6xd0Ejf5RUiOW4C1MrX
Z9iWS5Oyrt4b6c4U+38xv6VcEnGYiKA5XON4e4aR3Y6m8wkOMukzLB99uZW3l8lo
F3rVbxXPbHFqkG6DNOGceyHBo33DDZxIuSOa3gNdRSAzTXgc4BM80ZbUcbmqHioS
fagTnr/o3hswps1WIJRP77T4L1gtcqXW7zoI1uX5NggprwtegpJAewsQBvjg7wsl
uVU74ZpjjiGFNjGFtusTfE3k6VFcXxZ+joNeAcyap0cLqheUFrNvYbUa+sItu9nK
Dzp66KaOvPWIkOQ+B7xpd2y1qhPsNByB14Y8VcgJDYdPUI+2sss02Zyl7C1kZR1Y
21IT99hdgX0h1spJCMmrkVvByxOfIGWcD6RyqZm13S387AkugSAvHVXcoKHAAvJ0
5BFGi2MTBtpPb3WCpxxFGTlCVWJFVTgl/nHb+uU+yiboYwKRVNv8ANh9g9QpMh03
3w3KPR/2Vq/O1Co6wVI1WYWeg2bQ7JcgcwdYlD2407/UscgbPPMwBG5WC2J4p0L7
3ui4RRTxNFRt/oDugyYC2+sT7p7YVPLvsZZZe5mSfcHMXrlpcW5ZzDcP4mnqE6qx
CVhmSAk4lXFqIs3Uo66uVYZQqU4q82HK+L6rIYBWS9bZ2conLpQs3XL2dzHrEMX6
YTkbPShJQwEeFZ94/7g1TqQdyXPeJcnOPUfNNe1EsEp+KZg94ObM9Kc+oAlWuOU8
9oIzK9kfEJtWEutXxse07xiltngY+u9saGZYbNMbBLhTrc/CZCwzZsMds6tkskmB
K+d1fX0CLhW4UQUVCHAdeUJRRKGqYeKwYxcRwAK3q41xGENy4mEEycraL/zBaL8r
eefTJoMcS2PBrCTMBdrmowQUdXq+ZQyaLqinwVF4PKetU6GD+bpQjod/W94iLz1M
vINRbBcwdkEYC2sbUk2L90frBcRUg+1GuTGU8BuGC+2DUJqAH7hKUW0R43pyqZfD
ZXQQoAuvwx7ZJLYFPdR0AI5Qxt5nsRvXyv1R4pCFjdxiTVwZDRDoMfSparvIw9iP
Xusgl/59bUMTu0TUBSFo7me5IktTC3Z0nIIRZYzqnGOUZLZyIkSprmssv3jWg/Vh
XwO1atjLAZKuT7rjD4P8byW+2Kjy8ytYRGapU/J6QUkY/alDFuF0SBlBMFaenpcb
/Cze1XUp4BSbFsvNptUdQS+iss6o9AuzIkc9ym7lW9XDfxKHfpzyhOeJty+/sAWn
6Y4nrHL5hvh2MGPXMA1i3UOFR+MmZeixAUerFg7O9QSiHFC7E15OxeWxJhg0Kssd
mb9fyr5RUlxlAf3qm6NowN1vX0BEP6rV2j15oS2cGOsmWi6wJY7nZD4aL4N6aXrp
5ZylOCt3wSWwgcB9kygmmf8hDaDvT0XqjIofwCf0IIe/+RrOc14fuPChiHW+waVO
EXu8MzFT77/N/dsbAG9GR7gLPZmkLSBEBph2iYG9drcCseU9oMKQu6gE9rZBkVBA
S+YQS4mAKGNv0vagSuWienHwP3IdxmpbkB9OtiUM8MLX37tKXEEgOKMyniSbbGwn
E35TvLvNDj7AeaBgpZ9tyyyIdOj8rT4U7afpg5kCOu+ELOXnsCDFJP2Gop3XVQl9
XJ/zLI1HrebXlpIbWSLnSfeHMNT+CdbmynD1ZQKObl7RssY2jkSbGmfGtM/oJrNQ
DJr3Pky5wn/Ard2C1inKzYES9CKc2URuQdVledEeOBuvbHS/ALRs5k0t1cLOlgDI
d1QDCasT8H/Wo85ZyRtEpXvDqE292/EW0KHYhTE+NzYOY3SIFOYOM6qnEcHrgzom
KbzcTttjvL5HKUsGqicOlwHh/88w4bp3tTXcxYzHruFGkCnKf7S6o4gV59i0IZ9X
8zwn7dkCZ0wtfqWiE8OHMZvRab8mYBQF411w0d3G2keSJh9EmGt9cBjHfmFBFC7U
UlB/8QfJ/1TJeHSHLIeDnXne3PzyuVi7cgLIB3sGAZ6Q1IyIu2joCiu9L7LNRRgn
GT0DfcsGvpP610teteXqoV52dXDe0+PtKvL9839dh/SzW9B0a7UCDY+thYk9GJot
gQMrMm0FeaV6su7XRjwdhJK+S+Nng8Ao1P/CtV9a+ODk1aNvY+6/R7vWbQoVAq4K
jrNZS/ESxZ9GIxeVoP9ff6osmVhJuK23NEjgqdkWZWHDAT+yx/2mUpWKg/r23V7u
ikeu0WH0guzjI8a8pNGQ/thZkYcDqA/wF9d6B+EI/UD1SLskOJ8nKdXeo/yx+Sw/
gLAqgPzptdkPR5YI5xbZxM2ryOKFajCa10EVVB1b+BQc3qq9OBfyF5sPZKnI0us/
zU9d5o3avcCCVoSy/OGnqWpITmCcM4Nr2bL5oRJoCX5XlU0Tda0ki/+aAaJv/20e
gAOYyu3w6EjQJqST8TYipQ4CuVgc2fpsjlWVAMxXmph3pxCQIhdloUoHbjG+1NmA
5yaZnxnUJ/7gBvGQ2ZszmcbZtJoGcMI3DswS+Wyd3x6MYI4NVdeNZNSKOOkuDNWP
kY50zJYi7XkZmoTQvhZY6vDfOftcod7CteT3VlO/iEfvG/OAAXzaPsWiMmB6Q6NQ
YcWxmCGwMTxJe+J2YovEq6F7cqb2T6218MTHszHt9ok5SnIX2DZp6EsYAkIlNrEU
05+AYCSoV3m1WPbuG0jMo7wvkahUvhf/H0QGYg0o12cSIhuX04xN2bUgzne4QYbj
b0f6DzG6geYoKbYlQ69P3pLIdIcm3X4wo7pCtGuBe+JyW2xWFtvThAn6k26bt+gS
XSXpPZx+4S1oDi0+2Zh/c941WNrTaAz/epO+hhN0kYRL8j0XiQNby5JDnvjh4KqC
2uZNXAD9QwlcI0cXSU52PWVqXoOxR3Un5un7J6MwJrcbDJx3Pbb/lXboSXoQc8u1
BMy+ReUxWZRSG2goUIoSUG77ig0XyGDnmUbUFq2jojzlNDKFWBEzfmv139l7fNeB
/iycrBzkXXltBEOTQZHOkijVeaZbrghVE1qQhn2kYwgmQtJ5qyaJlx52ycZXkF5M
mMGz5QTl6k9lxfmm+QRNxluIbsqGgjXTcdV4LNxHB+uEhq4SapTQ35kJ03jZfhGk
DVzXkb2X1KZBhKo8hRAI4rXx4MPJ4LWjyDkvnVu2AYidVdXDxTHWMWgeG835e3e/
39l/AVNyfx+rZSKP+eQuv5xj/zvkmDxjiy1CEZpXejc3W+Ymyifc67uIlp0Nlm6S
/WPPBGvMp0fGMZPMXcqOHAnNOKQhF90TZmMas/uvPVAU3JKdiRntTPIj/h0IkOab
581lITjM72drviERZE5y07guHq+XX+ISwp0TAfi8Xb5klHXJr8PxZNIgk02mLlzY
PZnO0HdspyQEiOwkUpwMhIUBIQvZxn4qYnFqpbwJL03nCpGW4Khhx733eWPZKzkF
E1Q/EyaVZUplCz37ithAHlEQUCrHcg0HiJ8H/gn1OlwxY+hGBjk5tZCJsfm4EiCk
QOMG5AaZUtk+V8/4jEFqUDrHCH4HkiIA5PWP2esZ5QleIq5URmgmsPlP8K0jAAkm
3geh2H8dtgTDq0aI3JWuoHPaOWFFI30uAVOguUOiImexmlv6WLd5jstIlJIVmXdA
nj79GdXTF/aUpIJEbCtvsCpe07J6xdjgsogKVNWxZPnn5GwJ3UADOZDzi2dp/xy8
XRqfdLFVVvcaUQFR+6cnHSnCNAt+34WFQmCNRzaKDRhQlggw+fjk9V2QUD5f/re/
IPLOTwwM2j62Cn2/DUVNtaXCLTNRxKll+XRsaO0tv0Urs/vNRyyRTa4KZ7O7tcmD
d89/WXBjvhzAHrQCztXeX0AtPX1itDqFo2ldGOwr7FAaljvk1Wx9H87b6c/rHv9m
Ale2kTzdhaxrnJYM54UicABdYdgoqi6NUFtGKLazm9XUGJZXhCPi+dBog6tSdg0S
4GRULXZaBGqSflLt5+QqgUEn8OaE/XwFt7q7DFSSCf/ue6mWDE6Ls9WrYyfH37yl
KCp+ujzs74qP9Jos9+24x8jLvfG3/IV2SBypj6EdSuwJ6iGMZJl3GPDm32QZre/j
Be6p5vHa1mdv9Xktq74ZpS836OLtT4RfI86wziZHBxbKcb0l9q6Ffyb8vCa5WHDN
XTV4r0dn3EBd1B+4cEyF0F4kep6QVYv89VTT05rmWuZjPpNZH1QDYupkm9IIHm78
OueiyIabFfE1dma/jQIxae/u2jlOEaxW2VfwYdGKNaAEn/olGxuZdaoHPj6HY5Rk
6TZOu5MZ5nVU1/i1wZCObuvWF/0rU+krFZncgWZuP6SYRxlunMvzA4vbFmY9Udxs
TFcRu1hhyA0qqjilEqh3cGp8x4KAowufQO3g/52KdBfU4vzLalVQopBneTW0sjCM
0pMEmCcVS0llKX823Z/nWkTOTm+BGZblcD5qGsPu1tPSs+JS62BPvHKXWCM+ciTg
7ffcqwDVL+yY6sWJFsiFx9mMBO4Rw6ORP7XzZ3cevtVQCc6SRlCTeKpH0LrpBvqU
N8jNaN4PH54QgP29F62coZSngpTErBIbml7BVWdSFFYg5jIho4Ko+NCHw9RGFXHe
5K+HdEUgJ5CIhJgTo9jg8+1mf9pSAnUO+7kwylEh9I7h3sX61cXySegCcagtxxZY
EcDQ9CRy6bgeU2bDiOVMHqRitd+63UEgBAJg4IqfeAgLKU14Po3pFOOyVGB3uLse
C6sfjwFqeVwQgozFVB2b8r6APXNLVydWNqNBWI8uInSZCnYnuPH2gRqKoK3nFZmB
7Xw+HJJtr9dxM/iXuf/zDKXn8c0K83q/w9pOAwpo/uOxbMasuLXKvk2yoE9XrQHE
t2bEz1GZozz+DET//RFGLpJh/qapxHrQ1KdVCEqYmRmMvbfoILZfI+jifuCZBxW1
HtjjqlQZhpxmODlEv3o2uQzHSzPGI87rKTJu0VJSMPndROc2pU6EdTC+ugaFYKMb
UwWYQ2ZSf+JWnz6uhLR+BuAarjf10nolhkJUSq4sj8sZNZBaRZlKzls02zT7HbPn
g1TU+JdL+w/tfB28dSVMjys9vYENuOgIIvwy2W+yq0CrojKS0n6AdMDQpJci01q9
xI9Um/RcRFxTYSULWcqXogfgxVfbmb0RKPOq3pFIL3A+9fFUIYVsUA/qbtZyFxGp
PUJuqbOiPFBwOB5gtxiJxU0Wq3KWKqvhKQoKQYA2e+2wukdr+VeN72Ctx1Oki2tJ
UtG+fjqXsvG8wvjgxPM/TNXtiNyQAPDix4GUntV/FTkSnIRT/a/v2rFmMzV+GnQq
lMZaFlL/EesWS3QJimteE0/R4lmU3lqBwGqhh0T3UShkH8XpUYKrGy7yh4IxcVcg
d0XEesbkEJSaf2/e5OzbelV7Q8+hkMR2WAbjmwtDSbFA6rHSNsALT19xChNBtLik
xtnL7KzBMFLYyWiWEZe8e8E6DGnbj0+hrx4klYe1OYbDytX246cfPiNyk+0yLPA+
uEh7eFhrVFo34DGwtbNwas9M0MAEHqFp37MFCrBA8v178G+YLizugRu5DETa9k+d
Ilxzd17j+8222YiP5rtNwVr0Pnopj6fqMRxjYrDdqW/JD5S7Gt8iGYRsQPZX8HmE
Amqn3DYfWWCet0yE7bt4Iqm62T7GrtuRPMypGIWDpKGmR/eJURnObey3SaO7K1wm
qLRVaKLRlFXSgy6lDu/mrS0NpthZbRkhxSCWqkX6J7r7nYa0CJplkfuO0klMtmLQ
nKafif1hXUGAcTJ3VEAL17ZWyKcM/DL/hUzc0edISQaaya5gv2bM2dWPefsorOTB
+NPxj0Pq5ZmhiS4i2P6CcoGAlcc8IosfSHMo5REc/eu+CKebgMaSunA7ob+ItY66
cb1eHNYMikgBiCFR8HfGK8TbD9MIGhCdrq3hac2WfFP8KAOYvApQVVelxR3BzGWK
ubOCv6WUFMBbYnMHZ1EU35YZoctxEXhPbvh9z88km1W0AUSZc27ZwvjNfin2/R/q
TJ+9bKC7u7gvO3QFyaidpB3utvL7Fitoc3Dt6u79jgQhZHTK/oNaQSz3M6ANH4H8
sPkhMt0pZwyjKEQrmEL8ZLPL2SKM52JqvG90OZKijm6R2oKM+rw1vT+zJkRLhpcB
ztFQXeHjDza5sGScrh7OP40j8rMwkSD75ARb/KpabEZncn+DEGBPrp2rQG8I4y7L
Gmg3HtsQ3gaAcB9TRpvSEUe6zzeQ9EA4crJj9Q2qbD9hYe2xtO/DC3SM1zSMi55c
Gn/bNlev3FPWQ5Q+CqPIq+ZmpNU3KjxX8D5E4RRanBq7AWj9KWbT9kKOq9gZU6n2
WqVVx9U3Ot+HJwlhrbNtrBC/rBh9F/7O53kMmoLWYIqpPUEExlC5jJCV4x2BOWdq
fqrXYaaCjIJ8f+XIJl4meNWFeUQE7GLJeHCttwlnx3FHMVHLDCdPaLrRgvm//5K0
LFoi+kSA+KoFAg7PdTRO4QPNnCbD1WsJYKRvWf3dIsb82Z5cl32OVvolSefZhiRE
AHGiQ8ieElmmdBvX1axHb0XSU7aUPASi49wfcqNQ9h1Xg/7M1vh3tjoE0twFAgTW
J4pe7zidjtsafVTTQx5xPEUy6kybIjnr5SZ9uQOqY4ySa8JWj6zzOE6I42swGNbh
m7W5bNfbRBQvRm9Yw8A/AX+mdnrgn4JNUhDQuH1tPuSrSwfYWVgK6rscKLpo1cZE
YZVyedxAJamFy6GgSiD0qaXiBOVhuRjlPzCj/jbGHpOBYufLOyAxB2QjkhqwjzYU
M4YH8W3L1dyfOkZ27bvqcIzT1NeVBkPlMUSFbW/1bPWnvlQR6gl6QRt8DPrqgwzK
4x263RDtQT2htSmnrkFai+jwb59duTqHcxIto6dFEVIQqoLrODgec3CndJ/PWzPZ
oGGVFIjCODQgA98MYaZ1gEAFjNR9YkT+b6uI/uZFj1LL5F2Q60vxOt8/qGb7bhC7
W76Tnjdrra5q3M6yhi1JGxkPqL+eMeHMox2jkt2cM/lKTkytV8Pwl5Athl+166f+
OcwKRi++5sgJeIz7MFZZHGvu3jE1ZeCRxVgpt24spMiafnwmYDFVlGEyBmuvRNxS
8yo2lTbIG41UAtDHzWgg9CPmoTrh5t20PI0/IgNYjCgdhQkBStFeVcy9PXP7rmpR
zhXLuUyGLgLRsVfeIuGSryQYyZ29x8q4QLzoFdsHH+9N0Bzmo/hgN0AzUSbsXlIG
DRduiZjLoyXszoWYHy6YHIR2BDhxI9HgY+dczzfi4lQUFdatVH7EeKOEk5ussV9q
jmWcAc7odUrZ60OR2U+FzkmPhLKpFQGWCXUwhoCdflinUncn5ITd1dulp9dlhZTw
Y0BJzAmAcWd1FK06Q2MRhYW0YYoiKQjVOFvZYFb94TVzz9oHQb8FAdS2UnzUxTPb
GPfIBd8AYuZy5KLeIVo5DyWnLgRDZguVgMR47FAjc52bedXJtbeXAoB/kP1Mxj7b
9hxUDGPctL1cQGd1Ui81RZ6CiueHN4Q5KN4HyFbFbpibEyrOSlZcXc4sShCjIEWx
26Qvz+Zav+sWsyF0mlbUYWMcZRlF84agEEzIgmmwl/HDZq+AZ3fUuA4MWW5YYjwX
U8uRmbDOF2fM2+DA+11arq4nnAtzE+47ssI1mCYoMR+b7EwS2/k5Vx8bR699D5Qz
3wPTi0zk7I/l2r7/J/uOm9YdTIy+gRFAuUW7sdOLNOEmrA9kUsWaLCungE2KZCI9
qkIZdLQ6ag1jf80a2Bmr9HWKZuSiIJTbwiNQkLpGtb7v92vomZ91bs6gxV2uvW29
kKlZPxtQDOHU9f3y6FfBhzsnJmO3GefK5NlAgoP8yuIgvcCoYrTUezcbVWnHUJ32
rpEog22bwHa4QUnkTu8dKtgWmpojel6Apc0W21t/kDg17h+GL5Ni8KZm/LU1Oc+C
ENNHqHW0u98h6BPwhaRugx54uC81JF8w5dVCLB9BrKpyLOY8Gj4lf5+GBtgx/soM
mqS0kljLLwxO/CEKv8cWZT8D9Jo0jO7gf6bmfWLVTQHfY6THsEBLgAlNyJLerk8N
GeXbgSYgdrLasGwB5FBRXSv/zQQBxGUo8CDZGeVIMEywj1+K13Hf7WHOLhisTa2y
vmiNA3ax4Toq0PWA6tU6ZQHTnB/SkTsJhtM7/ynLH+PvAGYUaam/4fO8FseZOyB4
cipFR8j1Ng1rFQBR917UR+xrcDdns88MeHTFpYyCezqEo+aRKsAe3Vx2eO+gYhc9
EEHX4S29ijNig+fuQJtcZQOBAQAj+PZbtck4w0v3kLWXRt0LIW519/3NR6BglJGM
oahgwcK6+3/UH+2MaedoZBlCzkQetV9fvr1NOGHuohybZFQbNpDcuukVclpAs4Jw
T/JUQ1YaBXKP2x6Pp0eR3MsnZoMwn9iO/wzw/xCWQTip++IyXyuQXljMqEG1sy4q
nscwa6zYvQZmjRsa2syiBvAGxfJbZLbtItmQpsusnEjoVOjeOM7rj8bKDFiPODh6
QUJYbYBnG/BGB2n9ROgtMxhKvtFXGZBaPtpUttnyrTx/dBIxOi5lqaoatZm1q56b
t8bSCLySQMrCX4CbNS6qpaEX4kqwL1LCeqbAnTLaS/qBRMTrvrBqnOWKQlt1Yu3J
sD7tvd4XtSPP94VB1kbR7jUD+N1sS29TZFAsi7SXA/KfPSVD/eEdATk7Q5OZltht
6f2dJpo/3o94iTAjz52wQCvXzK7oqKhOY+iNcr2cV1+TwilHTdEsMTjOPHi8SKfG
2nW4auhWY7IE1t1S/DMSq/kIcr0LkO16KArH7cO7D2tUOaUXQ0gCyq8Y3Pb3Mqfz
ser+4xUNo9+1n8HUMdMYpG/2FOZk63LOI7UMPNj6w8tM9jP0i6N+LKatBneLW2pg
N9tBLbFpTAkk3Lp7GS8nd+snA4Tj2LANoB+CLg+6zY94WZaSAqhx7voH51p2VoGy
FE9sNWHqGwSqfbqOJcbL9KpSBIbee3aH8H5Mr6Cqd5v2gEiUrpmS6Ox6NjDri/qu
5sdvA3nu6KxZ+stxyQMD80P38JN4TgcmZCzgzDtUQXNQcm4XcvnP/YhjGmiz6OTH
pYa/UlMONxHW8GcC0BqadPH4W9CnUJWtogP3syGRMDOtWVXyQ4knf9am1aq98JNg
hClD1x7QPOP7fPyDu6XgbmrOHeHvFbXKucqLuBfl7uw/9UqoECbSceUfBz4XdlzY
o6Am2f00Do6ZMSjj2AVY9wz6Lg2/xNuhJaE8hvdX299qiD5lyhKs1432q2nDAroi
XppvR3qWU/MZFQt80MfcPv/zpRwA7PB2kE9tipGNrpH3k91vAXp5LyZSMMlK0lSp
DCz45GbGoZOBbP3i8QaLyWKDVus359RT5MGHUZMQ5bo8BtPkAn263MNMfkxtmWLJ
hkfBDKCnKb2p5gHmwfK4eBPPcpzcBWs9TPIPschN0KxSA8UnflrX81xcbXp8SADa
Rksatrjh1O1mpDmjspPQkv7hp5rKk7EKGr33D5+pJBtnhEY8e3+5gULbQJdhnnJq
KSpMbf1mDRkPBvMV3hCKA2jswDcd3PFlxLTLd1hqH12q56GENrbcalu2jIZAG8FM
wZqZbM6ibX68WydIh6YVl/gL5Nl+ghDTG/WJGrxNTWn0AZa5pcjnlvCy3sc1NyKl
tjtS7qQBWZnYJAchHtVPL01VAwz3qOJ1md23j29wWsP2YrJKf3n3Ld1sKj/1lxz1
7xzMlrO5lZfvi7tmhRafTOsqwdw2g/+Ihlep0Yfc48attZ3r3hSfmqOzNBGnSVDY
9AlcgmuPuT7M0KP9EnhxXB7lwDZzssx+lDO9LARINkuNAIbnC5+qLshwF2lvzLiP
fgUFrkHPwNVRf+2fD9eDqm0yEvKfhvLrrrEluEPkrUuxnEsp06SBNRmzMJls98aU
jfpqS1RGwcQQ1Qkss/rYSJWIVfZcetzmIn5Q2fIjCNlto1z5Y9S4i4mqGoyc4bxd
aO0s9lbhGQgp6INn/Dq8FksmISOiUqnkjL8kjZdwpiWZEdQfigwmoc2w3s0o6BAv
i7mrrmTI3huBhajrd9To29ghpsfLyCuL/eoTJFIMlY1apdrr5Zt+zZWU2YVfr6l/
SVQOB1624B4ox0DcNppBtp3DdF3v2IxSsXQcGPEFk1zqMVXy5t4c7hs2DARJlVbf
TGVnZgGVtKa5GwgUX02JDBSXWlZNOBylOVRJwJ+IXln7vIEBujGaTRrRVxhqr9BF
9Dpzdvm+AyDnACxTgT+0mivRtPixhr/p2yvwwJQy72xa0Z8+kSPjF0BpruB8xTB6
moD0rpq8tlxk8Gch1yDUTmYCpZzsTxqZF/XGUTtIlRfxz9Cx3+4edzpfm4LjGmLI
v5dTSTzJDNpf18r/DXslW0pZzp9kMrsSeCyAW2Dlsul2M/9dyCO0Gv64OD2BKaXz
lhZ20jzRyw0gBzOeKurw0YClWOdszfdlsJyg0MVHZE6Rjp4QNp4/umKZXb5cu2Z8
oE3ZXj4O2AvnuL89LB15U+82LioqVEbAgtOl7AWOQaEdu6pTwIkAj6tQfwRP+En4
jkpra061l5pC74z0M16ouWiJ/2Ug/NTgGDCoRQAm9sXD/n+HN7J7GqgvvzeDT9XP
3IyxD+fe3aAdN9hzCdv/PDOen5sk7lFD0xq0dLYtDgMyYIQVfqVLbveP16U/u1n9
14SldHo3xShLR9e5VmtceraMb2fi3sh5BUaGEERhufyD2lFBHp3vevXKkItRbGHW
bEU7lU6q5pvyc6Gbod4KcsdQlhov8Oeg2L6eTcLdd7YQLc5chhVkV3Y3ZmVbnWec
HsyTaNf3zh8dClFRZO9BbOfSi7qHzKUqnTPCc5dMkexZkCG8lVOWBcech/7kqSOz
X1Jtjhcf9xqNBlGB07YTT4aofQVN4JrqOvnxT3CEWwsbsas7v3+T1Sh+QdAwFoJ8
qB5rC/eV6F/ba4HttkRjbG0HSjW0ThawOezntEnGnr3n3RBzNRZyVEGxEhUvB8DJ
SWhNk4MOin+ovgh/4jZmm0lc05ucpgtw8dbAkRU7gwzL+q9BAddrKquFWiKT+Zsc
hsYgfXYYEqPTgh86YNTyB+/nij/QgFuo92dIcII/DoHYJ1OzLrOtsf3n0leZbXZd
mG3Z3A6O9M3K0Id3ECWkj8A21qis5w8A18z11Ks1YAUnT9FixSs4vjGXLuoH5A0n
13Bs6KZfQ5XG874CklcJa34AII1tnAUX7eXdr9PWulWC1Cvm7xdDJy7drsyU1uB2
6/wS9S6Uo6kDl25kzmenoT1lN480b8+ldRYwVI+79CFuByjOkbCYEmToBw1afp7s
tSjgeS4y4whWKjszICOZGdzBbWkxsIncU4/k0XbvydegFQAbNObAHw1D6tBvRqoh
HV/s+ijZYGrchzi/B0wXOmMryrBCyc4YDA3D+qrJ5qJsOKiCDiceEimMCzsE8nnZ
8MCyOw1q4TPC0rlIPKaNAWdJIc3bVkLyWASdGw7Il/EBTRS6oIHd9nyQCKcJG7mm
bMfVSyaJdXPfPRXRAK7kMevgb8stLvljcto2eGqdQ/JXJ3cRKGdV2sQdcY2iRJ9W
Xm1zIld6OeA409nwGfPvKIdPs7oAjke/h788aPoeCy1eCiQB+RAzYnBGIBNKV+W3
BOylK3UoRS/ixpG+lvWz7MNYA+tRtrIBLsJG8OP44vbJaYzvwzg0ZBXfaK/CqkuI
T0ArbPxLLEeZxYflek8cm4542ON7QqnK9k7YCxf93FGgyKAt68M1+2HbUG7+Z3jv
0R19hS0edw5dTRC6in2soIhwOZF2+ncNJ8HBXs4aN3PzK4VxMemEIbXqeniESVvo
0T7iD4fvvNqiKyAEtUADNZlrOaKY8bEOZ+ffNQCogAUCAuC7XK0vBxnMKOg/QEoz
q/0cLzcjMu6IH7j1qbsarKhMlqbjP3pIM5NeJGDqIQmlXV3bFgxMgYZ+X8iihpQI
PzHA6WKMvagp7lFYizUu64c01FdGjefIf2gZpx5gl9J/U3E9wShEeJfj99qN/L38
lpMB17sHx9injqQx91c4C/xJP18qs9xstmIC3ryYoTFpFD2Rpmy+Z531gNLwWYyt
D/Rywbn5kThKJ4O/AWIGF6pqoBYvUzSWMO3zdBFphwDjpZIN1a1qH9fvJOmYPXkj
vijxw4UjPFVftAIJZNMwmdNxXBYFqY/3+K6m3HOMcEip6XvbqeCjGn/EI2ogq1bT
opgGugvejlV4jLatW3q+7Lihq6we5Ft3aL0mDEB7OqgNO8BY4kdrYWKbZUGmAGdr
px2uaSfWsD7OohojTiRG5nKqCAhIpAlcdcGvNYOynLXL905SmzAOSrCAvP2CvYJb
jrv1FlbiGv1BvIR1/SSCBkcuNafNZNr8kMtSz48c4Gl1iVWK2zxEoUZJ23kUH452
o7zv+B5ndj1H5x/tOQeT1d39RYMfOgKuZ/yMkfCR6Frn1f2v1JzfPM2gONm9chRz
gjlO2A1RcRZz7J9aMfZdpUZvHJHusuXLzI31SLYzMDW+9LAIheNhGz2Ki36uerqf
7ey2D0Dce5nt2b5iKZ2lwK4X8iscJIxiDKQfclVO8v8nEqqo0lWyekyE63MPUfi2
HYdcM3eJpSqQhV0lbSJy7tx9UOKD6XY+FnkNcaslqh5THLr1XA1e/pyv7X/ZiP5W
8Y/KeBjlAwbtDt+DuGyGk5lD57wOYjhJTWXPI65IgSyB9aDgrb6XnnGBTjPhgIKd
uPpGYw5/cdZTYj48NVPTns/qrynGr/A6VsIKanSSxcnm1F5m6SrZHoDJi/ES+ZgP
0QTSaJ9bTf3vrkBr5NZX7jiN0YODfCUYWYTZNagonWrKp69sBlNzkxZGuegtp4ku
nL67VPEFuYbVBsR830j7/C+e4DdcqLfiWppTGuIYjtTb7cM1yqzKeQgm7jufW01g
9DLt+athQkAv1q/n7YcEAE+GrynngNoLpO/Hh9yEkXmHz+p4OWTqb0bKXBo0go5p
1iYdmYsirVu+wY4fRfTyEy+r+Kae3Y0iVH1q9BX/hxi3GWQWoz9jwyBK0PsJmx8L
+Q/uOYJbkjM578q+zXZWvJVvO4/5ngQywOZOMiW/PGAzVHv+qkXU7ykQ801bUpz4
ztX7fk6Dxz+JxJc0/XqZBaJ0kpSZAqdc3kr3dONc+vJcnjvac/vF99I5r+N9Brqb
f10VPJ4mAa9NnOBTRL54pGGXNdJHiFa4ats/MuhnVQhh8l/oGXPve2eP258YkLsV
JMwenHXxj0H7+4XZWdZYKA4lW7mKW719Pd0XGEsjh1j3HTosucDKSE+0EA01m6hR
34g7dDDHd+rYy0l6Zdk5y2N+5ZWvG/ThA8TU0ylKMUyNNyNrgobbhee2+SO17nTy
UupZ9dxjS692as5Eex6C2ZMU5+N3rv2lgL3pH+WCImdotqNcgMGxLSEfcZDngKst
zCfD1rzZlt5aZvkT+ZHpNqpbPyanWI3YvcTxAg0DXLQHMPHcyyfLHpbPl/XXn+UG
OuqlOjDmSm7VjMHNLouatyE+wfEY5Vd/jAREFPMzoR0VpORQOrWX2H1x6oDm95HF
wXFflUEZL4vL5RmojKSsoGFg9g/Dhk9b3MvH23JKNhEL9JvnlEUZB9+6U7r/IcmN
Cus894L36SnQhhQ6mEnuByJKCqJDs2C66L+4gwzb1zT8D6GojvYQFpawaN0hsjw9
nQRUFkh9eGKpWPYCNpCJ60Aqu6V7YLRrOOVS9aNmZ3sYVXBjs6Vk2ko6pL4rImnx
lnGvsEqGQK/bipLhAbKofiw8V8lXpvrFnD1XyhgIynbhuFo752jNql4cBAKV8ES/
N24au/Z0sfM4jHVoT1JajpupY32Pio4L6UrKnoYcPQIL+yJhme8JhX3bdeSQ87Jx
Db5nwT90mVJDeTiQkQhjLF5ePCMP6C7jKJnCAqHi9yy9RpIqETA/ezHn6rI4zXco
wcT2rSx2yc1K5Xl+n4yVTwO7WuimsbdFHICNPGb3nU95NRjFVU4iNMNbQHru8x0Q
/iF/0f0pTmUtAU593yDcnWLuOonp5BEULmKBNXixDizo3oMsNM4l2cTSI9EUNoD/
YeCsm2k0vrXtQVQQKGj3QDDIvwji1JayiW//TZM0mmZ/DzmaNwl+s/khQhnuBfdr
av5E/SbGH3DrAZXF91obpXP1WsGmnDS3OjJGu3qxnyqwEg6XgS9o/xYmDJUWkXN/
fAH2fwN7RmiR8+R6BLi1XEEfCOStXAvgC/5BJZPGGaH7QiSNL833K0jCBvl5lJwP
HyUcdbpi13/nJEmipeq/WQ1x4VJT/jsegEVKqYs8TPV8nhBipbh6vw1C2LijC26b
XxgT8qPrFI67XyNgyhf0/+ZanE0diVjCIfoFILWbszLCfZZ/DzGbAipM0/hoqQan
zPQW2bvZLNapcuqnAQnF69A1rcgyuZcQFAzcXDojlvRMkI7CmMDZ7mLKE4x84I30
N7KMI9zps2CUGVtIYupU8TS1aQmSe2XyvMHgapz4SIfzn/HRfHvQ/vKVj+kA0LCr
SsVzTlYPMdROKiX1h825QU1QWa7tazP+lBO1goXFGI/wVCpnXLFtmlJ5n7iS6ZXr
vuRL5yZwBeVlxDVUv6TLhi6+HnrzQSuNwgh7EZdhUseDmqyVEut/gDU2ifD5dmvp
tijglKzwJ7Gj+EZIiJVHjL24AceLNOJFUu2pTdWuA9pZhrAa5QzOzLR3Xm/DKXQu
JiuOjbATmotQ4iShuhbNQeRdZKSSCp61shFrINwuDQA4GASI/3SmjxV2wlnQIJ2h
+o9IaIp1Y09no8ge82ZO/MOqd3ox2APNe7wAOIUA8S72K5Xz54+5oFBurStet3dv
DFTg+cnsMh5Kw3BdNq03csfqJMob+spu7Og2jieFHBrrMzkfoopb6S+Aaec3Gvfz
bWKP8pPaRgcN8v/cTMKwtzFKK7JHCLl6jzyaN2N7oob66dGOmuGMyele8S+7EwBw
DcdEd0Q8UWmbXj4bvpco0+coI8U5KMGNtpWq80dhrO49pvmSPWW00CHRwZdoOAXx
gyLRHEFFUMU//1ZyqWsZJFjGVjGajIX4WiaH6Y2lKLig3MCzKIQeu65AIWVWYRYc
H409e8TTK+o/xss4SJwjPiOZTO4pTcYR/CRtacNHsSPjhNovHU77Gol0m0gINDEL
EexZBF509OFo18dFtdK5T4CZIGpg3vVKIlYp+1yycJ7CjBSpviu6/z39Iq/5WJRs
TE+yMbyOxqLEQLZuUMeWsc9wj12QjcShbAqbcXYPkVV7rfZ2GFKqubjKzbKLCZaD
TERvGi4ZwRBKRHzjEBW07fYdsYN1ubHwfa7B9/cAUOhnrZtwjkSD/8eqeq7px/9n
CiJSV8S7AJar9cLr2S2A4s8CX9h+YPrtmeRgNrRlFoLFZUJLv3KnYxqhKacrl6L9
lfB5rigMtzLre30c/L3YYo7BfyvaDSlDsfdZR0HrAYOPE9SuYvoGuU8rPoqu1v/I
FRMbfuDpTPbFZ1smaA3OdUR33VaIj+LZOnB56Z3OMc/9/e08NKimetjnncH+WEyt
Th0I0FgcNA2myFNKZEvY2qcw5jinut3NAQNk0XcDB0gYVswHxF22ve1Lh/Sl5mnl
qvVXBXOeqvp1RbdNNmB4VVeDxr6wvMoBLSUcKO+woUTzrQ+tFlTSBaTPcGJqJegx
TCLjmM2dzdEMmLQ2HiYFe/q/i3jfocjd8lUyAimZceqMBx160Ou41rVjBVbD+PSq
8NNqz8mZfRwwJ628Qeip0OKrjuTJmRAG+kHyX5tg0iaDCvbKIS5D1cs3ls/YPzXu
Hl4CiTNgm4N7tLc2G3QKBFVHS9+V2sBovBnEFIHzCykHRkklcGC+f4+Tied21OVP
k1wBuuwSQR1BakhBsM7ycF+d0YVtt1kqw9ro02IS7Vo3b7uuOGE+Xx7xQTpmUc46
vEHk6whK4VKix3F/OfaF4RzvKIA+g6Fa8yLGyhyTn0snkJqmT02xOBlnl1eLwnfm
FnHrWsTGln8czWECYJkmDtxFodc5S/j/VvfErqK2swECoiHETrDlIUt9+jJ4pzAy
Y79K7OpqPDm03Z1z+jlsgOpAqwpisHH9QqxKbf7jj5gnM0/UPQDeR4lKEV9sZghA
325aU8i8+1XRb0hwYh8S6OsMG3IEtU/GCzg6pTFGfEHEvx1Z+yTypaHUSULBOpWh
8Cqgb2Jm7j7RFaXh5V2TTjeYmO9AULIi/VBmWkklR6YFlMi9VzsTNbssqEaAHGEP
s0sMBLuVOV6V1bfur4036x+NJIXskJ/9K1fQ9dCjNg39bYcnxM4E2jHe9HtsXqNg
MVLxKSrurJxbBFbQ6GFKk+RqtQbnLrhw+DMp7GMJbOOSEkr/FMmbo/jWWT3e5T6x
ogJwI8m2VA7piRWn8OV+pZLmHvgj3fqnaI2XIFtOQ7DeylBggiT6w2CVZeIv68Kz
N7VfHnsSPK6BdsUfMSDxTpzlU1Rc2+Vpl/Sn8yGKUEGPGSkmA5CXt0Wdql/en4V1
yAL4lI2paK6GJPUuWi3mMrVFNRxIDYEgMURju07uDuHXC8by+5OZkmqXdcUT4+5R
Jc6yzPwStWzjGpA4WZJFTXwa4xRMnsGePNDLAu76i3PDdfHd1kNLRasRDUg8ok6r
+ph77CTKozB6n1wbXz5D4WiRZA/GjkGL7IXEuXj0iv5sBoYZ3iqCOsfS2wZlWVny
e/MMcpK/9p/mncZQr46Ynpr4mwG7/5X/SI4osBo547RulmHePw5fBL6GdOJJ6tk4
aVq9duPK+nUna4EzG4cMlL1S5hWOQ4gOTdIEuRe8sMTaLfmGE/UxtZ05KIGB8RUO
kWjdyYL2qN799OKztFy/NRjO5Db5WZcAZ27OtGctwROTc2/QsWn8+h85WIrzLEF4
WoghR7Jfg30ytMvzE1RX/vtwWpcUEFwOoqyfpcaxk8ecwsIr1+n0/oHPFONFZhG9
Npo+qGFzKvyU4W2IGeqI0maMb17XifME7ue8WUxxHZjZVEW4DGJwJ61gYAuDb56O
yLua5r8IdLXoINy4NOkR+Jxd3xrqJ+wZJipplPcNmvykeD5e/60HoS1FmekTi99L
d2mhNE40huX5Kl+vVry0hCNuCN7oHZKNvqB+0QlEUP74l7VZtF+yyHmKiPqLJ5ro
MvCmqam1rlCJN8G9E4gM6LuBhK9k0NLRM69wOSLtt+VTrWdGcWOO9ZC5wdH1cf80
82KY6pNut/oPy9/HwJeXGb+54CoHI9y+v8T9WuFdKmUYDWAlbx5U2oUoTGilibjI
PIxUxpkTqB5OAF+ktzgLTFbp+7L56p2Q9OlpXccblLEWpbJIyUlFoxQ/Zfrx4CPq
mUzeXLV6QVTQ34kpzdmfN2162a12sq0J0T+zHthxRbzuj141sCGu6ZCvrnO87F4j
bBa9YXFNboP1pY0EWoD5KQcHqno3YeMZKd2DkJ55rqjL43L6+v9i4iP4sw2fNS6J
81hrCLV+HXI0w//dPY2PjOWPiY/eAtO7kPwTrFcvBNqFbodyh9lhxRpRxbB2Jxjp
XBUUpdA5rNRB8lXDrbPwSucYUr2sFqVhIMgSsHUXj2az8NQ8Q3DqoMDv1caonZYQ
nUQ1LxSldDENVp0qJeBdyxn0LUdlVg0vCLeMI0Nl/+5h1E5wZ1qJesLaakK0+mwc
FlQ7tebv2qDm2CKPsxeGIKuhtlL3yEjyuLt3yWuV0W5LSXGeqhcBYoPZPPGjrYht
t6Z3xvUG2ijrO3yFLlutZAlpngzYf7Nuk30EUbgaynQ29WDe/nuiXC1akVn5YQ6n
NkPjNRDJ0/MOBX2UZiaR0xZqFTrTDSi4EK6Sg2CS5xNzXhh9+Pir8MrjTDFwy2Lq
FL+P8Yv21Y2IBQbGPZgAzkIuasz1djWgaAU4yUnj7xmyZbSpIa/8aE3rX5G3wsN4
69dzwhC5Y2ztrHjKf3+c79a9KVRTK0vb0Gy1hSKbh55r+BINLf0mhuGSGcwyOWTO
c3A0bV9VPEhE1CeBSwOdnlRKX7xFtfgFX1nTPdrmXxAWm5rjoXr3sxYb7HGlIPn7
C7EsI0jOA3miqh0b8jM+4C3M95oS3/nY2UYbjcCCJsF1DyQCU1nvQw8T5hHYeoU+
dLBT4zbAAnBPiPECLaPq56SfxB9fMIU9/bEjYYUrcKWhnf8t8i1POzGp+f69W0uj
xSs/4wVySc08nTdjRsl21vVqxARPp+bXIDtO0Nx7cCaN3/URPVymO+ugQ7MtvHLM
YrWV5t8dUMk1DpKvrRebeGFxQ2fevdB5dTpbaNS6aoUi/57u9l0/gJSfUG8uL+L+
q1s9E+YPo3zI36GaaNuq5sT4bgO9oHmDu33cTiKCmBVI9GendEvU/S/s6ICdn7+G
62JwnWr36T0QYoJ/eHBDifGP3/uYkIz40TUz/tn/UMt3mHM0/7fi50R+oQU9dva9
DmUUCHyefaw5f42As5UmGb5/RIQSYzaRy4Y9vRjsPZTVjgiBLvdJ75nsFhD0vXNO
gf2XGiMJ69lnHicMSuc43gnJyX5WlJcajD77djdoRuBF0JzIAX8+Uid3KXdLV+ba
tHQIPKxkEqJysH9sEjgoPI1mUjo9ygoNVBX9uv24HEoZcQyaZACX4LqxsS/v2Ovx
hbPbIJ8QofWCX5ItdnBu35vPPs4+Rvazy0yqfjqJ8QAj35FoXMAFF5xzE+NjCFn/
lZ09aApanBOLs5qeyEblAdhHNo6HdOCdzmH+23wQUI33PBzVCEhskkrNoOEC83ue
M+FmYJyfCu1ifBNgInYD0bY+wTGhSCOEmujTqOwc5LuIIp2Idr5Hf6Lo7uJsHlo3
65Pu77FYAN3lxYE0VtAKH05wxpEX505VCvj5RSECy2nPKsGsrODjxlY8Nk2QaQwb
sSGh0q+IpDL7hyhxeV6K5x2vB6zsw83O2mODPmvgOvkNdVPdFaAAFFJgZwRJPS8R
TQ9YN5DbyXdHGC+IcF9uaLlluF5fi+70mJl7xhNQRh3VhOlkU6jxsZWiCFLvtUOQ
7bJiRderhjmblVQjmsLOml8wLFJsHxDDV403c1stuRX5lhSyzzyKaEAUemqP0BjC
HYsPa05T+lsvqDTaUD0L9+Ra3lLH8Wb1Z593jGUGRD5fvLCH310FuyAfUTpaFfvd
CU/D9UkgPU0o7QP/ZXaUjEbLVVP7J44lFfPMxYULbrtHY8FwWhk77M0CVNb0+fm4
d9SCLULakAqLwZdcHOa7XfIFI2+AABYY8GVu6OsOkUjfigFaqYtwdidgnLneLbq7
GI+ja7sUzcEM1GqXsF/0UhLNv9THIspzZB7XKiaq0OUgemwQnDkk14R/s1hwIA/R
Jn3HOx9F1VQDd6soI10vV93+VJWso3/WGgVKOSPKVfKDNJixlJGj5y+VEiyTPQ6Z
D5ga9b0xd/tYLl2pUQGUK4kiYfpdfGijzsIjMhtr5dmcDGH37600wQ4vsJ4pB/Cl
qRsYs/h0kuOhtls5F5xnOMlrkBSVYu9PFCwEj3zJ6eFGRiCGKnC+9jXEzm9rmqsu
fRqNCLf80x6NEgUMvnJPj669TezHwj+JfFVfqRVJRqrx2BLPBiuboCFWUaYoC77d
WmORe9UKocYa49S178asbzyC45m8NsVeULVvQB9dFhZOWLThtDkceWmk6ZvspEGp
sZhSIiAkaDM0yPSAqt5ctvwAgkYBphRMmt/AR3ftvrlLWMXCBu5lQkGEzUKJULT8
W7hpttHZzHtw45do6+GeuL1RT1OL4mIZxavKAXQsjN7zY4DjAVCGAGUR0RkwG/B2
piVfQ6uL9uxIUrTcIOmfRVTseUX/WeLYQzEAyzQqqsZT7Eilqawz9QfLbiKWcnfe
goLVy8pgw9FWjD6j83kEq/73NUsjTHgiorxcVvROwPM1CSCcZFKFTov+DqhpvXxP
n3QAerCi3+vlR+XASeLWi9At3wnsseGXBYrsFihikEvg/Qz3ACGu4DhcErmr47nz
2XXqZ1uXZKZ54CDoAu1Xp8huDx9lBqXn/irCYcuTp58pAsBN5XC5eNCL8KVKiRan
OEJ1jBDYcllRBW6thTT/ywmJ//FCyUxDdk4UOTJ4f+SITRq8ua5MYvvYvdH1l4M5
wCVuj3hu+Soz7G401PAR9rWdsIFIaMtQQjyqI1/fR0RcsjA8age1an6OQ5jf8V1B
wL+Bxteg/iN1vxEIB8Hi8Ve0vp2/Gg1hLcB2ihM/l57SxRJJ3RIp327r6Ax3LRES
yIpyeQdqLVyTBbafJxUFsPRuhmKqVUs9NfZKNY4DQb/0egk+IN12Kput/K0gMvfn
1GY1Gqzs6z6qsSiAuoigzEW2yA7PeAAIjsK0kNR3OOvdfYCCiZbG3jD1A6LSYhB5
/UESYGfHwtdiZf9fTEIwA/9CZp+l0nTHJS3btV1EVDWIeOLQFvNGsjewFqD9XCDX
L2wHD4mjrA297xiAbOuH56rtAqFwDVZQS9JI0KTZtpmZMv4e4kUzKfh27SbWMqM+
5V+hgnVFyBzRgke5N81vsZEU6tJs6r9dkY3s6M0LGnz2exGNGV2IP5TC5xY6/rob
wihT+ZCUy8rEZX74NlopfTQMhjtH4qE9yIdg/WJE+4Tw6huULovg8IMogoSwU0ny
9qpFO/bfRfr2DgKj6BzZR07oDNB3yfdA4NExpc05/zhklfIht+89PvKJzPYf33xY
M7TboVFHHsFczkoPVZRtnWCwbk1D8m5db6LCj1cDVDYVtdUzg0H5SQS2Yj1F9RXn
BzzY+rekniOAJrFqAztuOMf4awxrsbMefqHgtd/icw6QL9h6uYp/mmBwnvyke7wt
/Kkng6SERgq7GczkDtbVRm+5KooOMuB3lPJedMuE1wdVqWFprjH9IVfdB8JcJAih
xz8kDmCsgnWss7FfmyY+HLRCF/0fHV678qZw6RTjPjE1PQf4f+D0z5yxsMnAOFCe
E5FMcN4CfIkhyK1XnCY9koaz7ZCYmZMpHhkR9VluFfMUO29WihkIQyCCadIKLWrp
atIFJ48egNk117NMU9NXU361/WLeK5FXWaYZ9TEQ4o0P040TzQDiNbOHUASwYkor
9dzkN6d+GrIaKCBhwXE43N2ZS+OYtXMaDJnL00uysvKwgAPhzlCS3ZkP5UrAinTE
vkxGIuVEhy8XWjX30hifVx/PBPUzsfnF8o1nfd7Zmvf6z7PEZ5hc65sGWUdN17jB
RcANTUgeDfCqI40vXNcCd+hQV+ityTcWYwBc6sKGJbb66u3zOzHBGgwQ78SGhzW2
6PMBjOTx+5R7H5z+JA9yDgkedx2GNdJAztHm52eDncBk/uig/BAEcetqrxmH2f5w
fQq/uloQi+E0k2bHSdDJC1nB5fOYVUYEh/yp1M5ePmT03fs4hcQTO6HSQIAJ3CN2
Aya2LnM4754RIWzMRMi2/6iAFZ9TvNProHaMjrJhgSIYbmB2tEPv+bpbIo8EMkYH
lMmsa2zqNfPzcTf19hTlYtURnGMsL554amkpZSACMsqVeLfa4rYEnKH1ASGlAf1u
YA5tXnnrD16VhvJeFR+QHPeWG+++9BcpNH87jBACS8+FmuDQ08h82sUeOtQrcNdz
HGh4p0SeE5XqnJzLWCq0zYj9pHvNnaOsP4qdfcEHBBZGnYM9iIg/9hbx96B//45H
uldw5Fqioc860cYysUkmd5g2zAVARMfEMvB4B3CXfRjqVs9GYWRYRlYigMis/Wqe
2FTqI9O2nyjN65qo2lBAbYBnAj+0YzV/s2zBq4NQdVUakiNTDl3ePx2PWgHd5GGc
ikmlpItsH3YLBdoTXjMPl79p9zOK+PCOMMOeaM7dC8F4lB+VqUqEne59Fkk/IWj9
/CkoR0B+avrvKDjEpb8IvtrjgOCBa3JXg1z1WLaLIF6gNKQt2eEGpV0Vv2FAURHP
ngv/fOmv5YQuipxAbJdbQ3lEKH3ts3JOH//sQtAL4wflC31ZMAKP4d4/9ASY6U6N
D1X9rDRAeZhcmUBYbQNsrY58ciV3HoTUj0v7DZKh+Z1ZpSG1P3Z0W8kLRbkyAIfS
KuM6f7WIgMTh5f+4IjAGwXwOdpx569RpM9iiHvi/SwNMjjrW6SVhGuWPX88V/47X
oCnqV78cZwzJI8kZ1FgwD/O5OG6Sl7Vswj5UOpNDS85vZmo7ZTlBPXFz13ue58WS
K4NclO5xxUdkill0SafN9VgJ7zyoUE5otMQxQTTEKuk6uWElZQ2klb8ND0qNVmgG
0Zi9OzbDRRrXc5fYd1XyJlujopaWXDhvF3UCMGFZNi0wR6zpe7e4+i23zXX3Oeqm
5zE6cbVm93YUqNvsl2wmDd2cygq8XnVr67eP2q3/pxnBN6oTokgf/WdHX3Gml5kb
DNbYU+AR34CG6EubIsme0uVKyeWB43IEWoJE24MDMqSJWKYtp2u+jhcpOiEwPQBg
cBZzn1RoQhXbjWMb16T6iRDTAcgUDzYsAmuZbgqJ/WI5TFhkIkcCL7NyPR5PRbnK
h7h9WN+DJ64NdagAX7z2nj+5TJjmoQDRE6lKV0nSxnSXpfDiVE8BA7pGYMkdg5o2
wrf+wf+pP9WiPlqkOiomhv1Dzs5t6UsBA4BOxt5SvtEl+5h+KnwQGEx/5AWsYnO6
K1UcRNmdkFcsvln74NiCcR/owD0tuEilRvKE2JPvJ+JHy5/58ALoYIaI3lsJ7Zer
Cp++knKefZ0jK9VtJ8e6kWKOaRWN8RwprUCc7Vdv+2aD7/bsM6tu+ndMC/FlQTt4
b2WkBJTqycWQ70ytHDA/8/YkrxfP4TVEtsEyUaCByiA7IuBkcjDbzhRsJ3Erh6Uv
xpA4fWTEQlo6Kf/lAv+FWA==
`protect END_PROTECTED
