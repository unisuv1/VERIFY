`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
je5ZVrvgCZejKe6pPzZtos/fRDvvHM6EG5Q/0B5WHN4CMnnPVtVky36+I8KS6ePe
8uuuTa8vumgCfdYcZcIvJPDYerA8x7gJlmemrm43hAONuqbaTS7gH7nuU01LM5KQ
ZJX68HtbPJ0zrQT7n1B6XE5AAp3j76KrqlnG0KaCYSTew7qxWpGZrwwgyC4HLuIR
uF8g3u6FamOFn5aZuIRnQ3NA7PWAxmFnDCpUmmcfid9PzhNGgS1bktABPVWd1CXR
xmXnPZwa3kvNAmJ+FcVuGVIt4auqVx/0yHlABq8/qB9p5VsfYNdNLKNCsFA/AtWB
lIxi27OC2OlkFIE6nUJ31icRWKdTrR2vQW0x+W39aEhIzIGBaN3YRDpJulfib2qD
ozqIaRGOgWC7TJ3zRWrGhUUdSMiNtwS1m1gBiTsfY7dal4ZyBV5vUStEvKnJ7Lmz
UQWn5sNFvORhX3euMzJqs7L9aZrb3Bi0OwuvoYHqTFuyxW3yuGLOudT0j5siRk6B
XiPT8VM666ht4NNw+epGRKS0K/vjfNXGfD8h1Iu0kVY5yZDVQ2miEGTA6a/WKz/7
Ss0f1P61AO266I/fKruTi5YqLLYuIYZL6onMS6ZQ4F+7RPTPLBjYsbJQzQkx4d85
82J3MWp3LfGccUcQsxy7YzH12anK1yHRjMTXv08Va7ZBNlBe5dd4TV7jY4ct049M
ONOYzA7wmlA99sH/K4CJCgFC+gKMiQ+qMOjTpVJ52kGrLeV7Fo2OuOCFYrXFxoQw
PD72w9uI6Sgx84jZBH0Z5gmiI5bialb/ZOO2mGjKiMxG22dlWQJnpsZwOzdbiaJ9
`protect END_PROTECTED
