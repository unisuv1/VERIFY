`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
D+mlAfpqWfhgPvQcUwQilfH7EeCFGuzMcbLhr38nd5AE6LDFVGQPk/1jpGWVnOUj
inXfTCpbrhMjNTcuO2z8WE7Y5/6BBFoN9QkTx9pLr9oBrvan3QjK83taKa3sS1F0
us/KWXoqT5EO+GlYjDYoaIkd6nb2KhZApeRjXPvJEulmcKX5kIZI6uGF/+ln4Zbh
osR4uJxs36QsMogWLdL5DxPL+3OJIAWdCkVrfGhBgTlZ3zY8a39X6/nh62yB6ONF
4hko3LkKMRlve9Sv8FYf8LQJSDXJdYtuSwavVr1powdeDxBbkV1Dd7hgepr+SkMH
ZrnvDYjA8Ju8UTefqNMgvTvVD5fgxDQNxdQffLPQ5SG4yZO3y9wGZu9gLUuRell5
RuhQqA9c2mDdJy6og1jytiCMv7nc/1/HvXaedCOp23AK0BxzX5iAg/iaUi+RDH7V
JfqNpByuKx1V8b2kznftqD80vphtULzLWf9kDvtN15R0uLyDZHLwo0s78uM/pAs6
EvqypHoXuQxkGHSKVDnccuWB8L5z0hClmAgvkua7n7pQGqK8IsqKTCOdhMAGYOy6
+zBYzKmPvQ+y9udXmny/ulTtnVhpoCrS4mSeIWg6rEDvd9oQ/C4EsW48BqjIAH5F
/06DZrscrvKLRnuGdvgn5lWvyrsa/0WwkzCyGusB7qnxxCVE2u5CBMoxBAagOUAx
lMrWMTQlZLWFgAmXLAAnuStQHFktdJvjE9ye/b3XPJ7oNgPE+1pzaNtRRpCVMIGv
mew4iIirusUyMT5LRnkw8y2/hN/bBNCRFaLBJKknWLCHqzyuClxQ+uxhnAz+CLcD
W8nopWKLDWvN/NBvbPy5xRVGk5EsKaOcjoD07JvBBuy8AvGPf/5s1YET7FDmGJ44
Rmt5mMbEppQocBf5Pw0Efv61IZtprr6cEmM9h4OPT7kX8hefLmBqfBXTggOu53yK
+AA52xRlWW4puzrK0QUZZb/WZInlfmVlSBljGRA4kPJOk+vjiiMKisoyGc44VCzy
P/2IJPauljz1TI9DakZGQcaq/EeYmFO1ccgHBbACH7OwHPb9isI2BJcUD9qRtPzF
4wFhbBCuHbvCINW+iciQgS5tQBcFhAgOwGyrEMVcpG4Q3f8CmPIXxLZ3nR7+4aGL
4fCex4f8Vl+AXI0F2Tg8V2FnOI5kGrb94AKLOGa60E/r5TU3p4y1jl+WnVPwDusM
ti5b34P+miOyvksfoJ0zUV5yD3Y88jtdBBL6h44W73cM5h8zlug5aGyc/lqhZdD1
bYPvorniWijsytGT9oS1yXQmkSooAUYjhrDAjvyrCnxNW3JnQIeDeEOgIWebrlJZ
SwUwTnibEZKCXfYFiVXEXB6pwExY56tVSneJhnGwimVQhqxdg4dgtEg84qKLiZpS
lelWoFKxzqw4OoFcYhIpfO1Fd7JwF7oAoRsOPH/ANuD/UZMKsEHy2LOzyIF7kbD/
27caeMOV0hRITxQyRN1UyxMDY/mz9rnP49mDhX8ElPstOAygeO8PDw6/oQhjWQHO
KkK5hLr0ccQE4+kY/gumkUJ4QXTzgzymuQxjQsyUtvRT0Nlj8XnRMfULyv1mACtf
sxc5bt2h0o5OTKbCH7s5UV2mhrehU6cLjSWVI7Bsr1Mnhb1FIdEpc47XuWu0YXrH
g2sgjh/24Zikt67F09Y/56yBtEkdwJrdPEZ9O2WDkY6UU5iOxR7ZLb4981XECxfd
kW8N54huY6DUA66Va+7wmOED2L+5kpGrLq9DXpQg9DejXJE6+XEeXvTXSFjtWX2j
hboWYaFwAkWLA0yuSSXQ2eOpwp3CMhjdF87IkdZxULyGVraqzoWD+ZV1GVCDmH0T
7z0nOjv22RQoDAPVoa2TySFwlT0IZDDANnoT+0VyTrWZqXuuxXbb1BfcX9xDOPgp
kPihjyrQsHrPHpixsUx+n2k6piKxpjmoC0tSszPA4skSsrd1IkxqhPGNZCX9hle2
1LVpwp5BEzYHztB1pEZrX9YICGi53DdNxXXASMNpSSzVHCyQ/iTxfFAkF+Tq0NuQ
C1NrnxBpLuSAp+8CZ4Voap8eCOdNkDKNnjExjtnme0GjD/Xs+Zh+yYgMQcwntytk
K0m7RRw4B4QMnYcAxqGwQBSURPRPSE7eeElFfkFDL213FtNrxzB+G/erbRFiHYeh
XppfDpmZPWb5Z8I7FGa6RB5tLrJrQjxINns+Q3c/9JLK5HI/VDyGQ0YUeWrhkUdP
5mdDNXPplDJeG5p3XJUdswADSJZBcRE2gDlcPQp0f5wDDDgUAwgRxhVUpWAmqYop
RDHQxFbdfLxb7Dwx+QqY7xoiqBHqwHLFLQH2UjRW80t4++5QSEJSZQh2aoU/h1Co
5czCKnJwAmlewNW2Om3wLFf2LJywGlH/uBgnwVuYSOiESeCc/KP41umABdwv8XW4
A16BNXyMMbIwAIOmmzpJ4iSKw8nogIMEItYj2oyOKFHg0GB4KqQ4szkw8njgDlwe
gwGlBl0cl5gnrnuxmYE1H/2YmdWhS3MurimnfRmDZddMkBWpr7uSyZjPMc9a5Z1d
VAhurqH3c279/R07Rq5ws+IGLHCw5MHJuvtvq5ng620HZTzHoCa/TpoTTJvg4O4H
Izc22yuA8pYLAlP8P9rRq6UH5OvqEO6/suajYVtJ/LskU6PYWyRgXbLYYoTmwA2C
Rvz/pJbm8fjuntFGTGNYmG6fvG5dcPutf2rk9ka58oPK9YLpwXNVC4pAHMXH2jtK
BHXh8eURxbTR2dKLstEWt5Nl1VrlmstIjhxMF1seVc8Ts5wJGnE8QkhdvxxHbTBG
f441fJI2fnnFyYQ98BK4TnwzFltIOP6mGumgMWpwaQAxeA5JpvglQ8oxVmBjWxVU
Hmwxa9wOyYuF/vw4eJRI7MAUnOpvYF/seCJBA1ksD0VLaghUPSQ41a0yfW6TVhOx
N1i/po768D9bORujF3AVZSnli8TYiDyojQHQBjkKK1eDUjInbSGmbazaIswdtjzk
nuqPuA4YpkR0dIcXHIf48I90RQHTbuTlSrPs+kBzORxxJ3Ibp6juOhmBGErawBmF
C6f5m+iN0pvFltn+2m1DPzFybIi2irDn/4DJyLzeN/mozmFb8gdIX//8artc7nl+
WPT77BI26uKwPEhEuMYj9vDxBODnspgKa+Oc9kIBsYvoU3UjMWMUvI2JzRyKRsTx
rzlW0MEF5aCm/A/+UtEQsijJZiCS1VTLfSVjo1gPyZSHtTVTFl0krRPKOUivTFyh
npiW3Wt8mtrlVElajfyqsRGS1HqSP04LkerExsZb4oid0981QAbsUs2r/G41k0pj
Q7++33NRZJPpkPtQr0iO4HTRJ4zWS+Wkny9qIKc9nuPCCKO1XTUB1+e9TA79KmJO
pAbutbX/qJDKzDxYqBlvcBWkDkDI/fdbAV7GdUNfyOJkFV6ycQxgedo/z2WvBci7
fsdfxYh0uVjcpuq7neZznkkh7C9QFcNCq62Rc2jxt8S+w5CNDifOJP7NP6shm2aW
DvNYgczoCxVzP10UPLm7ualo8w+kFOMM9GffanSKo7Q+xnppYB7NmzJT3169NBtZ
G43uZUeH19kSlEQvsMnWODRZZZ+3rsdjEvCDiYUTeqUxcx5LNMZtKztS9CgBcJuZ
hFjg0vYwjjubcKK+jUJAPA84hPutf6WV2H99JBLWFnnwbqT65YNTLqHu95bHCndu
SjrgT35l0S4z6KwYmgEgqZ9VwPHrTVs5v4OVI3iMKdIRbsgid/slOunWXv795wpL
vQQ0FDU7joTVxZGnHsi2e0z7f8IyIGroq+jpc2wnx7GKslR1qLgiWwzlh95dTLEX
v8i0tC05p+t6tTp5Wkw5nPdtFG7ce8dU8xltgNvxpVk2Dt/cgLZHv5BhTfA2s0XA
5Fbwq2pcMkDeMCj9NeZw1QvCDBJ1Vn7OzReVGR+l+3Rn407BRh7Zfp4MpIMvr+BE
iQ8/FhvMrEvyAvqp/OvFxzNWrLt7T6+i7dlZGrZLbQO6rTeqk82BESAK7AnBa+GF
QqnHVuG61WkzKjpqJOCHVO3GgBWB9bk9UssefFwMgdW033T+ceU+olvAgHRZEOjr
Wk/mgLH/UO0dYdx3GfVrZKBkn4HAbmzYQZPI27iTty4gh3ohOuVmAcrEk6+lbo89
kOfilwoDy1HsV9ngH6R6awe3R2E6uqt8Lr8i2Sc6we3dMWPfOy5hYQ978qSxoMTc
5HU2Ae9DcW/2lNrkJcdftHIy9lqc/pmH7zWAjNEhggQGrdCLJ93Ob8xFw8tnvnzN
AObPLBC5bU7J6c52GhQXYyYhYQPw2AGbzY+CRrY9bfLm9NGYUKJ1yfN+rrbnXS2M
y0Nmj0dehnJejLPrtBfRYJvNy9u+s4TjgGLa0xq+RyQ=
`protect END_PROTECTED
