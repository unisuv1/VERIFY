`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gONNjs7Y3EuFUfwGbSIb1bmLXa3H+smt3bdwYBGEJucVgWT+aypTcVWeLzDXoFUV
UBBCz8jU6LBRcZpVBwsEbR6qly3GoiZn/AOWoFubgH1LUb+p1UHRbly1jA6hLRBc
3fymLsxa5mrGNi85767LuxPd3vvmVNmqneOqcw9lTOMF12DI/TTiaedAykNOVrk2
oUV+cvMmiJN/5B17/CAG6vC/Kd/X0y3Z0bnJ+3d2oB7D4G2lfjUufI5shxRd0H0S
1gKkVPbrb58pRun5w/rpjGhF5LtjckUGH5aj7Mw6bMow51d5d7sGn8fNl7l/XFNt
fKCgaZ/vE+Bhi3zIQogPq2BHtwAVTq2mCGZqwn6K0BPQXIWlwq1iIthVSp2mA+Hg
sQhT148RaqeMnWsIEjOdkeJ+xcvBGu13oCQ1mLAnhOzrIfHzXTlPqo/dl8DuYrs/
gFM+35f5VVcXZy2kljxZa+rx1wMHPl8lhJaApRZpzG4sdHiZKdW5tXV5fE4J2sgP
ych/K/sSv1RmelaAkuIzB4khcv591wzgiFB+BzFQdc/sBPIp1/MmhdiO+5wQqjbz
zWbD87mzcIRWDmznB1z6WU6copHR79fuXEPblMLDTnD3gcw+/WePPZThjbjA/hWU
Ex6n3eW2BHTLQEfJ/lhP76WQtkB/OePDEQROphGxxormYnO1osWBfnIrtZ0mXQQ4
No/9zHC8ORqFJHbSPDIoKaQb7bnTrC6WB2QtgSajhWw+p8+ggvlZh26HjgYHViZ3
fD0CC/uEUXnyI48W1V1puOlwkeUYdAirXpmheNjmMF9KQVCVb3/qBkBgsD1LdLbB
5iTcVKVhfc4tXHstUnICOZNp3CPEcT6mR+PWNKYSQhX843Q0KHC2gmz48362HKCW
544YntzNrocO5JMcIN5wJtV2d22L/GE1BsQi9bpP47AV5yA6RO1grzoqBKta+K4Q
OGp+XpsnUGtSaIw6DGV8MM1fDz6qAIjFuXrq6yscxJC1+vII7sa5Cmv6wAGuK+nf
UKCGhNZaE4M12Ivk0q2fgrZL/J0Ougi68a9UPPbzAFelePmP9FMeKBP6p6qzCsVT
NlvwNp4iYn2SVAHTMT+xd/s5du0krSQDbARPKF7rmTdSOXFwxq+baIxxWs52imHj
XEPKZBDNp5HBS0jjoNtY2O146MAdxnMlIqZnGfv3L7yFTA302mt9/7gFyr7RF0FS
H12PXZA0MN+m8UHZ4Pmy91e85WYeOkB8Z4NbFKo1c6AaV9XLl3SwB7DfKVyTjy1g
jpkY668FadZRD5ZccvrPQ2gT1dlYRd9InN2bZwk+BlNnnxIUnPtww7vXPZZ6UxbW
bxSyd2GWq2kWds/YvXhG8XHnkkHdoCnkQQMfWVtkPpdP6igjRuEfoTXWLMzeVeL1
AbKad3nc2TRhkKEuvjse+bJfCisH3mDV2E3r/j3fsaFUA4r7HSNB31aMmlITfJVf
34nakr5XThMuHNXhqsft8H4jJ+/cHV38EttPysESR5t3Ng3AZX5kMWvqavCYGS9Q
6FxZ/tSerbV8F5kOTNL5PGsHbyR+yJPSPWWqgE62VuKViIReSCTsBQ6ELWujhKTu
f6KTwMZdcaa33btJk982LFrOEW7vI6hpTxRpE2xtS/8ZQ83feytLa90iaH4iew3J
9cgXgld2TzfXnXaxLVUkZbr4SrGP63G0oZoCWJ1GTtR4ifguYobyO9yrjFrc9mz2
00djqdT0zHyMlFLaWRaVTWxfCUT0teuzvPetrGlOhG1osFVoEf1jFWh20H41OlTC
`protect END_PROTECTED
