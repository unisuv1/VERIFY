`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TipmwpGHQFJu+q9aPD5rVmX0l8RO+grdgmlPX50lucC9+OP+fHmuvX70GVNNIiWn
jOD9PNg3Ksb33HRrDcaQ3cwDj/qQiu7qdwdEhWDkUbyu8Yb1v4vW1ohTkt5TBdU4
jDYmWlJj/yDQw0nkNTP4nHK1Z0NKzAR1jleJSDwhelcCOviRHPxMfTMhbDzFAf2V
exZjEpwJ/0ZLiA8rYc1CStuSYocZV7aahzJx6UoInsLgdCGlSXSkvDR7B8ox6VH9
mpeCeO/QVCOb06Hj/2xZhqk2md05R+vA/C1ciCtuLaBr1WOIpbeB4epMzUdEug+i
0A6Aak9gyiDImHt34Oa36RrESMoj7jcuVgnCZAD0asXzrxsX4wWnh2J5nkOlfCeo
7Nk2fqZcN7gzqwqkgvl8rViWmJGuqCB8iRvIaDrDc5F9bTbAbNIIi9yaqpenyNpJ
J4U0pW3M8GrCcXYDH1CxSG/rEDMy64q2hEkGcmsFtgRxMnIEpP8HedXOzSPmzcGm
5IYmNrVS9ap4JsTkI4xZQv1MGj8OOgNLW+cOpPlCQeEfrQQmmpT57pabodJDJ9Uq
YkgySPwqG5xCsauc81F2I3JcmL4dRgtgC1liM2LxTcAz2vWDQw3umZuGh+TyO1HY
PxHMCGT4JljB1xcNjYhcb+jXnBC3HBuDnin1KOznhEi1yl7XcTR80lJrOmEgag0y
PX1GstjWTtzWb4EEnOWxcviS4gs24QO2os+ADBbQmmWp5dpQmNLHP8ypmKjKQ6dN
Trgt+FNCnO3gCgspfiS3+mX7FnOvrx2t9oqo0ncP4ALbig2oGddafMqqx+1xb/ki
7VXyVP9kwSBrjh7z5ZqBfYmESAwgNPUsGzyhWdrysYE=
`protect END_PROTECTED
