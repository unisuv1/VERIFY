`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
SqHfMxcRs20x8cGBPUaOn9Li/iVA7sBPHyic3T6FQkQyHpzOPy4vHFzL8ZmNXv/G
/ZwTv5f0U4e4Y0+h878YIYzYPiU1ZOyQcWlWnRbZBEJ3BXZIe3yzEqEkJctSwZM6
GS9AyJZB/MOCvxxszRyECeAbLqvIQjV7q1tUu/wNuunlpRoxKOfVtQlhhI2aTMy2
Yv7qLa0CKKXdg9NA4a4aym/JozeZuKdWUroUkluhGUbRKF5XIGVkNoLUZjSR7//6
3Vzr5L6dgV3ktwHCEb+IvxzkLjwr9zdu4Q+mOPgegEJI9sjZVdI6kw2yNJTLkz78
F8//EOFWgPP3Mxy1K//r/C4UYnjrY8/lA2m6dr///Eghzwm1oise5qhqeHdua177
CqfsGQl6ej3pNMqZxu5bnhGnxuymH+V83u25Povxy7OlzntWyKhaJiVrwJ4CA4Uz
VgsXXRwzSjJPxAaxiwYBLZk1UYoNsCr1bgeHBgH0mcdQIIxAZDXX4lKZ7e2O+VDk
pmuZ+sp+uSvgtJ2thlQ/Z7qJBrV0F6vcWQWYrDysE9uofvq01CmrNmIuhh+hE+c1
yWZLpycjU4eXiULsh74q17mAvlBwTkSPmSeHcsLBqQRhqwgto0FJX9nWisJ128yc
9QqK4rbYg1ilGnGuyLErTG0sQWtrbvasuqmQ8hBXXfZzpZwGDq+0Cim5n1Q9H1FA
489t92AkjhF3dsjCsTKDYtuKo9ssReDWsiu6N70FHMQqBdrgt6+s0mB3O6g98Isd
ogyH4JkPAOiTywyax2wNZkWjlRyLbFOmU6Dx4OgW2hgaCd0Pdd3DVyLsFUOM9FXD
VCeHAmWZFqpEB9psCPZrl6JaYytmQd/uTF+ymmWRqAocKWrRn0UaQqkhGdjB5Yz9
Yx/5RvWbV3ib3Mep5IuMtqfmA4q4KyctF3Qpb4J8JhZR3hscJMvUgqMAaBm77z3j
k68WzckNPzR+7/NhzFy6eR4sM6rpiWsgX7/3YlqEBaNWr55ZIJ/tHY8mQ2IwrrwQ
W4gu9DCdyMR9993/STxKbgF9U5ahyHPJxsnwRG8sBfQbafVmHrSRzbngqiflT0R6
NbLtN+ggUmijP3oV1rajcE0D3d0aX0Q1hYjjgH+MvRvFYxKBZUv2Q2jKCWyR0WkJ
jfCafc1Z6brQV1FtN16iHW2rbe2y2S0L3Or3rajNhqa8uwbIdxR1+TJN6MKV8z3J
sBmY+djZviCmPzL+T6DdI6brlvLIdRRYbTOr+2eYFjY5j/pC+/D2deuS8b8svqSM
`protect END_PROTECTED
