`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YNDtiM20nJEncY7S/Uo/eoZesdvoyrBNOjurl4X/Q5z6OfuezO0Xq7GvJivqIMuM
E1VYRAtILYlINeGKnFX0mnFKjxobhls8DeS6WhFdhCkjxJy+NJzkd9L4hxw6D85c
r36FsAtrXIvmK/eMEke0ng2pPJHQW6G7pOjEiDG80zEim40UbMBlddI6QcBukBib
ab4VA7+sjEDbED36l+7Ef8eTVHhq2zGAwVghU/4fSJLSjW1cpDVHF2/FcpGH2UNk
/3NEoG99wEC42ewOCJLDdQTP8aGXbKSWQTUDDbE5hb6KepCqa7qEod8qgW/zZZ1/
CNbpUAa1TK4Bd9UygWdyixAtLJ+e0qBkgfe31JDhjCwUMybjTp+Ggpl4J95wANeW
Ke3KHYeyZ3zYl8VWbPWGoHiBPQ4h7Oc/6krARaIQkml1b9DPdI9zWtewDmBDErG1
EaeWtaJGIzc57s0M07BU93MV9pR76VTqoR8MQ/KHFWW6mFbx9eEtGk0Q8okxkedN
hyf6JesLJQaMTbkaMIvx7gRSO4POGbe2WCjUavvcDzF+q1fFeuCI5gnJPwVBO5TF
444vjkwaE87rqfKaff9I50bErSQVc9oZoPG+qxJZudk3cWUa353PcaLUBJ5eQg7L
38KKVxPdiGor+beHcYyfaJAuJtblgV/zp9etvnuIQKw74+649UoszlNBbptTWLSU
Rnn8Qkic87xwGvorHYha88tBxrwG/EDBSNnTd0PX342S4rGF5aSA88WoRSaVI/Nx
eoT1JZQy5M0HH91LiS4S9kYGG5qif3IpY1AGM5VsAtrSHysWI4DXwZCJF9hKWDB8
97jexOCcGZesTvs4hUXFJc3iPCbMdutv+IhIQUFAE1Xm719TRolTGEy9Ix1qk6z0
cygo0/ChM2NnD9jN/X5tzib3yBcQ8qicz0vcta7g/jF3ooyUkI0ohv1rqb2c/Iy0
x2X7lf02vkRYtqitOGDW/o+eEX0XLVqqtXmUWkIlB6GGOMVxiW09mOJR6Q+0gYas
Ctr+Z41BAfw1//vvD9fXFpLfbwg4rkuzlg3vfSFix06ftOGWGj304My/KU8kdAVb
jOrBnyb2zS1zikCuitpDtIt0qh7pjkzTA1aIQQCwoZqRSSSEN4xJ8xUr7tXlPUBD
cl/V2YUuNSGyelwfyiTEper0erxIpx55oYPQNwk8KMxXiYg21/wnhOAMUCRDP1AA
6+MEsY4Kd6b6kZrsJnDpbk5mWLC81Pw3kyGwQDiOwmxBpgZY7Gi5rIM6G+OU2XSZ
4fiXOqvO0jvXD+ywMdXAVJrCamvFO0xdPzOO3chABBHJAmCDJpo7oYYLY1CT5VjM
1LrWpRiiBfB4NqSVQHtnJao9JxqjmQ+QmyseO+GQ961BjZDoFKtnoD+hqUBEGLhR
r2SX0NIeGWd9qMTtX6gFfnEdcmOLbhQ1OK5/OgImj5gr9j13KOYq+fNyRUI/Vgbh
KN3tXqToXA+0BV++u8ng9fqzAiVxFCt3yjtfHN3MlkzMyL4BsLCIbFQedElf7lo4
ABg1wLXyKSjDJZQg6LlTE9ZUWJHty348Fk7VL358FHxfg/EsjfaVGEX8Ffh7P28u
DTM/05yx4bLhpKMwm/T+PLTXaQImmA0corHwjs6B9TOKfDQPafrwrw6khOs3b7Mb
C37NcN7YU2JSTBfU/Md75JLwf20R9mQdUB6U/Tvm+QJIneIHTsp7CFwRvliEC2h7
7p9p4mxz+uq4CBDmwszWPhnO9l0N4c4kfkThvVWtyllD8cd8w9ow30EckHp4s+Pd
T9LT2GX7+Vtx36vJ9qGEWaAQ+rzd9aaGD58dFXu7pmBH9a53s37Awv3xTqCA06oe
BGjLx7MuBC18VXHyd+kigkmmWq5v7+6ywDF0DdZQtzr5e+wJcE4DHkevCEQevIXK
UUI7g7kGwcYhGfJXhJC3z8pJhT35ufTm73ofU2TuRqwnXlu3ux9mj/LAXw2rcCrW
ILWcTIxeF+MmUYeUo5mZyBGzGqWxhzest0NAvAyX0LWEzzKL419DlV3wEDNt9kIj
wHfCAB9nyAAUaC5IvCKgbPAN6a/mLMLJphrD8cplhm+sqaL3/2TXscKPLCXTqZpo
QRpAniIoujC89x1n4Q+Z5FQ1JmcV6GiY6NRjBwfDO3ejf9VJIqGW867o5gZd73zM
CdMyobTsgDvU+hWKTLUmWaJgnwf2oI0zu/lKHAkVQxzpp9V0akUbZ4o3E8+Gjn6h
9tOJIEIgvDOeIOix4XKJxYF1k/v5oxOE65x0AQ1+5hEA44LkVbqUE3qM5ahWoebn
37C6/M7BK8HqIdATxEIRgdsIhkROM2GC0ScTh3mDirIab2e/LaK5Zg6zD7+CToQn
fvk8lFyEAFsZuUeiBTfZKLyaMEJrOChqfbOzyEKs7kRxwZFx183CayBnCfCdgdlT
GgGpF65LnOdvPzQpNssSkbNSay8Cu5A/KRc5zk9kELE4VhNc4zux85MXB3vTBkHD
F3/q/K8Y56rqWKbOV8Ods7YkEO9vDL+18GQytLg7SllAnF42VkYeMMWubcC+4wrX
WbATLgmzh1Ioi3uW4cOH2EvX2aqizvwG9L9CVzn+61niX//RYWVeV76TqlT90f2G
Gi7O/yBkyWKGlzwkFvtALi0U6WbOg7I4q9X7HElPpkBIbU7OAJEhM9azXfnuAWZ0
UAp+pNDfDzXBi7L9/aLOERjTCb/Fdc6aW5eJBStAJnYDjpdz6bX8b9Z/TL3B2JPM
faQRtw5XGh8c2wi5+cFu3Ey4OlDnFLB0ATATwRXcAxYan5HAAT4H+ugAGNKX3RFN
cFDK9lPlidn0bAz6Tee1xUJ8j2E6Me4aawtsECzhiMe7z4bo3ZUgZWPFBJXiEX44
UsMie2Qy400jsqlIlQt60r7XRwDqAANVpnV2PP2CEJBWdfBd4kFTw3Tfsc4JBrgz
ya9kWM8WIjy9wbpljmbwjmPdsr+Yvzt205XUQOLz/2eBIKy/30FG8nT9YcUJiy9g
tCF/idk3viqpJsOxbMQ41zPfYa3EkREq3DELOZ8KIAZPehgv0O24BBGIqdp0yIkM
/IVeUawG0YPxNIanAsAsxRgDgB+gXoSTPZuw/9LRbFamVvkqpo7W8gWxQh7qmHXv
DdeLZ92d6a2pO2rY6Fwwr2aG9LmRZ++Ina6eyRKWd1r7IocwSOD+AkrXj+eD+fCd
dIGrworCsqbFpyTcAs34DamZOpWHPu+WiD1Z00b3QzA/3XvHWMN205jHjlxUEX7d
N5aOeKQ658UP09wFBsN/7TZeliHOboCzxSHjnAowbBpVTKSYlxFiHox3ItrYK/Gx
tEVuYBHbUcXFUqIAv1h8tnR8ifSBJFOZxbsHBLWCCYkBC5cOLrB7DA29orDuzzOt
7WFzlCUZpSqo7TqPViQ+Xgeo66iJhriVemOz+xqsUoBaLAklYknRO3Raf8oFaAzc
VkbNzc+74Lz/F9kg7nVQrIWhOd09DWZLJ/yM8IEPgBgDDuQIZt4bynwFdvmUDuas
oGktk+RopP0VCKCaP+xpNJvpbsdOuqmkjrdYLbMk8uLsZ97cxF8gSOEGIInt+qbW
YJuMGQBWwyfLrU5u1bdgUWIEIJz3M4g/64dI0TShYmOd9s9EwyYZVKts/S+lUWDi
FADZsOqU5KKCjDPxT3EccktkqcxREV803gzplsFcn9sfVvjGskuf0ebsWRFBCgzR
8EZtS1LFzE+b/WeDg1E8N2l7Ks82ylpMubVYuLahvnVCNzYQa7v42YojYD27dZVN
Tn5n1hbUSxPesiuV+QmnWYvfVa4sT6bTiy3ThzMf/rqfRfa25BaX6mGFGiBA7FYl
bMAD7vsuDdZ95oJ/h/65LrHxTlntdvZHMC4yYKFM7l8cz8UFz93vT+OgynUnjkKN
zyJwa18w+d1F5vC0YkTWLJo0HexFSOe6bcmegCGnH895AfS+GOUropLNPOGXDHKr
kxraxXLAZwtubLhBER5kJ0MB9TfcNRyve5eUZJcTqxZzXA/03eJrzE1XEXQHw2dh
iiyDVaHm5FIgBiJcwbOvXTpt+rAcIy2JgSfOlXLtnnkCR2o6vgvT6z0PdPPMdcyg
jlIBhXNXBd+jgPH518k/c8VzkS+r4YK0aQOhi+0Lht+yYf+32+xXPmpTzM1kHJ58
17oPoEhWh9jaYppxddElkU4CgFgnrj+o/rR05LRmQnh3vuyjdkV1hp4kVsiBIkyh
sAZxPR5pyjj4RpeCL9fyu9bDRRfjGaHUJUR2Q7jqPzU38digDndcsyr92/t65UWt
Kbe7BSDYqTAsFEPkUCgkG4BbEX6lO1pzVq1k7uOiHXpGnobjuL1LxIM4H3rE053T
eiZ9hblvCRZWHMAH10ZfGFaOcjb3fIOhjV2lgKZkUTujuebVi8kF6xSg4Iczqkns
KO0tjIfpM/dFlUB2odtva1MSd+gv7zIfqczI8yEv622DwrQtczv8h9pEUWgf6dPx
E4IaLlBX9Ws0b2hclqKZVF3UnRbbw6PsrOPFA8rxFe8LdGsXa1eKIp1JBD7CCv6N
wUGBOCLgZ0xwegxdglG4nvT17Wqori3zH9gWfF3OFl7ab0A0kvkcOPMlo0OuDF4e
0F7u4oS7GWFMhLtzeRU2XAFJZF3tqEHEZEmJXxCRWarrOvYMayME5ZF+KhRQdYzM
XR/8rv1xOMMJdlTwmFl+jHBGNrp/Yq76t0pjWuaIwAfXOrcon6KQx7R8oDr5Jl/a
cHpej87En18pfgkwI7XJcWnb77UGs9H4ZaczdB0wK9n6zeUrcbst8ch44S83L4Yt
Jp+xtM2uUlga4kKhM7WJLo+ESeKluOtV0LxzTuw43ZNnGNwcdaw26SxStxp6zdBS
Y0/Zuk8u+Lq4OPync+6YeLNBK2A+9iEdGwK+nVHWIUqE8BZnCARMj1XwF99iPH9n
a7a9L+pYYA1+3pF6EeSQ8y3gkV2bA5AIgX2R2oOdxma3YVk2+4p6j3MBBxhNLfko
M1sSmfrZLLyQ7wTyQnZR3nUNZMECgLopeezgZM+1/Mf83fidaUEahnfppK/IMYrG
rnoc0mgk7NZQE4Knefv1OY2AhDtpJY5JqnjyjgozfhhQfm10fAw3LkvrkRRGXQXO
JB7lsPuPcVWAVsYN4k8CkOiBnoveqgbD/cyziAAZNSUnHXcfblPzcr0ZH9Yt3BqS
PPgwQOMh5xpVjEQR2ID6gkZ+hSG0KCcx1lZ7W78++a+0vcfukQKRC211k7Z6n92m
L5S7eVdSFzagwKQAHznYe2qDJuALRLbDx8E/x9NK+VW9C6S9f+mz5mt682XGqc4a
5TRGAiLGFErRbpI+GuRsLFrbRqLN+yTbweUZMr1whpOHmsxPGnrxGY2iPuP4y3wQ
8KsSFI8piL6BQrB5bGhHK5zolfyWdOQRgJYcM2Ms8XuINIXe2W4Y+qVtshx34muy
GKqk+GRvzrVtXE64LfJ74hHB2bTkqXO+iP/xiaQORy9jPT4rrm+71HSn3zxuc1eO
iCY3Qv6AsjYy1CqUdWpNPKCeia/k26305UTs65Ciy3ASsp51pG12Oy3vh/wbadJy
XCuOZMGg9dTBiKi7NLRtiqOmtZP9MifhWsyEorYVxE3uC+seFIGVqvlidH/Pv7x6
mDLRZDhZ4jkUh7IZehN17IlfUui+mSKz18932WMXFTK5u/fIziIk/+ox0+s8o/4C
mzh+9CylzqQSvQJjugn/h7qWBDKWDjfgzlWWqilDQPiPRwfDApFBTXrzDri01lBJ
/IQVMTqRXSatITmo+NbxdTljtYkN+Rp6B9TKybhpbnqzF5KXA/2BjgVDCllDVBtN
7gNYxnPs8dx3+c4IABT61UXsOMuj0GLLPEpGdNqjnXNRbLfDWvHMKh0+xpZReERR
ksN/9EcoEWHg3EbxJ/0tlQLr3nFVHWqAmN473M1rbUaAkvDvks0HdTXaqEyvMdMX
SL0FX81xZdoKdGgiZ9ssOt6L9CM/BPYO0Gn307NeqzB7goul8YMACJkKJqzFJU1R
WzgPeM+wWxSvrqBTX2ZgdngjP1vy1Usgebk3RR5gYpC1F4XePSqBYU+Xbi554hSU
hkYMQGFbMTp2WuXxguEb0CpZqNTlckfINYxcJFEfOZCXOCTmtHynD19mca3Qu0eC
P7xFTK1qRo1v5bwEMuJUZvKIeMXllWLoNaApqbka96jI9GzNQ7rvgBIC8eJzADl0
qojCZEYfGYpNS7z+LYaRrULgIbzRuJuFGTjNktF3blCRkutQYBx+lNUjdHdyLT/T
SCWWGJXkZmbljTG/kvMHPwi0Vs9UQfrBgw+gDHfBh7PQ+lCBBgf+jOTYUwIuO+3D
oLxjyif2qvmxaBia3LJuj2Zjm0o7HfiZhoxQqi6vSmNx+SyHYuk+Kb4Nxq0I0JBC
2j8xKHS1wnYf7oYPyBp1dZPvoSOF6GKoKFG2xp2GPnMXFLqEE7QLz+4tcQKW3d3x
MtbMv9t83afp3GfDy4eRrCBX87R1od5FwidE+uNXjMB0twk8oXUYLUN4wsAbkRDQ
Utn12M9PlLCjicEYKVZssE3PePbvhhN1b38rLhEys73gBMaw5CenBQWJ4IY/2/4B
FZI03XshgPM7lV1jtlGoxdovDr/GNjwqymnbBWW2Mk1KaVM0gOV0x4WU+Kk3Vxth
jBVn8rg3y2mJFA3de3Rx1y06z6kt7ydfhQ9ffTmM3wjxSW/eFn6A6NwnIgfpgY7P
/Y+4Unzn1NcaSmJTsZFJD5aK6YogIEqufY7DHheI563FXume+saEx4L6CIfT3d97
Ca+L+gcKI0t6a6rhM47ifkwe/1/wRo0syR4vhtlw0hiSDetf6k/BdRk7Wlbgd2eL
hNx88bn+pDnJexNeR0G0PhY7DSsCx8TuYbH5t5qydWuIhTgpRJvt5Gudo5F5song
+iOt8TdqXA+8/sKEyFyHaMoJdbiMunc88SCgq2k+72EAhzOUT/QWmzI328EWn0GY
j9ibBL/S/vdVXF/L2LzvSpeAO0f9NhSXbByQOzx4Iti9mUlNOyNccPw5j4beZv0R
C0Qk3mV4dvO9Y0h/qK6d1U/ViOkRsIVZCTeAt+jSjl+i7u/UEg2pG1iogSCov+Xt
Kb+BzGnHap6ItfNWRglnELfBB0U/ySvU3dn8yG70xiZHQBJ/cQLRmixldX5X4UeP
48f/s4feDLRPUvqMLWK/zwt3BdGa2jNC0/1OQ/6oQDqQ6DXJPGQ+q6Wgb5I37JwC
Lo0bihxysUzla0sGEh2RnS3jqAe07eXVeRW9DzqOt54YgVUFYJ2aCpjnhLMpYQAW
tLVeXWO/48CoW0NIzwD6JKJS7Jw2TRtFAESi/ik7r9qYmQ+jwoAg3fH22M9ZDcPi
/s92bmtNirUyreUIMwivfElaBY4hMP5eAXvMCci8CKqmPpC3wyfid+xW7YqrzLwp
Q1ak8NEC8gSd+oZH9iD7oiMvL1Z8oUUrtcgGF7WdXGjIEPoiH1L28bhusRVTy9dv
2gCMoRIW3Mw7yB1rzcCMbs4rrFu2Xw2iNaDPPxDNAwZAlixP7gqUzKVlkeeL7Mpm
a0KYbvl/Rpf4YdX/FzMjduhyaYfnc2jLH8Z11QjfPeIEBlbBT7ns19x1aZ8BPOl1
Hafh62RzaRTu1ZShprHN0pndujm+RGptbHWsVOQ/mM9PuNdEruX5F/1aWRT0hFs0
UB2FtKhJA+IRN2jfmgnj0sh6B/lKnefWlS0lbHWitOr5T4rNlZjN/YDJAZaEsCDf
DmSrXA8oHu1JtW3s5uInjsPEz2xnj7v/REJTRY32CffbSnkAZ15K3wls4kR1yHVT
06UQ2WzlAWQZu7XzH4UM/MC9ROgd+NrtPjbq2ks7ier6yA2WJ6pYdNx0nZFn1tWm
AAxMrBIzMeVlWRu9zl6R+NphXqAHPXmnzrTGdQnbAXRuXoI8767DoC72TtPhkjY6
dsOwj1Ahf24g4ft1fjFW6TXOjPlVU4lYhMiaMceRb56lkDwHYBzVI/o10Nml5D5Q
7jl6irgSRsOrVqtyfx+THCzN9q0E2k1mIAwax8xPOxk3Ij2V4MhnGendtn6L12x1
MbA/EeEF/7ga7GSpqQ7eEAUfLYysK7q2XNR2oejJojNWb40frB6NfO3ZxUIul6AH
jBQjIFYkVtalGPFk6LK3kq4kkmjqVcW3G+OKMJvkCAZO+BGfX0eaKBXoAtH322Ig
ELn3CtP0iGB+aFjRL+A4HnJZFsWkc8gFZo/TlYp2uiS/2q9NB92mWNp44PV6x92w
KxPinc+G5JaG2zaA1ItKPsRPpZqd4WKtotmeNcy+ATINvgHXie0xu1flgeRdl/I7
hhvsJFK4sf6a5LVYv2MHXHcO3QAcYuy1cL2E63zWXdgkBnQ9T1pMGvMUqMQ65xGD
NN2hREAShUi7sXcsFHQGWWiRSvHNyxJKkDj9P4Nao7q6V2I2YbifJ4ZkvQ/jyYr/
YNWdyB6IKgvrSw6458pcRm9lxzEnicYhvDyG8HUliSYSxa/RNdVCfrOfCiALyPOn
wi0Q4KyBDUR7nlMLEda3HmAYMUhkNfjMc507ssr0yYugrw15EaEOaFdtIZ5dvcj6
XneEU3EmcAHw6OISHLXAYKIZk53E4rjx9LPwKxGbhSPQSv6uAkwn5BcCyY820KP3
7FhbWGY8fu4olYDeRk3ro8Q1eW/26FaLQ4GhSreI9D6M1uaaB4VFZTdqjjbMpWOy
sHo+r17w622H39couUpxpuhyZVd99SbiZEzJ/1K48xg0KoVQQbzmTtCERfer8FC2
oPtuDoWVgs5kMKpNeHS66st6PdJy0vBOM8T3gsEMBldpNMJ+oa/+6MiP3za3vOPJ
P8fG/PVlxaEBTN/7luy1d/0SasuYNaX0P+k1k3dVmy3pRp0L+/6fvZhXnw7jdnUy
oaWwAs+eDNI1B9XVz36K3mSqevMbJpDpC7r2r0+0Za6LFuQaD3El9KWc5gAx7ipL
X81oOo+ZKe3XRZfAg7bB0EMTpsbxxKr+7cOBIFd3ecYwHIHR+pHkvo0UGNLBFV1k
jnweRS2+eTePfqehXk43bTNBcitKT6o7t2gwLybIumIFByNF0FZqlpWw6kHLOvxw
HHTNNBz/iCcs5xK8xjMaBbUvlGXInsL7waVk03T1bQqYekfffzFKf04ywnvNFK80
1WOdvfZ00PTL210GXTv+4HC1/eFzJscTfg2uCPTYlbRxR37g+NBd+Q1MzVL/Uk6N
3xCFS2JdODfWzlEPEtlpYsoFkLNoOqM5OSVkSs5D7Nwb+c34j4U2RTGZu/4CU2RU
imS8RH8MfmN+SQSXrAZmrt2MA/8DsRZ5ivkD6dg4eJ1jAujIkR0gwee/WJWn10E2
9NYEHJPiX3kfy2DMGb4zoxmQ5e2U4nk8zwnQpwvrvvVUlSOymKx4uKUz/s934i3n
F1G0SnnBx8CX6ymWpFSu1mPbeS9arleoUdAXG4Z+EY6Yj99OsWiSz4zeez/ixfOQ
QNTPaJdCXNbweU57xTI6bldivevXyOKCNufEgq9nXvyJt5OWJBnxCro+OjyPdB1u
9gjMS70AlpJxVjkRRcMkNIe38cdj6WIqSgpgGxi77H5xP2pFK0+HJPzGr/9Y8pnd
hTfKhP3XCIzJOoYxXWsjW8krrCI26J8b/0qerp9q88c+ZvsYpdTAAJlMH+tUcr+F
/7zoiORbaFZLwIZ+Dm4bhAD6w48ZDvx8xob0ue0hPE+5YCI34Ytka47eXTcSqtwa
bnsCdNcmlbj+ucXk+esofQZwfKQJ2k8sfs6gr5W8UHXbvrtoVrZH/U2oCcZ2/xQg
80jUzuUMSSbG9Cf294yL6RfMvH/zUNA5Y4KrhvhaDJG9+RiAanzwmnCxG4jocn8y
STMYrpsZE5vX27E61AJi8pdoO4hx2j+IxCmLmCilCemDOC2WqPuZ2B88Tzc8Xc9H
y7Efw/5tjlH/+8a0RYZl1aVkmaM/7O57nD/B5dFGEFgzvhtqPp8T4zsGPEsx5uqZ
xIPXnckQq2eABUfM1BRWYKZr5wIABh7o3SH2eqIlTBig99BfD9WB5/43BOPEKtL7
F2zhUce/QOpUp3PyG5BhPmQUwOYWp5elMlZ5DPb3WLmauNTE1dp8ikXsXKslVH9R
k6WiICzrjzYpbPTo7kFUojUTyLzkjmp2QRAgi1Ve9uvK/gf4uxKrWCsliNl1HAfo
IX2kJsBbmy0nTI6huPZp+3Npt7ETGE4ycwI2KmixUJZOIowF2uDkCB7z3iUS9kon
WdYeOe+AYNFCuliQyaoZ9Uf6JlntbF51oxugY/0yQwvkEtcM+pYS9bmv70MBhn8S
pCGj8yLjyODbaHcLWA6x4U4blebC5oQG+khc1h/c1ssZ0ubJjN5Syc63mW+aEram
poq56SFCUOWG1pfgQJFBgPwDXvD6Hz9+AUdhf7cvD1Km2KI7LTwez5ISDWchW6tW
DJz0bXbB52wqboDuFLGBVLk0kDg6pQcZcsowT8hMH4IUafGifAjN41AUwKQxTaAf
yEZ+/ZivjeJMSKKBdi3/VauBva1KDedq6dufhsGPJneqpZTaD3BfPahj2gVONYeB
2sdBfydRZCweZwoQLKsZW8gTabRpb7Tz3qWePbyMvuBfo85O4OZeIcE7XAzKUcGD
hBocO18XUfvtFfS2U9AGPdo9ZSouDPNmk8smjnxFyYPTkKzrjyswasy+I2Ukll0d
Xxd45c7bu2c0ubIfW5eeWgcqfUuIXZ5y2n0eIQxhZMUHlzq929bd+URUD8s4zSgZ
H5X5X372iUFNPf78vqs77YJo0b978TwaZLWAaKNB8Pbgb9eHOInkqC8DsMU5zsc4
kT8AGAiup3/S7OQc4PcV9UNDiHsxEEt7XafkqXd89N5HishRzt/nafngKPCCuJ9O
M8Leg2i5B4OI4XsmFywOJz9VzRcLxUAaDAz4LlWanKLQakQmHomj1WsROuG/IOZm
+FNPpAEVwGKHX5xscEbNxT9vSKJA1SFwFlEORZLTl9n+lDCGv+qez1QyMQRs/MPa
7r2wC7eQLYG54YhrI6VezsR488Gmr+1AyEmOevm7PNOT56xGD3yzYFU3oUj84Kdl
oWnJMSUdyoAW0tr9vOCWSntxKpgPfgl2gemU12F8HMm1iYUE6gNzThaDpBkUgXOW
ruZfKyRBZi+N16sEaSOfs0lXSRB39YbjcbJQwfugDnLQ0LNMttP3TZBDdXrqVP9F
wf0d6xFrs9ArFdYf6BLqb1mF4jRBY33hZw/FL27c6oXd3QWhtjYJSFKsbw/jgHBV
uz3AFVuSfmMrv0YapN2x5YmqF/iqyYZgVb6dJuA9mZBw+vWeLHFsvEUDHpWUb1Qp
CBq5SwmKRNqTY9mI6iRCPp5C4WRALBY8mhfnpoLvkm3QKNkjAEOv9wMfuFGCcaCG
PQ8QPbz1DWu7dwkyJIwSeaIqKyP/YS1SyOV92bbKCLguHVQte+lyObRIkHWJg0C0
QVz6b5a0nXR63I8qLnFk2SQED15RHHxf4sn+xPlocRAPh1ciCUCFXeJiUEfBV1Oc
l3b1zxv3iSDkTqIhy3aeaPYz13P7CjSn6Bm5lIYIoqWpJPE04Lw3pJq3TE9lESHV
ZS/NR9Z165myR1p+pAcFXe0dWsDP0L/pQEYrM1rjESEWkAJhDohxihfgg6XADUA5
ikENkg1U5VW8bmkT9a4X7+f945KgETMbvOTQgDb3xFNM6lrGmSR4rOYVBeezWz23
ws937/vjA73OQYfqmkdGrWfTJrt0ToAr6uOoQWq+pfsB8y4VauinE3Re9CB9LDpX
X628yeRgv+HqwLG4bMRdKjznklLBnSBtarmET3ElZ6SDsPYlEDOo4OeznNhAb2nt
PR+LV0UvvMxX3uZWS33clHGy3JYH94qYuRFDUc8XMKnbTin0eMABtQ23bTo3TYs7
VXVAoiCln5TOQDOGssA1GocBU52dKxsfSQU9/wdRRTsEKHVhc5kFQwznIkWJjniG
QV8XFratOoRlS6Gji+NaBzZEeV5ZJQVAjMJxOILxNvRxQ/JEcvzAvwmggYqR4fMN
S0Wc05021GGmWj0ew7JLkf+z8KfCbY6s1uN8sdew2VY93RmDCiEKogRyPbsiVNDh
8PeqEnsl2dBYyI+wrpM1PnOZh+J/tb9LG1DUNypfLa4c/3UcZXgQ2T0iLqeJAOAR
3HWZBkAmRYQjYTqJni3QCenqWkQTL71jrM3frHROcQBf/Jjp5blXuqBOSQlDihCE
xUCspcqU/4H2igcGC0ieFTK+kaMQzwufiPjPu4AXo215FkgPq0o1JGowA1WF05/4
xLLQ+gTdbtq4SclztW9BhOXLne6ZL7BNRjHpx8b0Qn7+i7bV7lxeEzORw7uSqkDZ
W/gNYBVWhTV4W92iqboymco8Lq9E7kUI9bkIg/N+6jaPn1Q+sRlQtvKX5Kv4LZXJ
7arhUQzxKEJAtWSCEAljPZs19XuyQXZ4xx+5JQ1Lr3REdpiniIOYJ8wXbEXtb58a
EHCpKlSJHLekFASeHNLRRRMIQ82Ya67DS/QJd15a21uTys5IfDHFOLreVcQl4cQc
Xe/H87Rhqd4KyHsiBHJm2dS0ZggyYnoDBYWZ02k6r5bT5lTRstT1pOAsHxlGKEMc
/NOG/Y9TPMYbPuR/0UonU8/eifg3Cw+zGs8UTQB4F5h9FvlD6XLv4ru0Kcd2yJEM
8/kPYKeW6St3jo79hFSy47MUNOwWTOrMVJlOh0/tDmKGREAKZnPxn2atYqvxNhJJ
XdrJr3JBclS7FwSMeTFpHsIviP4abv562an96ukcw/4TfZO7JkEy2S/wHyQXKrlT
tTyFYKo0kYGZDjBwbGw2FwRH6VIVKqTOKj40msL54CMPudXiY+UJiIsXTMHJYDdD
1V5Fc72cufrIaF86x+OkweNqC3uhl3Hzm3dC+ikbiXL3QiVgkRuHfcFYj1cq15TS
JTbwcU4BV8L1UxAxlIiX2yvwkdjR6FGx0VauB5MeUO62Me1jJxB+9ws6CNuituei
DpO9AiX59zY+BYXW46t9qAmxB4i/c2zRBlJd3TPdfHM88Gc4nAms3lFhef/2Kvl1
TDUP+pUxbeyTodp1vSOfJ75EOB6j6jVpEtkNOSqloD0RKkZ0co0lO7NzvQsilQ5T
CYXpl5CsAfqhuPXO/oS1qpf/guwe+eZ15tiiL6PjI9Mhcn30WolzcC8A7auomtnA
OA2xQJr5D8jG4yzc6YceawaYYdCz3a1xaxlyGCbIq0u2uBkGDgoA3LsAdz1Pt7Ws
u9chDLgkjWETnWMscTcVQPMVc1zZ8/cJltygoErLBLfqdttt1LCF3NJ/J+yebFYY
C9w7gDHRC37TPMEF1IC7hcVOdh/pf65fP3JDYgQcKhfke61i8wh2raGc/NOpklss
0JSa9S9xvHV8EyWa0UG3BF1WmXXWwwi7KsQnPqfVY6eTOh1QKB655+fdky4z3izI
TPvcwCea/8P+zstrlGix5UXs6oaqUDWyVOYgP4Zmg6vM/olwuAHOlZ94FTRDmSnO
4iZRmTAfuHkbcA76wEerC65d9v4dIg3jJOlvX2WAIX4Lpf+JFs8lQa6Uc6S8VUQY
5JqMplM0a2U11uplyT20bD5kTP7SJHhQj2F7h6XnqKaJzjyG5IUNdfW34tme0xAw
5dPPusY29oG6gDbKK5pfYZ+NOuBzvGxdDnAApA4AkoL/a56iZZUHwajCl6h8MVlx
jGQcTwlrN0D7hivGXliS3NwBIpheWgJHfk/CQv9EtWhwj8zd9gp3O9kZS2fZae1h
agDc8AxG720W5HWm32lGWsFbpN9kMPkvcQNR7g9xaPEsuYhHwXeHfnjogq8UsDLF
miQRP76nWM/6c8ogCjmd0kKBBqWdctgSRjhPx1b/SU+WHQuvg4Xe5IPDApqSFP1c
EO/xFLdEucteK8zQf07Kp+JXgdPtMf5OECsA474j7CbhKhxyDmEquNjpLsY3hIR0
wumKJ1MrY68tKqrz3Dl9GomUX9ed1h1REdkixunq82PV7HGmZMRSIW9/Fj/G4MOw
ZxppF9mF+7Sz0MXxpYGQy7iMw9YYCJ8xddv1HtBOGCGwg4WelkwrZdll0+vEyY6K
N0piTzadHc9WkfA6Y3C6E/wO4uh1qJTmm4jfp0ZOMvYnZB94SkurTCzMYKNOHD0x
ksXJbtdonXohIopoKdehqDGjtWEsD07YeZScggCLrH+eNtimfVAxsx1rBLrW1WBp
hqmXxlB+D89gwzD6dho3pyzPs4+JFU8cdfigbSOWS8+r2bpne2k26X9nH8XQh+HT
m6CwHevFRdEEJaSQ+3/ZdoHV9dlCMbVzeCz6Q8wKOKbWgI6JTzAiU1zUY4f3KWed
Xu+FfbFK52lMYpBvb5uWYPyvy98nqIq7R+733Ne7rcEp59Q083810STOdfy4gIAz
yQ9NbzCeusRtQanhxrDufJWEfWlIic3fF74HCMRkd4hEonx0bGyiwXnyUrfvKLYe
uvxJmi5B71EUmhnVe9q/B7sFhhniD3ImP5OLxOZHXxekRIu/1kjq6d/r/wUnuKAR
5Ezz+gb5ztPFlLTp2vxT0K3ZzRrrji3oW+IKVnSgMFSDL2oQzknk4uGknrF9rlgq
AeE4iuaruXywOhwCGax5kz0utchBibmJFBILrwQaMP6jEC5bUeckk1Q3v+UtHrUe
JJHvcniaN8366ogbOM7KXy16PJTPnWhWEbVxZVlYHU6Qrvp4F+DusmJE896BVyca
nbQ5z3dblPx3gFixIjUYJSBpswOg0ZMLlsikzXOoD96I2hKLj4glgBfv+Gjj5FpV
B+m/ECUar073/8C2sumGUd61cBbbBqBhaLIuk9YaMPu7UECbn2WZKjH1x5Dx3Flv
saqPLSYYnnnWgs2uEgIwUQzUcENJxkgRLEAmSo6/jj/D6RBBZaWEhbSXPsw5Ks4W
KaCB24qJhoMIsoDKpezT9cNfgTa8fdezVyiNjOmfWk4on9WeNyUaJAO6oNluC3pa
VWSCamohgxHA9bZ6jikRxp7Djt8Wak8c5SJTOu3OFGiJca43k4uoHeSRlv9kNO38
kQ9Wmw2nKTM2uWyxbzdUVTgFq3ZAm897DTmcn5st7/X5VIWNrXELmNhVkSKx/E9l
AW7IyY+wNRFpIHrxcdLlzMy274YEquonl27ZcWgjtcTTS3R6oIpETA4ZdEJg23a2
df8As/MbLWebENgUq8mhIwbazjeTKRkTJIGxe4D/cXWExMfLjzY1tKs76hU6Lyqu
6sSGE+PvVVfh8l1ptorOAlIWp0ngb1q2FBlgGtE0YmzqiLHPdogEjZPP4dhFsB+0
9DslcLaqow5Wg/KoE9/ymEA8VdWxbndTSFN6/kN+TR8ZyXPTX8aiE/FZKbn6H+Pc
b/bzEeQJCtprRtHvjrornV9VdRdW+x6Uq/5NWoH2ouRtZPwy/DdVVJEHkej1mfa4
udhBpLEt4VtIyDnW5uwTGLjkC9Z/fC0h30opeiQ9+CN+u3swUfk63wGDJTCEo/f3
ct435OxKlfBRI/g3aXOTK2kqpPNBrWAA2MAaqbASlMu9qoXoqtMbvmzTuX+lVqlC
RET6FwisXorVX2pjRafyswveZubw3138bs3JejxRTQMm1YRwvGUtSk2fEVKOjlaI
Ex3qa6djR3t8AwHjxslCs5tURXcJ3I5jwY8FFQccTtLnrw+6fFoM/ldhc1myQ3T9
FFpaIVpJAfvEBftntkEwDcs5dMh9JoFUzLZkPLiC4Pe90tLdGKAULArevcVfzdod
r+7gDGCWaz+swbhzr/Em0HQudDovvaKOvQSWHvMn+NH4PhAvHSN37p6LE5Hdljw3
egZRYPXY0LtDeWlkgkB/mMEP8zlxO10dIZJ4D2ptzg2oT1B4KUzgk2HPlZaQLPeo
UFIwGHSGbG/LaEVbElSmYseaMnt4rFxvKOTeEJnU8Lxs4u2I+gBIViL7eExTj3SS
qd6bHWK2eQVT1a8mnCGGZ5+3JZhrJ2vhz/yxnywNzymtWAIwKQBt6jmOQCpf+lkR
eoW/sEanvsSdpfboxjDNMe9ZZOhcF8Pj1PC2zXsbjG4PgygodnvBABUnsO9Ufh+y
LWNsnTcgAWJ0IXQDXFmdLUwSYVakTt2eBwHxruSYuKKBTNRxWclFJwhdM8kNtzuH
NYFpj2VvKNfvxOqN0CBxvVUHYS3z5FA4e+4093x29DzmGPDsHF6cojEEEgRRavd7
lvt2powh9IlD1mgxLaIE+LFYhZWapnEcxnQQI4mVh4Po8DD+a0NzbnET0cOQ+7xz
abeDORirrXs+WD95ojxcvlf4e9C1uEsRUWWw23BmN/EbOQjkCowVQk2Bf9mi7nd3
Ju3lrP14YJEBFBw/okixvOUNLim1NefhhGGAn/2+E/T6o/B0UK0imblA+myD+ioS
cBDAY/E1vXqBYwFeBkfhMSwJN1RTUB6pZOZbnaOiBEIdHAtzlTw5VdKiLm1FKRnc
D8nmt4xfy9W2HBqW3Er4ixyOiKq9jydxohpbSAMz5XBlmLmtQrlPw3Jtgfkltszk
cZdBshuvxgxIVDYBM0jD5sN211VMMrYmw+mZIOIuaSlwWqvwIAizN05TinP30xl6
CzMDzBfcC1WtGT3IJrejThqT/E3lsj7lP3KneGYot4zIw+VKoxVCajZsW8wsBI1I
d5+lr0M3ZvHy6jIXd5FrM/pjw3CVIDtdC+5jakxrfc6Pw328QGNG2R1+br3QtoPJ
o8SZKZbYuJXOBWSj/3Vv0cUYf5NC+7/uDFfjbiVYJEcdf+j149v0ku1GerJaaTE2
MArEJ2WmjE7O1NsYIFwOzGGM4vkqZP3fgB43JqzaSNNTdv4VpgKvAsyyplD5arFT
iNvdcxOigytwi13cXZd/lJOlzi/vf8G8DvVFl7WjxLvdn5npJ45FLAQ5Dow5N+m7
a0myi4dQSBDbR/2UgGEKglm+Xb+xdfVyfAPQmhUXdD41nD5dby4ggSKbqgXYwztJ
QFJXpCHY/og9tN0tyXSHNyFH5gXQSwZoSrSYFTTFEmqhcGaUi6/fPMXiYAvySXA+
UvKvnB864j86oha1ptglMT0lIryuDC6TUbtPh1tuyizpEB7FJSXPxbU7mT+B15R3
7TqLH64h50NYpM0KQGZZiS3A1Rg6y3/U6uWZ+xF9BCh4G5GCpiprnj91yUCqAyB1
b4xZ3gXKOUNMFFQhM8nFzT6MZnYgMhb1PwmP5JNXihToUGDHAWE9lP0SqEQZxjeB
ofiA2oTg6MP5btAX3LZzThZsPv1VkJ2GfgaQ0ZTntXvRNXmqoxJpC1l2+259n+H6
T94JQIlw6lTSi345T4uf9Unc9JkesVMBkHPBYRllCwDgjRJaZPfTN5My/iCa3tMU
1TNYyKc2obvn419ak9Z8jQgvnV1Vp+lCceT2P+7Yy10Lgm+i0bG4hUuxgsr7uNF7
xVkUNnViMCSJHwMT41tbmSlmoFY9EGRGHpqJ+xtTox8Q04xMifBU3hqpjfisOhpA
3gHlpgNO/qHxRgdiwqPLr6q6FesSm2Iv8CsxZEAbcQ2l84RwTSbVO9kl4Xt/tXVx
UAnBvouaDcNuH6/58pPyB0P7awR7npQVoAMc1zoG0zFUn49b4Sh7J+XWQwf7m30c
Z2fhLgN/ehu538gPf3V0D+dE9xSRC3hD4Zco7CgAhQ0DBGh84wTbSGSfueeiU/6y
mm8bTk9dcijus9YKDb9zsfo4+S33GvUDQzpg5IIEqxD14YHgZ7NvukrReVNv8H6I
VfVlVmF/4bkVBltTV5RrZaj84qx4Ey4hLnDAeSiNyCtpWgYzYqBU+QLCbhgzzIZs
pZJ3yRvOqA2/EQPpxewiVJsxtzZpQGnrYrgQeXQ/YEPyVfcLGyDEhKbVPWiYTOyy
9/Z4sdgSUhdfSHTtBgfWqFc2kyeZKrswtpDXrzQ41OGnUCzIeeIJoIdd4HBapcXW
IYe80hIBW6LP2yphPyA5teJJuQYJAYLWW68qTCzF8lJ5JkMT08/rXQrUHlbEicq5
K3VDYP0SuhKCdbnW3eOqcjdzr+jk8XHxgbMvtUM8Ht2aVE1G5unip0rYsl376LEm
ioHHvn0jbk8ISicrihsQPk6E6U16sCJTu/jJh/ZnHnaXfcxF1XvXHZtLgQKBRLys
9IzXfjJVdQ3yOlarmw/caMyRqng+QwW+MdnZ2uGg62xeHQt5nbopb5arhorX70eN
uXjnyvRA6ZDtsQwU2H6gPBPaSYx3DcT5h1RKGw+O3Gx5m4CC263xgZGjgp5q0isD
oVPxhTW/wrjBBl5eIZM2UvHz0VbRFRZnlbOUDb/f9ZiYFWq1B6NtItZC9tO8dGu9
VB6QFb6hR7BeGbbbYx3SZ4lxsUW9L+jFeDIhJn7uC1s2FN+oc9xrOeFQZF4lngMg
CEbMPJC8wvbzSSllJOZSk+fdJv9NuFUnWY5jyPYI/+DQLAigHfVLAb1yPasKSFLO
MUL0dwutF7rNVlqni82b5KHtl064mUeKTGuGu1IYq45aD9ce0ZT6PntxGMfEfukc
xpwVABmHteseBHDOXmIsQi91sMe6/detDL14M67NO+ketffug3FLaRzwIQjH6I0i
FEZv+CR4xRloRQn2H8DsDZguKzcVVPoF4lEgsxIr+iJ9JtTJyoWphlqPtvTZN3/q
4TVlQulFt1gOc0AA77YgQCKGOJ7yWmLMYXJM6A+Rx2TqDPbGS8XkSeR5DJzNw6N7
qXXxLHEy2O0OSKhQdHAjOsxlGfJb7BdEtKhdx0dxL9ESzgEd2GogOTc0KUFIYj01
aJigNKcBRjLeEdjuds6Ot59O+NfBaL0X1YgKvrVID8Sl9LVEzOYpzCswuL8U98Q5
zITJb4lHpZhaL1QBO22J+ZsN+tpdnmq8V9l+ByzV2srDMcVBNrRbn6l5UeARrTqC
gktUPmz+8E1kvRDkwiWSnerFB3eVcpZHqvzX3Rp3f1jJdCUid37h7SULfq6i01H1
er2CskTbO8yOMOqmeECSOzdFAipkRlx9VcRLsKFaqJRnj0Y36KocSZrzpm3C4tgh
7S7SjoYrMbI9LO+zSI9UvdBVFotSviPDVfcw7GvOOJ6s3AQ6tsYBonre3ZNFHjEb
Uf/jGTCxpbcDcjC13kflu8ZmnAXJzNvhgTDCqgNfuc5w7Oyn/Frhpo7I/Ky3W33G
+X/4zjQI4BEfa1iwwtFLnli8L/L4ichDV3CPiwlXU/R3Z4ndNmyP9Vp0WrtvL1T+
USsibmfUDV5zOv8iVODjdGYASDAJAosstwtNRgt7/UKySmp9ZcGM9l8dPGGZ1jZ+
TwOr57F1SbV5HFiLmZV+e7hFPLERNcg2CC4wgMaa3nejwUQyHBB6UDpmb7/22Mr+
4I8RmyBSKu7tES56b0HKYvmsWdSApXFZZb7e5v8qk8uUxyVI/vPXpxsXSZbHxEbf
rONfBAha9VBFOCobXxnIFAzeML6TsAN3Ykjl8p1juX4DwfeOPwY31m4dqovuiWQK
ymrwxVYE8KDWcBWm4/l4XBKaVk81qkCMx6wmkQKX7KdI85sFEvP15/HKVo1e7KpW
0MqoO8q0E1pCEmQ0oL4ruV5Y45jdoAPf5Y+aCDCaLq3dYMbqCUJA4lO98cE2/5Q9
MvO2onGAoCTlgIAxLR2V1O7uGvlhGF+4cMIJKKGscfYwFJfbN85XvRaUiKsudTzi
MaOCcOBM1Fx37avk60KoLc+vwdM7ETYUvnkiM4VpWP6fFrLeg0X2/SY3VnCE9dXI
ixagQRAWfP0heuxzlOwXtIUmkFYmEsLbg9K0Edatt7wOuAyFVRsTWvbn26/e5fAS
7aNgtAdeaJot9X95EvYYl+hL0AmsfqX7c8MlvCQMVEJqGdXgc3EBoIz5FuYCQ4pb
TyI1T1K3CsRLrCU8l2fcNIf38bVt5Zti0ztKbk7nyJiC9aiT1eMinCiN8pyf4HGm
KBaAWWHd+57LPEupnVGUm7f7VIuQnnDIkB7zYRqS/yvqIBcmQ4wjsoC+IJe8GAHQ
W8xNT/B/InCIRncDx8EHefc6eba8Ibyi0pfXrHA9+2tmP5a0RUFIhdmmAs5LPxBI
gFYx/YA5ta2ErvSa04tc8O4ME3QrqDxszuONy8XUaHBvhe9UfXnJY3UPBHuiLjPh
y6FbP8vfmP7TY/4qdDgyo0OQkG6MFcr4DBFsdHKMtjgLKn3IYhHlwOxn9OsbBP0f
9TkEjtKeRzIKwejTfHZo/3BiQQ+QctctLjJpYs7Ijl2bRY4pkFGYSA4P8PPEfw3o
fqXcmUbUtW+BNus4W++3bK9G+gxGXDBZxEAJopemCwanjWJ1e9LfYLOQR6kby3cz
i7ZUoxdtBBgMSIau1R9MUZw3teF/UwfdLK5yeD0HSWvyvHd3wxxGjbReg4gYgpEn
RqbRdOxNh9Tbq0B9EkrcJ4cR2DeYFUBRsljRlV+7ZyThJkVT5cVaKkAOgelqLCpU
8V4KTbRAzUaQR74EzrPZur+8KBTXNS0G+9ePsipXjUWX9LH5z1MAPYPXB0C80HSK
nu8u/m3ZKt/IpE+BDqZFa8eDwjk6P+niT6/bgHGZzSGwsNkkDL3QDPI4vwdm3U7g
Kuk/Q8S5DmY8EaxHXmFBgABPnq+RkU1QkoUcWmAlOIx5VEIdykYQAPGdPc4IkOVW
WLj1l17CPthpjYzABZRyFJdmRU74trXqY1MH8hyRW2hoWuI/2M/ab6j28Dr6psxs
21sDQOGhmoYsOx/9eulNmjFwTdqxEW3Cl983vKBlSz14fnue2TU0FYNsIbYGYHKw
liXHLx8jtkYBDALK5zmsOLy1A29SxPrslVq4EpnDPv9cS1LZ+E88BJj78GkCvlcJ
LkRMNcFzMkGowqXlLii9Y/ySZkKk0iuU29D2hNXbZ+MrKlsEK2jiQl5RxBh0zFCI
xa37Lh16eNGLJPpwli8L4xBrxQmzQ3zZWQqtTRLpXx1tM6b+DTXIvIaEikixsh/N
fgXC/27wbMTrUbe37k9/1AlTkkxty01oc/9dmiissPHDGMptlaxOxdAULtcgn86v
0z4YcJmPlpKHWRqw8ApJlS/rrhCc+0ORV4QLD03OVM3ob9JxqsMXuTs9AZ2tYPf1
jt+BWEVJMzWzFe7kMGSEjBKedYkwbo2dku9huTF/LEPrisLyDEQKGsReNY0GlTew
KnAf4Yzobq9LfNdYi5QLcJsqWhfMfFf0fHWNlZd6PLoXUKQYMqD1k/Tu0h1fmS8w
XDBZiji9GxK3467/46rl2VEW863s/apz7kB49PQA7yEyXS/CcVX6J/++PoKOcurI
phcmbUbSzK3ZKrEDr3hdNnx2G4RK/7uSvoZFmHGzFRlH74zmS0II+w3f3rBns2v3
p4tu3kx569hVZyw6zxzN7VoEusQlAHtZyLQMNUHy8/D9AahpwgP2MeqdIeXiKUeV
NXk5x2nb9JEg456hVUPXjUOF7STsjexa+CKOVr+i2rOBbWwBJSoJuT7DwL8JVC90
QH1LtcGZpx1QOmtwIaEt/raZCzVERaeg3q0nzKZAYkU7TDID8zceHY1aOCFIg7Ly
nkS5dH6KTvpf+hq8ongKXPoyhHK6N9AhngY+Qdbk7dDfIMgvP9xqc6hpfrweZgrO
8JAWNw+w9VtAF/M4t77vQ43fGf3yP3vg6lZwR9M8RxBDaq5ArWJQIvqGwS+ziWhY
K36IKUAanR/coAeipLjj3eYT9yKTVnN8guyvOfJHW98rbJVH2sYmVnvXOeIjJRuO
MNoPYlwxlYgc/gZcvWVcYdVRi68i7xzMsnUWRWGBr9eJoRxpkgekLVJ38KQU87kf
5qDtqMfiaL3B3e5646yQ+Gd5Hm4CZgH8YcvpoBIARCQRmgs7BwJCLqcloPw1IdBL
kKwTLBm2LRSrXmskgGziDKBQQQ4p2Zc834BVijL3WXVs/Vtx2bLWRnpxV9ijZZ0U
FWsvPM4/T+TozERTKY3CJ/JNDLjqpDlsqyUdK0bj/MuiJ9GhjGBXoG4e8giXQz1v
kLgGdf/Oy5watSZYHrqsK4X9aiPOpeSOxXyb628+6GWp760TuDAi+GcI4A0lWRnD
ZH9lCXbUOYHEyrlecQzOYsk3SzHvG8cnpnSe0BwpBQLNmUV8Nb9oeq4D5GAvzBGh
ouw/MmgxlTsUE6v3lm7GlDAridtAzWW9vBLtOth66Sr0obMUqDDB3RqAflEGsMoJ
gaES+W6784BqgAN0lqtKjOSWn7s7I2PbwQ7pm6KTwqKUgg1VnkNNrybjwSTcqMLJ
o4U+ILSS4KY14qhHPLPP3jV/zC344l/H3i6bZkKpFFSRvc3hxWNuBpadI2MWZ7x3
/P1E0rc/CDASHQbFPTLan+haUvtlhUBAwNWEajuK0TLU5rcrfX4chwMSC2AHr1RY
wabMR6c65vg9wCxx5J59ibVDlKsZEfW4RNirUVoOZCaWhr+UAVjutSW/LL1keEg3
ri+as2zfrYOtdjghQQw/uCMtDZ7lQFSCwSuqLPCGJZ17FM0zZdUrdOZncwBQgww6
rjxV0hh72gpKevfZtka5RaNlZSoqtEiktTqRVvnuZG+m2cvm4MFsZHqEJ+DaqreH
cXv/mA75zjy6AnyFUuJl3DfmO+iyf/9JtRxyEG2u/33YnPLNWXLVtw2Zv+SY5F72
Ar2zfjO1QMiJZeYXHK01RbHYRwHQGKr5yMveW0U6cqinRSyQbUN3YHCc04zEkS0i
VMuNu1ubMqbgJH0C8RK0QJyrmWJKs3am8Wq4bfj5gsq4Aic7rxqNem58Yc3IVN2d
++5bG0fqNygeM+JPuV6QcD4zGZv3LwXFjVsZt3vZzY3kAGJYmSYA0VKR7xwdqNKI
80AGKMzwCCJFcy8+d5NUNopROOPKLq9ktr/dasiVnazQcp6VwFAdF+DCZE6WQFFN
2GDNz6eGKA7NtzvCEZPvzivl08QYsUMVP/egTCen7oPwA/uMhpHBMDXinLVLXYMl
97Qam2a+bK+xzClLaJ0UJeYZSIzLZT3u9viOFl3YSPu9ofkVqzpl+wcY3mw0v5CR
HISa0yT/yzl2XGmV2eoTOwG2IUSh1k5uFEMuDvoBvCslKe/tp2c/Woe9Pyc9oUoz
jF6WJb2MyrG4DiFVD1dRoTptnINUAkA6ittfqIJtK5LHna7eMgNOPShinfjwkcxI
EJFopYXFYwV5Q59PIwVszNtB3jBYLVLwt7oTXx6bcRifYZQJ9O4DeebYCV6mRdUp
70r0QOyoipdoxLmbCmWzEk4oIyfPNMdtWrM2xIayA1BTjynIecZ7N45Sp0awC99p
EVjTRG9lmvxine6zsdAIT+nuAt/7DS/N5YhxN45DA+81N83kIdkFy3gsrfSTeXv4
iHX79qV+N9U77lEFjPMXnJ+PJAO02Pna1/Sv+LOK9uExwdrM/YhBFVC4zkjiN9dU
vmM1DrUYMqD0//hWMG5BP4VwzmvdxlM9URiaCXEJk8b4l1yao8NFhFKTfYNJ2eQh
gVPFLYMO/N4hQNUzmi5Sqtl6K0hLpOowGz2e/+G0tUHV6TxsLA/o0yjUv8yYsZPX
Xds47tNLfaTM9ZMLOurkVd1xNeSUhVXiFZ4+HcBWWz4nWagtS+vuSPXslvtTp7Cf
JtGxB7tF4LNczh5ZXXIE+Ttk5mqpmhyn0faFB40xnjTRMKS30UbXd04LipvC64xd
3mkomK5LXgemRqbcmJTNoPmHVa63t8obwx+3L9MOlXuNQC3m8mI6SOt5gtf9Q6fS
DBHTsEVBmwKnx1JC6xTXsHKZGuTEUx45m+GHDYoJch/KgKwIp0oxEqKxNHAAMERH
cDhD8BjkDRi5082RMKWDDve03Pxl/hbyiueqKtXwDxJPEPoikHmNjp3KT5FeZjNU
gd8GmEFbqLxOPGT0gmfKZZkl7nQr26hIE9gdzM45ZGe9tK6RDbqS/qOVjsoBsOZs
4J+cBQsaK/tK1v/VdmzGsN+hlLxTzJpcwyzTpaZ7cMNTyd3O0f2h2jJbFR8amhbc
EenQqsH2DykKv5U+y9tSJ+ca5Nf/sqlE0P0/+ZWjJcH0PBfsfXFl39+He9ekI6bn
NPYeCs2uPO7LleOD4O/A9ns4dnldMSqVQ5GgE7XLyvxlVW1626LnB7nGwMRPk8Jg
4FFU0AapQpvIC+OWBMnumqHsLhM1fl8ZAKFiSoY+Bnr9bQzKijmui7uEIXMWjjok
1TKrgSjRZi6u6kx22WSnsPZCX0BGlegl94qm8tKiWe0t2aGCDcnph3w6h2/Dfn7P
kcB3N7JpP5yQv8vOrMAd5LyeU5n6LG9Awf26VIrieMckcKHr4dvjmAEkeV1HN6jj
GZmD+R20LmXVI2l74DZFgsXdniJVOPv/Evvx2N8P+4O2fHw7L3N9UQTMuvXyvYpi
zIOghiQZloNqmiHS5G8bY80FgAFqhGRj5Iv2BsFY+ILA09JpFbcYS/tS9gaz2y3z
Dg7MjrX+q5mK00ZvBdodpSyNjXtzu6cGvuICW8ilWQfhQAPuYxqjcY7KQJ2gCLx8
+moFjiVTWZGSJLcqDkXTaIy0VQAgHw749YduF3lO28WRDp+PwVsMzeR0GPsaI2cN
yYoUCGuZREqPAumTa99okISX9NRPSCrFyl9t3FFD2KnFh4YVL8hcuh+F1P4wROG7
qdP/YefWgDlfYok7ay/1nn8I71Z2QMAXEPK7dJU/bcGd94mu1o7Ft4OA+xNi8g+M
MyohmvOwqgGEbdtfwWvTUOlYhr95FgpHbpadFKEqjchB1oqdXff1owbgQ/QmXB6r
f9IstPjCScZaTlHgPTcRONHGZenC6eVwVWxkglTpQciN0XO9q8v7HslM7d2zBZjb
w1N5sil3y1rkJ1TdTIxSTotcumQ4vzdSY/f/YTp5m5y61lvbN9Ett6XbMDZCsnLG
/yzFnuDAw4dIq6+UngdQkeWEWEZDlx9htpXD5L4bhCv9GHB8W70HJk7gTOg8ObSR
X0VW5fDcqONnrw77J12eB2V0tD1nhmK9FcX6RoiXY9G3HgNZDm+UUaQNTyZVea7Q
J53X2USNC3O9Yr5rNul4t46vUH3xfAzPLJeLQMeH9xK6ZK3rErCGz1PEpoqhbGDY
vi4zytwY/oREpgWJlhNWXjL0ArmCcgzhkpOJHxn231+qB4j7BZLN7KdgAP9J6IST
L2jis+peSiog0ID5WBz2RUKKLu86Uf7286mA3Veh7Qun1Jw72vYJGOM+wf8XuEXu
NmzJNkAR2kCage+9aTt7C7lOxxgBj5/MBI5/jthCzUR56tKxoNf5rmqhNOycsuaU
7a30Qg+q18MPiO/rvpzXA9eZtUAlKrjdVW7yvCLLcq0+qJY2NJgp9rSqpz+68+nA
h1Po0U7fJqunOtmFfIz4YdwpTxd3VcgO1VW0okB249W07k/JDXWSvg7OcdK5OVH4
aiV/LJvqINda80k5RF4KaESf7CvLitzG4qU2/WApE8x26OBgHUQPCCu1MvU9RaRe
NdUMFvDtUuNmE8Lbkd06LVZQ4CKCb4zE0yRc4X+rQAZfA2NEuXGthsa1t3vIU2Dv
Tt6A8qrVWSjRyNloGDeJ6EIcJ+SXI3Y/dmnbN0bsoT3of+29YxVltCrKHsONHESt
3qeFBccU0LJQGCjdog0/mz0g4eShuxg9lFMxzjdXiu3R31fg7XPr6IIkDN2S4szh
aYys810kXtiAFG/2AONf3Coejq2O9rdCdeSmirsysFmYDY7Ht+sveNQLyeBfksgu
4JXaewKlRAEqo4laxmtCPnnkNZepKLSxuFyk639w4lovb0QcXW3gHwDAganTi0Ch
e4l1W6xUXzpE6eI396foEUmMx732oSRFxXedKHmPclbQeH7qL8lU4qNgKMbMZW2W
1OgDE2AJAhh1s0Xr+4Ro8jSTx/OsFlRgMh3fNmq6w/3oWSj7CPsctpOP6Ce8CjjP
zkf+o+4ltBvh2VrPUK9uUtaaAVeJ4u+OAy0uO3ORmNQ5TJ+YTP5LNHKuC1BUyhV3
xNbksFWdNV+n6A52/dJ8iB8gVNAYpnRJRvS1Sd28OyaL3mrvh9C1W4VwWMYz3c2g
Xw5RRDp2PGhtFJblNGW7/lEktnotuCSYFdyGyY36EezszPVTmbrRUlbB8lvrdDRm
a54ZV0qszW9biqkARMr3o6HKqbhJmysGIICh3/kJxE5ZmW6KFVuTJxaPWN7M3VCq
im3h5mQmCcU9u+jAS85nmH6SjE9gqkxAXQG4/3Dxaa2bdRsMPNI0mJ5b+nGEES86
TM8WyztMak0fvJZwxTYqrhpntpNjaHCeq+Yp1diGFB/s4kF5R1yHoVjBWVp34Rnt
oq+N+fsS6GSn7UVQwuolGKYUxSZ4sF9sq2VkMh9NgZgn6gpB0H1BrRrS/nECslYh
aCwDtZFRRl6ZhQHlCiA0C0p6W8HSEMaNU8N1gvceO8IGyq/SQ9ah3yF2acG0pQ0Z
eLKx+QiNZZXwb3JsoH29m6eG7H4TX0wgSr7ferKtgKWxSMNxWp9/zNhsZse7pEUk
lY6PokNRN3jneHfBqYq33qBtU7ICcCB5XVngQZJ2vo/4A0nIFMomrNRlZhN9UBoK
AdeXVbg5QDQaL7SeOIuOeiAzcj1w9OwT/1Fd/TinOGN35tKRna4WgA0twQhY/NOn
URWyqrdClpdz7GCb2YtzcmQzQOFVZwTDIS5RvuhBC/oxqPHWMaAEX7Eiu1WgSn+5
u3t4aSW6JDximuMMpybKSC2ZyYCBWZxWMAT3VW78FQG2O7LwW9FA1zQVetxUNVdP
FYI5qVAWObH0Nd7DZlss0uaJcLFhYofLSj+gRyKDyxGDBDBCG+99cLg5v/WVRXTT
4l46ckJz2h0KEHNT4pJbV2JfRD4SHY5e1lfBCPeCawVJT7HU4dd6Ohr4se/+lXy9
Dn6caw+COCGPHCEl2UP1lNd/p0VXccOzJgJVb+dAlO2QDdl3d2lFvyEcwFhh1Cyq
YoyraY/av/8InEZTB0IT6caI76s6+ZrU1bHUkwSGUcKG84P59ynldM9jQrbud3ZA
Lbp4Zxm6c0+9YH9sNoRXS0j49acWd+mB/voon/bV1SsWvqvvGUsQyXu4BFXM2qvt
2NO3lE3ygWiClHdtuCb6GfQMqqyvPiQSW0luWPoepLab5e4xU8z4HudiDCLTSJFO
QVFWd1kvk9a8Te3/HyME0DxLAiLLQSY2N0PVINPtrxKpV2yeVNpF0TyThsKcbJkp
TNFHgQNc27Sr9Pn42OpSPJGPh9UWPA1fr1+skha19xJfVDUbkKDaLyi8pbC7N1Un
nc6lM8ndURZ+9SBcMDGNCfq+eyg2Y2KOAq4IcXACMLF5as+RwdfCBwdHnPSYWGVL
cumCysIC0lKgWL+W8UVbDwpnRMsUsVIg6WXCuZOJFiklWG7M7wxwZVxyCVrA+1q/
k8gxQwVZJF8jHVSbg5jHR9UoNbJTutWOGChmVRCHXuDxrPqeCk8f/stH5uIg8xfY
GANDGOUFziAE5cHcqTHLNcUazmz1HdsWJVcG2/9cevRTHbHURRCzYYDqfLHNGxZP
c+kF+vGQwHxrOsHfpn5J+v37Sp3MQxjD0/uTYl/1s8Ww+GJAw4wuwj5Zldz6KquF
11rcSgPmhe7a2F32fetRGM3kFCGFTnKTmkbt4Z9N5leIli0Ef2V4tIUE0UWTna+o
VYLbPq/BC8QoXzv/wzJQ61neAUyqLKXK0Yd+vjbuoGzPAhVD2FsjtfJf/6noszKV
k5psGu4wLrDuKHyHenHquy9tDgg9wVuvZyfi4AT++AM0KW1gSgi93BvQlSEum9dV
5p13uUvefatLXbNlhG2BjfJvsjSMgPeD6Nk2lC/Lw39CkWhgHn1j6YspsNVlOi5x
CxthrDAHbA6raoqY+1Y1W0sF6uH84ECWsDU0sUc+Qop2EU97WFfzLc2HftPi90T4
WW+8ApPHU/3VL5aCdHyHrzYgjj0GwmNK4HFB3h7IHki5tVfS9R63Ez5dxXX8HJr7
f7cIVdjUjzMolWPl0NYgT4SLs9u2wYAlJXikQ6mIDTNI1uwgzvGk5NhqOq+Jz1/C
sSTkbA6I8W58Xup+BO/jpRUiSncBW0XI0ApI1AKg8Iitb4YJgmw+6VMkiSGSsxxd
oHY05A8bfspHAcGVDjdLesIDgxT6GhRKeV9K8Dxnbrfm7/8Q0k61aCxBzKVwyTF8
mgDhkppvg/cNL/FA0xQfDDZb1wo7FMhNR1b2HUlUiGf96SzPU9+eOTa+P0+xlsea
sZ9mvhagIDv95LYUA2plIv7MKIigDHMbI5MpbcOYW2/qu0woFS8YQkIMd6BWLEzO
AJPzM4YWxkMCcqfQpNagU3HHzaFGS4NFecw9fTNs4ljDROYScYvGHz4ei7gGlNsk
qicRqkG7qZkB0ESxltU0hMJOrjL3UhdgyJyVR8KG7//0Yi/vWS2qQqmH7uRzb6uC
7k7d5LmOPWPFtt6CPc1qzbfM5lBLZtDMNwjsumBnKbJnFRsdSFaA7iQojsa1pj3q
wwFc/jXidbTaQfyBiPupb/H2oytgiRhMSyYV9+p/FHgwwaQigL1gr0SYRdQNUuZv
5Bwl78RDannTLao5xkTEjjxBKJw4M9JDZeO8H4zFsaMqRq5y6s4gsgb+5cZN/Kqs
wsSvBv/iIM5KnYhKGXJo7PGKIKDjjjPU2L5I0PV4hsRI8lpJqIZrHmNZ937t2Yhg
rLX8LioEsqi0lmm1O4Pww1B8/5fN2ns2ZvD1HocWayL1vtU53i+SeqJg4g1KJ7er
SdeuVlfUbPXhfsj9Ox//8ne7zxjFu1rUGoLG28urOluyW6VGVD7VofaaZ5sbFtlx
XFYIwzLbOuUzZCI7o5HqzC1BSIyG/yTXis1IdcF8TlQrpf4QPY3wqsmec5CZgeIX
h4JnfjfWZ6xhoQ+AHNrZpi4dvdzE4paicgB+Rz8ZYZyQkqhGpgQ60FXhLXsbQ9jH
KTD+7hvNgebfi2DXqSocw1LMFnKBEHSwNVOCo1vndl//z0T4TBQceuQze9R+PRWB
dpMrvhb9aok3xmI+Y1AZMBsQNplrkvmNxEiHytxhoQrFyTr7ODaMLmngiEPeg0px
Rf1kEvNwtHYcQyZtSR8DnpDt7YAtWVJaeb5hwQ3aYBru6tUJtwWcqrfvGaRUsrg1
y9zPpSKWCTqW4843In+dIuNOT5q9SahYL06w+QhbGMeFNkoPZRBxQgmZpsfOXcXv
4joM7xbm7/kQd2l/Ae2L9fys6CSo7RqWNYZ7SOjMAYMW6Qo7rLyoGpPIlhKryIAo
K0OHA3bkb3vuUfDcAf1FJnpDwJcCmDR6rKi9BvLgtlKLCL2qg1ZzcNsyaSU0yRLR
xIISweraXScUoiQa/NCs/A/5pyfOycENw+0IHUBLdIcuc61G3/hVELcs7xLKX9/b
E9tlqPpr+tZcHLcT62l+umcqCp+kJbuxXFpV7gJGZ77YzBfZnK98GiC4OdBpZM3B
Bg38UFN/30LBpqzrwUlxPbLCdhrH3W6td37qxZDCYWWHKXMnT2HtgQnz+h1Hwz7Q
/AdlKnKn4SPtUj/DvkoMjDoxmPE44UPfrbffmkl172gtcFAoxzGnca7KwemjUn+j
iO0xJOQg1JwWuDeMAYVNz7I1hvrNcpftP8r/KDZ14Y7+batRdAJlBQwVwJ0j5cln
qIp//ZURThzVopWH6EuStUo4fsJR/n04A6L9SeyLWh6hVltt8DIDlTiQtSdgy7sl
zTBxMUyk+ZDgxFypm4hFF74wsjIee+i4+XG+inWSdwd8EDuI9dYCBE6ONZwM6TOA
iQUsbQt+yu2IGIs7YPriDPPKhBSigsmLIrLGd4l8NAOlvBvVYr68jk97EFXBmCA2
fIke+g4+PWe7ifXNJP2t0xgr1su18lcK/UiTwAo+rLayP3fmQMTc6dG9643ujKUu
Cgy2ayVmE0Ff+yRJj02/So3SznQpCW6iugfGEVeuWZ1ngCy79V6zbcbD1RDeraLJ
wJac4qhZGrV0VGgFT0mVJF8S7eRuuINC//uF28trflrQCevkS8C8qocG5eEUyliV
UBaiPDAeG87Rb0UId6noEJuDaJpnSTf5pU5hExjyB1aQ+gBkjdUqAm9hQZX4waow
SJzEzV9tytUS+B9eD9kCMxJpiZjMzYA14e3hiBe2xetYQJrrqIdR1k4oWzn929/m
FWwm7o6XGkmPKN/0U80GpZE8P9nfTlWHvQ07+cBwQ6MgnzU4C2fBHvW1QEiJFpoL
P5DZb5uJWDjKbEE9JZRUG3fwMvNVP6k3ojgYTMNP5CSC2RY+MGLANn40aDbdAyY4
3BlD8fTUqoaePmUn3ezK/jO0xCI+i9dcQCJZ8btVylxEki6G9eHR6+PKoUyyo5FG
8sOIAp6LtlBpX2HcvaNYkOi+y/k5Bg+yUhv+ISoyuH6icW1B5Vq3GLowULkqD8p7
5xVWx7k/lJwEMILpenpi5y7N8lsKstUKn45YzH8yv+LR9ZSvItJXSwEoMJnDQpCI
gcSimCMxoAkxeetL75HLg7e9MN8/nsOYInB1j5Li2Efui9AIg4AaDnOZ94aUAqN0
1mWYptU9kJ25Ryf4mmp4CuOKfuueBujGI/0w9FrDUq/pKfZgg+12e71xrhU2rBeP
Q5dzS0zfeW8+EOUXAOwKm/pnZF/Xeu8bR3Pdg1pKxyoJy+9x9u08WaC3jxwPJAoV
xEq5UaT8FGzKuvIpsAatzBfGXa8b8900WNHhbLqaMk1VuU+ta4A89TMZTeQAo184
hYQb4q1HGxukX7czplExECAhSS9jGrV9Qssewjbj51VDbEpctF4dYExp+5xyEC55
DCdHfTDxZwXAT+Oj9WKjIc1pVEJVkZYFjSBA+M+p8qIzWAgRYU0lauBtgPn64QsI
4/BL3ib88JN9QUI9sl+mxm2UCs5PZFMGCI94wGcSiKbCOVa6WaEsec3Ew7UonMul
6i9HuSsRI3vzVrOfUgdxejjRrFQg4oFGaIFcfh1yYH8kQ8Wy/Jn6pMDpyzyqbugY
k9jeHtJWVtXpEpizFkdlMm7nGx+eZk7c2eW+k2mjmff8m2zEMuYbpca00WlHvbcE
1xinSaITn/kNFhMaHnTCypUBDhON0IccY73LaMh/uW4uPiLrp5MGd8qEdyeZX5U6
fXD3rl1J2knOT8xZ3gGSeMcel26YTKXaATLaHQtH9/F9QxcwL2f1UXdJzzteWbEX
zF+vvNzxprVzBhe+s+NvDgH6InVtumo9I3caCwSaEmMRZhE/c/am39CrI/ivGuL4
HhOBNB67spqPCeIS1a5QfZWbupq3JQWky6k6W8OxnErzAkF69V4/kWgj58aLxRl9
5uNTZhddrOmL3u8VRPnerZIUzvRaOZzV+QH6hqNbNbT8A6XpgrIOXapRAdLF/2LK
ZnOdFUEeYPRmI6BQ9qz0cJcCjtGCHyTIfG2D3yOojZNj0Wnv0lv4Lwukv9DNpV1z
pL//yCcBwGAyYQ1BVCD6NNSMzaEFA6Z8pPOYSRZs+x9eTwKkQZunSZ2bGCYqEpTj
57VeWwHH/BzyJR3oSKdizt1xL6IrtmvSrofiPFC0bjVXjM42fGyZZEXMFhcSJ3Y0
syMqtUjZdOOqWVAVNxbQ0J3xayad1OE0fW/6PpJp8XRGqOkS/Og1QilEGTqBtsBu
+zUMeWYDlkdWeFL6MV1I0stCSTsnIHY1Tmp7WbZ8ywj2S4gA9njrHUycxGtBgf0a
Tkr3XKMpHHKQc+JCAt0spp1dMlsT49ZDcmrUl1OzxdVuoJFxxRThKCb/m67O7ox9
zsuUtfOd2c4SUhNTUlIi5Q6XSxXJ55iSbnKQr8S5ZcnepuDx18bRqdEHyOsbInFZ
IHA0txyz5eHpZaSxGcBWNCQCUFfCQVIfXUaYOAr+GHme4HtFfcosK+qW4hgS6+o/
Ieo7TytMLfmSGRgUOIJqAH/hxa/Ie3ksjXN+PiPuRGcPJxZoPXzAeYNq2JvhRO3S
0Q1OP00b2LI1dd5S5wY4Vd5/Q5EufpLNzfgUY+wnY7RapYXYtig9DjbmrSsgTndk
A7MttVrBZfBSlQDRLEQ9MN8/7yc+/eKVFrO1Fbp1eo5yLsfJDMgNIwic02wUHbac
tYkHHTIwEv2k/vFDztV62orjAsak692jfrHb73Sgzhn5j2EnFyyutDsq/yU/59LK
QJzZW0cJ6mADaFqAXipTgHWHJPskJQvFWjfcOsCrqF5YsORziRgh0K11qWE/2wZ9
7NvUg18qNJ+LCLPmjwdUF+z/BxJlZsRftLAggUb3jdcyzUoXvi9KTIbcsgtHKXER
tLl94cxID0HEQDadqk3Q7oI0ELrhIEsFkjU6aAavV2hTgcLEMudwKeaOeP3Jr/ff
G4+MI08MMbWZ4s6yzWpLBWMrNZDwB4hviSMIp5mgUTXkkENmv0+4L+gK3mpAyqhv
asytwIT/Xeadw8g6bo59BcoxKhvn/PzdcXzdB8QV1dBhAu3zV71oiRecr2zKNR3p
p0I9UTsaGYVN2XKf8xJI6/wyxvZ/oeC491cSUlkVH/s8HttrR4gVv7QV0aw3jMIB
9OY0xmFKv2Us0pzeq9pyTnAbqJPaxN/CF9kxK/2sVOAjNimlEWBp+69xYojfw+VN
Im9Asf1hwKbq+/IvtSzXr0WNPzwtY5L51ripMd2VvvUdvpwxKETP4RS512DK8S/x
QJY/ytesclvTV0Qd9OgEc97IoScKzFacsMQuoQ0NyB6wAO7UolJUKR3bIKwUM812
9SFjgukv8XLfhbIu4ukHLnnDHiVB0HZh33JJzbvCNEc8fVDw8P5rt29xDSK7IGrh
uks/RHGMEO40cCTRf5b7VMF5ZecL4EVtPOoJz2m+/ayWCoh09AAHPwF1J+bAe+z4
4LHRMQvPFJ1EibO0hMdf+Uq+JWyBbA15GMIFuDEwLbXdFzgtMkdWCfX6jfBXabsy
1FU3utwUDDthmd3CiXSdLG8HGmSp8GStNraKvbQtGtQSLEkeqU7Mp2ar2nWltBJM
ytKtrDbr5h6fzk1VZ1Khb14u5mzpP+4wu3QabBRCzeBcbZIMyBe+UJ2vSwnTcgpu
d4aMqytA3mcXxZTt/Vv8v2B0PzYN78cpnAc7LFwd/vt+ypJGGY3cQJs9fKTrfLVc
cawLu8YPS7iyWm2bqNsjIKTrxffGoed9wNe6u4laC/jxiHbTqKT3ThYCEvdqs/SJ
NMpXvxFOgQBcpg2Of6hrPZCqSO0naqt59lzxyGcdWrAWT1OJOCfZ5nscnLdzxNaE
dnVNWktdumVKGy8yVCsSA3xw2gGkOhGH/ehggd0Uo2gMnmZ8SQcPA1yUTk7NMwgF
ZvVvQkM8bsoDYn2Gvc3iON/K4e+756xFsjAu++P6Zcb6m2Z3p9cRvwumtlkFujJj
C3Du+coSEy9XT8KJQBV0VBwdWQdr2U4bVzvzEvVVE44yn+NpF/0P2502s9dvWkHg
/sFzqtz+9G8dc+7Za9fLRgky5qK/AN9QYE1L9s6A85I09uSkT5f2X3PHU4JaBddG
2E3pQef0Z637NFB02L973IGcHhtaHDtbyv4j5ByunTaDoXReUhbSx+gyJZV+ejAo
pyHBJ+mZF7msvhFblY8vp4UFQHGx7/3qnt0nG+YYjGLl7tLx2Ns3jpIp6WHjFX/n
Fn7qUjsP5BqXuC7SavDHFtC46ppX4S9ndoSQNsmduSXiYlWGKiqimuC92BTNkgfe
j3RLEG2p1nW8jwbq9UHYq3PsZl1xOj5eQLtjN75DFx+3MpT28h1a5+8ykTUJekeK
URMk33WjharkljfcdktZwsNwJrg/gblKfT5SmsmyZJ6MT/oqFhjNcXvnOeNCTmJE
LrWFOl/gVKRK60NNCcRbsZ786pT4AOhhSECOpSbxK++GIZIbx2kLoV/z8a0LyvlX
aMz2DO8W3e9P8/OfN5QlSkGbo0i4VbavwPLdJHISYfPkSs5MhAWBgFdVS7Ya7QD1
hbENEpQKMGBe+QzNRIkS8Nhoz/1ZRoJvy5tgpOhvWDy4/Apg6n+aH0ec66CiznIp
Ml9aRnspDAf3BIYHxOPHMbI+EIJfxHvahSBqOO+w8QMDO7HsawVTk/icQrMoStKI
SCQ9bC/5dnezV5z2IirRZMrooe3vW2Gws8Qr0ozyITJ3suzdhMYNHe67lM02G9Dm
ujfffBo6+TGH7KLj4Xe+g/n1NBUV2eams0L7LFD3CQww9rAbQrqUErCUQzyCzdkX
N9foig44PZg+MS/IrVo77RLGLdLejwvdLPjFu7yPI4cubONV/lIlTtw9Aq2l+Kn1
hZRKQOUxlZG01Xp2KI/D7K2KncV++W3Kht98pUCSEs51TwOjWxzdC12uBBkvfzgG
jg9s/ME9yekN9/Mok8N7EHipHDFrbWvr4SgcBn6w694+nsdAxktGq1x45Ml3DvF3
0PpAlnJ+BCGPfjB6U3XQ01rNnEe08k5AHq2Degj9WUM9kIJD/ajFBMEjr0y4c/iC
eYRL6bNIsxUOSBu1wuLtXbA2n0gDy0S+xz68F+XZY3Z7EeSgJWPaVD0uCBINyt2m
2YaJSgSfgIk6ZBg6cCRTj67YVTIkGsBlzmKXz5qeJQqyDROQZWtQZ1pfvYJT23e6
kKlxg9v/Cck0TIauPqNTRdC86qAbNo28lAOpjdcN85wv0gaClEeQU9jJ0FGvBpvg
y6YYY6cJFplEEfUPEZYhwrQdhj2gRAA3wb7XvvD+W9DQ3BSUXGEnxkbOqIyHWM1M
z+/mjjn+RngOGdVBfm5jrQCBOqWWI5WDbdnx3jXdsCWORI/jFDqmOacZXvVso5eS
8glER4V07HeWXN0IaEOSjpsBlKQDn1B7GLvXrIA6+mEiXlp/beOBHup3GLN28B86
wdRbCZeX9LAdUz0UDjzqA/aI5txoUzmq0nARDcFqN64+aWSLUeRyULo8G3p1rgV6
VxaEbl+mT0LS8fmKMCtawhsjObVTJV2sZT/XZOmKn1vE1ITTnqHbZZ60TC/tb5Df
/9RsM15OqQJ8TBv+aH/yhJHHYKMDy4+59myiQ03pfJc54c277Znf7HI+xKvuFYGi
1GvGXm6lVcOxExz86bWs7IGcwlZi/v6LCkinYerg1C2tWV/+h1+L+3HdPXKa0BuJ
iGucGjw63UoOapUvqDj9IU6GrkX9g/r3fas50gNxbEX69Z/KL1rOuTBtUvQv92w9
b8CL4MOK4QHyw2z++gs/i5qdkwAcB+BDuxZ9HqsjLxmVsSbPfr9/h+qJ8IlOCWJp
eDgnm3qN8dnTR2eRqJhHBVEKXq6sZ+ve/bLpoikiCDi9Mr9BX1Nq1+TzEPON7gO1
R3zmoOfGk2bsu9Xtazfev8ZNtgGKB+sB24o7vngy3MymCiv9kwe7b9yA4Iu0QccV
8RXIvI10iEtv6OwJRnF8Qt+zSlbq8agNeKeNHA/sPyQ6Gg1iKWZn/04A6mXWRTT3
0zW+Hc5fR9BUK+vomNqcDnHwZOikaXed9cOsKdQP7fblP8uMJphwIFy8hL/SZrSv
jtSDLYStVjdNcOpjiogDWnUT/lA54I1KNsRlnyir+05ZnWb1unw5OCJxqM9MM5gu
ITRZ6LzwzLBj1/Df55RYwGty0DPO3s4JN7y0ztiCNCfL3UMD7OvFNRe4Yvpv8PCQ
ZrHIRY9H2HDmetVwdaUsKDlrx1961TkF5Vcr+FC02gkVFS7lyLIOVZWOlkhTaFew
4OEqXgKFFzoRCX2JJ6CS5eYcjsMuZqqTdtbHwsQ2otmNC3PMokaeYfIWkttMn01h
4uaMj/dygfiEZc8gwmRGY69I2cFZiY9OTuZ8KqT0KV11OOJpUv8F291M0KmYgSPo
TJpmJvBg+o/P+ODcnv2yAOtjGLr6MmrDYDjHCAYnZHkOinRy0CgKOoD49VQ77RXQ
AGHGY6gw4FyCoVe/BJTafRjpOKVsrEHsIdpnN3MdnhzTOECv+r4/bEuGN35IkctL
q2NGeKNHhbMLEumw0qAS/5jZP6K9O/iP9IqFnZQE6V+BUmkXEshXNPgqWskrLRyL
YzD7Oe2s1qDkb5z75AYkBClWdT57W1sd9iEmIkJKrMl5VwE5D3JSrRZvMZ9e3Eh6
zeKFn89jXojl2/6wgDjg9HEUoIKaNhIc9u8T1amgB05iU2GViVcjQ+ymrEYoD9r+
bRe6RWPR/z75wcmyFpOnePiutaA+1K2nBj21g7TjHJqMF4y0qH2BIo6+Y1aKnKaj
wrf+1ravI8mNlq8kEowHliD4+7AFCefBvFhNoFOMKdknbio1owAsZ0tE5Bt2RzI2
PU1z1nlQPlClXN5hCV8RkRjxvm3PQGZxP77l9yAOWWCH8UNCwe4fPOCdpz4iNZR+
LBWgz5Lv+en5yS2h9BIGc3l74xFdGqSwn0EIJG2eVaMMBsqYcsXhIN7WHm9f2lw1
xHXhilTwzjL/v55ZoC+yw0zPXdW7DlugrsxxiSJ5WguwTv92zvHeJ2n5gKPs2LRu
dUneGwla34vgwBq7xy0Xin8U54smWvj3q+m9LfbCmdZx3f1vWSJs2bw8hze+J/Q5
/DqglX81NEMQkRP7oZrJfdGAc5Bg01JkeBq43GnEasnKQxCdnikpI66VbIkWnhj4
2KzFa9xVieXbsHhkcnn3QYUD6ojEUp16J2SD0g/PCvBlo1Tk5StIvSoCjhNYf8G5
b5cWGI3jGMtHzOLZMpp8468svyT1LugljMl6LwcSYSOe0LU+XK/gTlGAuJTsxgFc
5aAzZ59WmbAa5KUOS/djD+CxahOHtaZmqx/2xbEfPjURiKfEODhV+L/9hnDEBlGM
w7jsuHBNQmUN9M1g5yr4xZS4dpwx40FE5ntsYNVQLbCcjD2BfUrgx7Cx71cpt5ux
hHkCFubfviUPj3+ZmOZbjQV9scsy/aUzZprS/JxF+a46LQz1kQkmrEAu0Od8e4W6
9XlPVPNTNQ3iZ8S7FFAWOwV+mVb069fgQI45JT77ve0+SWVidyFJCStqWReG/5Xh
z/kJ9WfXcvPQZcdxdRBGzIDEHtUp58MgpRJw2SuE0bxIZQDu/H9NQhEKJLpVy8Gv
+V9zicJ2DmnG+Eoxq0nRQkgLOaHIBK2Umq07ulHIcfAMlqe6aU+eJiY48lPgJGjA
sQQf5qlLlg8IwJT+y8jIKYUSv4/Vq8CuZSVp3BMQQOY4Ac/Zvwkm+LXbH6qa4QSo
FPFvi9VPlZICufMzg40H/BOHfYtN88qf6i8xC1ljQUMz333Edj4IQOUeM9nvrxEL
bsCHohJgh4zpekh4YqmQCbIZKt54sV/1Y8yvxkccBc2K6s/iI1IJnvevKdGew5TA
fdV/97ZmYH6gV/zRYsx4psi0J+klh8clVzjKGGZpv3fVD3NikBxsCGJ30mQaum1T
YzsF1wU4hOCcbWWbJzRVFdqCEgFPftYQmQXwRx2I4SY9sicuB75vH0JD4CCsB7nx
75b0hjNEklhXAGFL+gf4oRGlqj8MU/gbhghZa8l9JYoJrmavzLZ+MX4FPgIevYAZ
LU7LOPM58ja++gjENtNfEMWGIYIbFMokDwyTPBhHk21EqzGqabiFztpGiUcFarpD
vZnUtipmoffPjWN6yZLtM8oBO5fPjKCSCnJJwub+yWRDg8py2D1z5pVORANrAiei
SOjPV8/hUK8FbyDCSbXXu1o6Vow7oCunOy1a+LJDX20lNeE0k8l2DIrYLSYYDbka
g1W8WasnNXNrHP/c4127A1RUdGboAO3Zc9IGAh0tB2XEpRAchNioSLLel7xafDYI
lWplco4xHSNfxuzgtzWI61WPFBYilIoYIYo95KILPDNXlthUEXrhmqWJZUHOWe2c
LFWnEzZAP3hBE5NAqNwxf584UMFTEguJITZF37d41hJOMc80UH6TMJfVKlZoSpop
M3qaHYXU/M0jZM0tQOJFppKGAUOOrILTtdKlvVRwci+Sq9ENySY756PeX4O4UJwB
KKenrZBvjJlYnz7xU7nYf2u5vaKO9HIymBxkU2jeodKmd8jMLXH/nq+xtSCIU2IY
MRznd0kTmxg5BLS2RnQ7DFrUk0dFNnZTqU4wvBshuSodUa9drOJ8hXEjxKVDC6d0
as5v6JFRyOOrzIysOstuwAD95g5GmUIEBYUiNzyYjxF2f8fghKVrAvH8xukytKhB
jpbAjPv7FVLrFGNTDbkhR55u1KyxvGKorpsGDzdoOHAZi2px7GKUkAeQil3KXU7i
wmkVoMOKqxvDCKFc43H4lcEKGYiH169BedR7LdxTzCIw31fEhZyyLyRuOnsHFiL0
gB5JSZR0ubeKtXeF0iXvLxCKJBc073ywwamF5SIPtiInV+2Qf4urPYP+VCdv9c7Z
uMUmHofaciOd4Dn58oBmZR5P1mai6kYSaUgZBHbbR3k46KJOnipS/V9hYuk6kJ8J
MuRaCtk/dpVlWidG2vQQVWsBkMF8nzDHdoTZrd+geoqMXtJXOJbS3jTJIoDQXOfQ
zCg/XR1iJEy9qVF3Tv+W7tKcdUxXpNlCWhoWw1oE0sfRplZGDij/Bjm5Q3Djy9ri
qWXMKYFi20yc39kU2f6J2sxvqx1FYUD4tGOz+u6Cp2MjMxD2UJdQtEpK76+YgALS
nNlg7+0TXTnI2rVnQ0D7sNnaUIPxVImUQakW3nimS5CZN5HW3I5EIudo84KpPA8g
TrdFUQGkkQIq7gi+zFc/EqHtFTKLPPpia0Eg6unvr4jFC6n62JJ7pOjejhXOg+7E
us8ldLbJb94zp+qDWZvUxDPylTukSlh4ogHi3DWjwAFcwHIrErJQ5FYSOljgsrwI
ZaLUbaTBPopRgBGPKKkoV5JLSQ5rwY5Ja/OA5wQJu6Alz2Z68Y8CQCst6z2UOafY
KBoG6EhCST/zFUQwMvaGCDkAoy0fL27ouAoyT91qarVlvYVhyA26arXP9lnOUMtr
Lweem53HcIDXxmv0tWjfJJGj0ttQkWJdX8+P2ewV+5j+2iidktu2yyBR8X1rUA/P
c3Q1pGAiF3UGyVgHN9Bs+nzn09L2cHwnZubTRLfYBwqiEXOJXSbImATOH86raPfK
Upu4ZoeLViRcXA2eLZocstHL7K2XXP1B7xGjU5aPoE3Ch4SoEsS8IGXHUwcG/XqT
t4TsxzIkuczp6ABZM1v/EwiLCTYvYkwCMM2YGCekgjoJqCNP2owmnYRhWugmAgsL
y4nZURSTSGDbqNu7OFiapbHGmEWyzwLZbZIOgXNf/hAAWpZIyadHe6Y2u+/sga7f
HA75DxEZDez2PA3IPu2wc4FWbG2KHSb37SGPkodmYU6OI2rUH4W25JCmtDG5Wg3T
QmBzh4UksxNXpoxjqNdxNhWTP+6sfW8ZS71KV0HgEk/ygspSQbb7bnBgYNQXweq4
n+nM6KD3qEaxVHTUteJ4ymC5dWJBt5aXEdLzBraAlsXazm77CQgOpkpsnD3hhoQ5
wilT9UrqbV2AJuRQiqZVKANy8EgKaDGcDFeSF77KYkg1bz79XDriDEfG5GDyCDnR
moTtF6VCJRbjJRIXhzNPHRBx5xndvBryoQzTjhZ+HZseSVooawJdpcUe59nCHyXW
pBSge9Hnvw58VQxPtmkauLHYnZEIAPeyljSIVMZH8C4xt9JuxFnn7k1BF5HEbiM1
GAxF86MQkFoH8wzMnJjSbJxYWg0Xh84cTn2Q4Fv+00QfpGEEZ2oSx0NawbvpYMrQ
3uoqC1LQqpbh3MkPnuNlqa160lBSgkmsu7OmJDB6yzhzIrMXykLTvgJXRTA79z37
ShHl4EFoL/UjtAEo/nOB/3ODyf6hY9+QC3Avb56ifJnT9Xa0Bv4RR1rgMSKzqn9l
U0w9lAkHmoIsanBRx+98ZVxzMW+GEujtzvQWdxPqGSEWyOCT2oei/FCHenPIrA+h
p6+EdQeaUQT6BrsXqVVbVBSTdTRMMHIx41Ju63v4GhWmItbDxKLQexZJHSwfnC9m
YrRkSaeZQ3p4OTVeF5IVtGIusEKnwS4VAUtoLdEG9e7ArsHSrencDnmjXvMBdOKg
D4vfvWchu7b4qh8rT5vP3paledzAFCu4oEVpNOW9nZIrPuNv/TBvWgjRiJq5Q6bt
B0TqSTTZ0NAQEznngxEBTc6lh6V8m8mcGUcnHeoUQEolaAD5972P45x9Xetly3hi
csDJYegkeRJrMr04oVwzTgL4GpvwXGlAx69D6gkFsziDALIll0L0gYEemBlHVTx9
ZJZKXa3yVFpyNWX4A77VFGyLbDgXZfZY1d1C43CWE1Iz/CLTVL38CbM3odEabliV
NYJhaH+rMAMiONJNR+5I6K5FsZeOWnnWHfwT5o6cuEvNC/4U2dm89MmYKhzzcaOa
s/KR44LldDMOLqhlhdTzLo5tiUEA3A+XlQR0Gcbol51g4T+6ABTJ7xJo+oqS2Tmb
qHFF338C98hOzGor5QKaX62QKxIKoddkILpK6NacpfecC3JnccF4N72jBcAfjxDW
MBHxG/AH7WN/2LrfHAE81lWIHIt6dKqwELD0ywM4iJ9Hmr+MuiOj06NsNewb5DYS
6ioGy2o9DEGcncrgkRYz6U+lnw7pT0hcLXKsuAgrZlE7DIIB+eiGFXuXWmqPJ0hc
LNAZeCpjnbUYvyBd1X6A3h2xTK4g0CZRZKfwUg5Bf3qFFU+d9dfhsfW3QNhAX2OZ
B2//E1wdaR82vADYKtypDOaRuwLGmqh/fA2N52I4jB1RSZDlqfInamzs8z7RtkDs
xGvc6j9HTGqjfFdG5EFi3hjaBD/3H6x3F/f34jjM91vzsUfjltu89kohIC4ncEpm
rejNJ3vuM7Vn3Fffz7842o2eEJJXgRGJwkFa9uHHIxKNbpofmsRaHK1mtvJBYf1a
pm/FIxKgdU2BZAwbAVWY5YfvFTpq2tJqbxmB0HHz1JR85Kw7NaHOwlpjaWlMZ9t1
sPndTQyYs+LkZSEJ6DH52fLoa3aBEDRhMXiBloD86WfPzkCY+NpuD4XxWZG8ifwB
z5N1Vsy2R4UfTaQ64GKmH5U55nmUGH90CnvjUS8+sHCqTRR68GCvLGbrslNL+dFx
E268F7ymsudKNCcPDsU/RqOFhzJxEIW43JFhUQFyNKk3hmoyCJOzLAqv9Tl6XjZd
NB81J3Y82k8feaZHWcJEfY9MHwEJTT8ihkFuOWEBofGkil790+g4VWSuHqXpFW2a
exSk2vefBuYGY5YRmboRn0aVfE2rH94iC734+L6H52D9LRUwKAwupauD4Tl0KI6J
MBxoWy2DS7XuC32GzV6maSp4PR/qgFTXFZYmNTq3T2/EDC0telj57F+2BPNaSjbg
TxFJ48PrvHOB937MPbNpUlN5wCFPQhueOijUDvLzxKJ9WRSuFkMXDXO6W1pNs3Ea
goo/6v7d97T+MUurnNHi3b1XXA2sUhP2FEE9Zgg5FZMrZfxRIuoawgPKfH5A2MEU
3qJR+cVcm/ZLN9lXnRXzhfg5fQvr2xoEguOpoC6biK16DoD3z8m5oyZ1Xolo9mfr
khRM8j3ygXG/74ZSPsyquPVQJE/tuSH2qnfyuXM2Vx1Ku9I6j9rEjmA2jROgaxSd
08kaPM2PnHSimieUG6bDhEh+7fYAtq2sMQkjqARtstMgdoxNomTMjZHqE+0a6glX
6C/OJ3oZIp6GxjvZBk3KBzJVbvl8urM9MV7pJk/9a9mbut7aZRxMhKk0AYs44YrZ
C0vZHEk+9A5qSRArGLWFks0wkd2zeJH8Y5rF2mxhIdqm6xKHnGq6dc6pef+ftIzT
ReYTBq79Kmjev3acg0SszzCoEz6Jpd+bekhrtu0hwuhllPmf4hj9FwEsrmsASRyU
DzZwx277kv7b4YdsTRuiQbIs6zSE9hXUuYZomZ/vr6QUcpKhIGaGEb1AXjf1xi1N
Dl9XKSnJCx5uSRDF10YKUKkKDQecNbCK38ph/33ekVOScxslVsfyUSaVNkifwfhZ
br6mFUwa/KbPDLooH98+9nMu2T1TjQuMosCK/RTgJRoyRRNEQHAIYFS4LUCqg+8U
mxES44A1Djza/IiM0S3bVdyCEzXtw6YCxD7OJChWOv4LLC2g7f2xi6DQd1NmPexA
Bz4txZYb3M56CjNijiPMOzFT3BmaAXWX0S2RtoJlQClbd5Sds0FaMDRutAfhqrf7
00s7Jqki9rRhcEQKfz3EApGF1yl5bFWeaGkrhMnsj9lQJGJCP1VtLqFjZS2qAACx
+VySeOfRa61yKklZcBtzHrfQruDcj+c3IhZMdUyHcvj2Utcz0yU0IlqIYUAYPT6c
LokE7drgOzdrgKtWRmyTLa70tlfsYA66GetKyPP3YTG2i/SKH3e6zg9Fg4/VVUyR
lBUPTb3vE/+TgNT0Mf3qjxpmwQ4tSf7K/V2TLwy48Umw8rLeiyrBKj2wzzD4Qt7m
c0HF/EmOGdXpjboCdk5bZneYTVadheqhnWU4S6XSOA7Ij/6iqrYQ1Rgv2rTbk/um
e8UYfjLS6CLr2aP8uyu4xXL+pqrc+/X31BCgEsmqlzCCdPNuCKneJe95mDxZ3mXS
xMGwbz1ZuuFh8MNrIoYtR3UUc+63ovahqKmIk15SM2UsO6h3VWtymXSPO/cj8QSl
ewUYW7Pe8z2fNeg5WpJZF7kogDhd3lQAMLnjUdtw4XOGxTuPc3cx2HKn3PEgZzln
8h2TNoLpDzKY1qtuXkSqRaZEIzyT+OMd6PXxSEiPl4ggR+Coa+hmFniQSuv2w+Nm
MyPFLtDkD0/LbfI3zL4GiLNk+dXHCkC1VVFzogAY2Fcval4ovPSqOrT2UTeJf5UN
+xMQzXMv6cMSeGYQDlWlrKDqzRBT1kzYHsNj4grLjJ3M/NFz09kk9Xl1jIhNoPiw
4RMq7RsyCuTS9pq6WkWKtDMZZYItZKwa/4ekRMhbC4rgcLTq2jiLKzQzlVM5Sqij
OKXJP+qheS4nPJBDNXjP8KODqLuVnhwkzaWZ1HAThYsqS0zZL0CUCFyX+qdXgnlm
r9p4qIfHC/28dchm8dmKN1LitvkwAgFDR2asU3wIxp/cR/dALKonDIZ52+wu38Vo
joInbX9/Uo/MBzfeZy8UP/V3HsVpxldxj+Y01+u+oUyKleHNbG2D0MBphP15pltH
WDHDaU7g+WqRR/HQUZzExm8hGnp8u1euyzJQXikNs96mPmg0ifOpVlCzrWyjml5+
G3egSqgVg4efsxm5WErB7WmKSmI46sBBai74WgzaYYdkvbc6Q/ovXCvTscWJcom1
+sLrjSPOKk9zCoJFWdoTuv2doR1eJifWqkiwUV260AyUUggK4d+/MeUXw8He8od2
0qA16qUYuiXtiXqZcibkRD0TLT7KIqycq804bLZdzd1XyUcPNvF518jxkth+ljkf
b8XRP+s35nMBg+rSkyEwqP9Upsr9P+EmuNblGPC2Yd7Q23QNs5A1Wm503yY8IJBK
0u3eVomt232/0FuYVLYij6grB4ebW9mb+/n1ivLU/jqoI05jjfthZhzTrFHHUFMr
+Ekep/DvmJl4qcN/nC3a9AEEMZGbfT2Ejk3pldEPsOKOotFKG2Ph8mlHGWkzQv/k
W81ZvlW70q/nRcXoRdBjpgqfODW84FiNiMltWOXDAUtbd4mON9YdF9JoRORicjCE
5jIaQY+R6fdoNweKbE2/WDDtUG/pSTYmXstdb276xlYw2eSbsjIHWmHbvJDkf5vB
tSdGB/kfn0Sde1XpGgcZmulBbC/OFmYW49S2tj6K1Odo9QF50sKF1dJ8UV8A9dkL
+Fs5g5KT3gbHPZfP1YwxREOzEU2tAndSAcoqtObWOriKcOTVbpaVnuFFpy3bp/47
2CpaMeisEXddyg9v29wZshTryHwn79aL1b9OqkYqXG19k6Y5HGIaQUqtDdCA7x3C
e+THve3JnsuG514I+XuJxqEbPmrvJZ9PRDvBDgC6Y7Sckbu9pGKsD2Zty3bLRtzD
6wbPRzkbDV/CZNzWxlFcHOIorfE46+/wgEFRSspgqqgyA8M66prrjB8BBhXPqjEf
BarXQUSnfzjvEEeMdQx5ceF97zSh9e3eoufr/m1Qx86E4wj66UrgNjEZ2i4h0tAe
Fyek5ZA5dQpvxmrRU0HJQo7oGxzd3uTrec0ZYlYK6VvmHTlaFXbDgHhEAQHfEqkk
v1rigqkWVibp/X3eixf3b7ySe4Jgd2NmKoSI952pYxnAIKo97y374o/+gDq0qhrv
ZtnvcAHqvQU92u+XtxTd5jL7aUGl9ZAf+TJrAnhL13XAkikVVgkj198f9HwDhZUO
WYj/q5NvFeJMas9cU5HJGWuMS/JZFrkjOdunxBvwv8dG83bGGyxTN8gcCKFm/qTs
RpximFbwWA6oYHr8GSn0qmKP/U5K+zI0aTVS92wrVCVwkhs4M/04E+2OHYALKEFW
qTNn/Dqk8WrsBHTxcEAGU8hG07tHCSoOcjIEtEtXPAmr6bHbFMJPncSnpBR5oQf7
qC8iu5IewRVrsTsrLNBOq/lvXzcOj5iGVmJNKue39eRsDcFPGRF+iTcqc98pv1qs
Arrpb3hf5DO7CjZU0YhsL7FU6Wp1+IupIir2idL3Icb0mHTJViH9uAfxdlvneKbA
YLp8TjIXzcf3LbK9MGIDotyd82wjkk36+25dxS3J2Q5I1y4o6TWFoPtPmCE59Njn
19noKBvWyNNSQK84L7iUavf7RhRAMKahgmtjqevPaF8erzphoX47Qyrvpi2Is9Dm
CtGG5razmT7suzGn0cFpC1eGpPl8qBGJuzfBLmJRkEPiCGZqzJgL56UlvPfM8aY9
6L+/EKjBd4koKGc60pjvsWODH+EOnLmWVcVuoeUPCgCtPIgFU/MWg3JIfIasz+Mk
EwnoL6QEOu/uHnsRTt7+pA==
`protect END_PROTECTED
