LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY DY_DLY IS
	PORT
	(
		nRST					: in std_logic;		
		clk						: in std_logic;
		
		sensor_delay_in			: in std_logic;							---��������
		sensor_delay_time		: in std_logic_vector(15 downto 0);		---��ʱʱ��
		
		X_Raw_A_Filted_port		: in std_logic;							---���������ж��˶�����Ͳ�����ʱ��λ
		X_Raw_B_Filted_port		: in std_logic;
			
		sensor_delay_out		: out std_logic							---�������
	);
END ENTITY;

ARCHITECTURE BEHV OF DY_DLY	IS
	signal sensor_delay_in_r1	: std_logic;
	signal sensor_delay_in_r2	: std_logic;
	signal sensor_delay_rise	: std_logic;
	signal sensor_delay_fall	: std_logic;
	
	signal encoder_cnt_rise		: std_logic_vector(15 downto 0);
	signal encoder_cnt_fall		: std_logic_vector(15 downto 0);	
	signal Encoder_A				: std_logic;
	signal Encoder_A_L			: std_logic;
	signal Encoder_B				: std_logic;
	signal Encoder_B_L			: std_logic;

	signal Add						: std_logic;
	signal Dec						: std_logic;
	
	type delay_state is (IDLE, COUNTING, FINISH);
	signal delay_state_rise	: delay_state := IDLE;
	signal delay_state_fall	: delay_state := IDLE;
	signal int_sensor_delay_time		: std_logic_vector(15 downto 0);
	signal int_sensor_delay_time1		: std_logic_vector(15 downto 0);
	
BEGIN

	process(nRST,clk)
	begin
		if(nRST = '0') then
			sensor_delay_in_r1	<= '0';
			sensor_delay_in_r2	<= '0';
			sensor_delay_rise		<= '0';
			sensor_delay_fall		<= '0';
			encoder_cnt_rise		<= (others => '0');
			encoder_cnt_fall		<= (others => '0');
			delay_state_rise		<= IDLE;
			delay_state_fall		<= IDLE;
		elsif(clk'event and clk = '1') then
				
			sensor_delay_in_r1	<= sensor_delay_in;
			sensor_delay_in_r2	<= sensor_delay_in_r1;
			if(delay_state_rise = IDLE and delay_state_fall = IDLE) then
				int_sensor_delay_time <= sensor_delay_time;
				int_sensor_delay_time1 <= sensor_delay_time + '1'; 
			end if;
				
			---��״̬�����������۵������أ���ʱ�󣬽������ر�־��1
			case delay_state_rise is
				when IDLE =>
					if(sensor_delay_in_r2 = '0' and sensor_delay_in_r1 = '1') then
						delay_state_rise	<= COUNTING;
					else
						delay_state_rise	<= IDLE;
					end if;
				when COUNTING =>
					if(encoder_cnt_rise < int_sensor_delay_time) then
						if(Add = '1') then
							encoder_cnt_rise	<= encoder_cnt_rise + '1';
							delay_state_rise	<= COUNTING;
						else
							encoder_cnt_rise	<= encoder_cnt_rise;
							delay_state_rise	<= COUNTING;
						end if;
					else
						encoder_cnt_rise	<= (others => '0');
						delay_state_rise	<= FINISH;
						sensor_delay_rise	<= '1';
					end if;	
				when FINISH =>
					delay_state_rise	<= IDLE;
					sensor_delay_rise	<= '0';
				when others =>
			end case;
					
			---��״̬�����ڼ��������۵��½��أ���ʱ�󣬽��½��ر�־��1
			case delay_state_fall is
				when IDLE =>
					if(sensor_delay_in_r2 = '1' and sensor_delay_in_r1 = '0') then
						delay_state_fall	<= COUNTING;
					else
						delay_state_fall	<= IDLE;
					end if;
				when COUNTING =>
					if(encoder_cnt_fall < int_sensor_delay_time1) then
						if(Add = '1') then
							encoder_cnt_fall	<= encoder_cnt_fall + '1';
							delay_state_fall	<= COUNTING;
						else
							encoder_cnt_fall	<= encoder_cnt_fall;
							delay_state_fall	<= COUNTING;
						end if;
					else
						encoder_cnt_fall	<= (others => '0');
						delay_state_fall	<= FINISH;
						sensor_delay_fall	<= '1';
					end if;	
				when FINISH =>
					delay_state_fall	<= IDLE;
					sensor_delay_fall	<= '0';
				when others =>
			end case;	
			
--			if(sensor_delay_rise = '1' and sensor_delay_fall = '1') then
--				if(delay_cnt < ) then
--			else
--			end if;
						
			---�����ر�־���½��ر�־�����Ƶ������
			if(int_sensor_delay_time = x"0000") then
				sensor_delay_out	<= sensor_delay_in;
			else
				if(sensor_delay_rise = '1') then
					sensor_delay_out	<= '1';
				elsif(sensor_delay_fall = '1') then				
					sensor_delay_out	<= '0';
				end if;
			end if;
			
		end if;
	end process;
	
	---������з���Ͳ�����ʱ��λ
	process(nRST,clk)
	begin
		if(nRST = '0') then
			Encoder_A	<= '0';
			Encoder_B	<= '0';
			Encoder_A_L	<= '0';
			Encoder_B_L	<= '0';
			Add			<= '0';
			Dec			<= '0';			
		elsif(clk'event and clk = '1') then
		
			Encoder_A	<= X_Raw_A_Filted_port;
			Encoder_B	<= X_Raw_B_Filted_port;
			Encoder_A_L <= Encoder_A;
			Encoder_B_L <= Encoder_B;
			
			if( (Encoder_B_L = '1' and Encoder_B = '1' and Encoder_A = '1' and Encoder_A_L = '0') or 
				(Encoder_B_L = '0' and Encoder_B = '0' and Encoder_A = '0' and Encoder_A_L = '1') or 
				(Encoder_A_L = '1' and Encoder_A = '1' and Encoder_B = '0' and Encoder_B_L = '1') or 
				(Encoder_A_L = '0' and Encoder_A = '0' and Encoder_B = '1' and Encoder_B_L = '0') ) then
				Add <= '1';
				Dec <= '0';
			elsif( (Encoder_B_L = '1' and Encoder_B = '1' and Encoder_A = '0' and Encoder_A_L = '1') or 
				(Encoder_B_L = '0' and Encoder_B = '0' and Encoder_A = '1' and Encoder_A_L = '0') or 
				(Encoder_A_L = '1' and Encoder_A = '1' and Encoder_B = '1' and Encoder_B_L = '0') or 
				(Encoder_A_L = '0' and Encoder_A = '0' and Encoder_B = '0' and Encoder_B_L = '1') ) then
				Add <= '0';
				Dec <= '1';
			else
				Add <= '0';
				Dec <= '0';
			end if;
			
		end if;
	end process;
	
	
END BEHV;
