`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TbTIXoihkihLj2lQzl8GIfjqmcU/anP1Fz6NLckPCATjUp82z+KB0KN8gPssOOxh
pVYF4VyLpaKfj6WutgtWvdfmcAtVMJXnp2BWdRmMpQSjw4VUtTir8fYYDzv1ynkA
n/3d6WFV9aCoo5q3FkqW+Z7sQ8NHgwh1CAj758t0SHU=
`protect END_PROTECTED
