`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
rTVrc6fwmHqsFc9UEeR3zuBRD2+YhLIbdiza6JdtEYL548Wc8IxIp+AGs5QKcUJo
maHhp3yW2xMgh4ru7424tvcNun4K0h4BY7JBLFyKIDYvjHk3HvvfKGCNnKgClY/k
12lqD761Kd0FyQWDyeTEceM5cQGA0l9omj7SqHysbTk=
`protect END_PROTECTED
