`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gkdFXZu93R612Bu5GHiErJvkVh7SS5tE2KzeTgXepFljVl8BX+txihRuE/tmmaC0
LLEeVCaoUtv+Bq68H9tF1EdBDvr1xiKI2RdHfqrCs6HZt6AZjVvR4sKQBqIWQj1y
dvBeWQRB1yuETxWRixhaFrK3kZFbLAl8+J+Hdf/vasrpkN+whqa8aSnYquogB7Fy
fPI/AosGNQMfvICtfwme4ZGFEKN9tydBEuMcTpdyHMYJ8rwNGtYemmIZ9CydnN9k
BJy+1knndvid28WJIe0HM85sThF6fKlPm+8qECpcsHHY5r44Rz2pR3XaOEqkHJEG
KchNegvMomFl1oVNQmf0CWsWoCKAreCoqZG51goWTwpn8qEfk3NjFxd9UGhR4oR+
1z+FFCoCoHkmuePNVmvJBLhJlr8gMjJ5J7xoEiQKGUlejD+4P/bPQ07FIOIvs15F
20BsvOD5yFamU0GgCKR7vMa7ZSHNI1l37ecBY77lEH2xH/t/B/MvKXW8LF7h7Bcz
dzwlwQxKA9OAJYImJ01itx96MNMvBdkJ8s3+h5pKJPGkdfuELengjdQQQDJLxbvP
ugYgQEWcfhFUxqYKhD3PqtnjDAePR1yZpi7PPCWhTZjrF+0W4ys6mOfRRguQXw4G
JWBSI6lLgZA5KQQQQENh5smF2WVPuI31EMaMjFApQ6GzRd3oRinpBnDqTo4u3YDx
56GkY6C2iPVYlQisArjgH4CAeqF3RBs12hsannjo0q8MFMaICAahguhmtX09yg5H
svChU91lArV9WE7hvPPf5yPYGiy8NC60Jwu2rjeqre3Og6QCTNr604HHoeIC88Qc
F8P1+qXSjmGz9yynCPm0iCn9cK/J9IN1BHo8FyW7pjqXijSS/xwqOK3uYMKIvw6n
Lc+JQwRUVtVYPYNBwimZuKTJ3BRJUD40ugeNMiKb9HA1mv0Y8MRb3ESYtvU9UWNb
8NE94oC1JoTUdkYHLtbHi2QT4POo/gKXstE3vC44A703jHGW8kkOQ87rZqm1xa9z
cvVts6K204KvsshwhTP9NPkTjL4zLzMKCC1WPIEq8acD9Ld9s2T68T70cpiDoLLM
vC+MQXAqJ9P8vMz/ki1/sLij8Dcz58ZNFAyWo5Owf/8WSzuGCFQdRvsmbPXRmBeU
z/OMbL5fJDdVUGMPeR4sYAsBgIZGXzMH0VEPnK8aSGgaM4mSyQLRIakPCwxed72X
zIV5iCfn/ci5zk20oPCJxYpj9J09KnvZUxqN64B6SsBlq11JJfIkAl2uQb+joLh/
jaNFSThY+n8q2hFVVGXxx9VJGFfn533mw5oAPRk0vULkAHu+959c3Ut0TbxaZkM7
Zf7US/6RIlSd407NFabgUsy67zRQ+K6wyeqdSSl+vPCR6XNFA8kwwQuNUt9XHlU5
TSg7uj6z8kZluVy7L7+a42OTRfab226WS0mY5X0r+se3EpXnNXTNs49lhYMF0mFw
l59bHDywz2q3n73UmrgFz+LCNARO6G0bFyLVdtyaiOGQFVnlusCOMvN9PtMc3ko0
Qbo20bd7N9BF6peBmGFvvGct+DNHDBL+Bd4GOlh4hM/x8xjghUWnlhjOUiLF16G1
+8F+ZvRzwlu0fGO70FemmKKJQGcLvzt4vwY2Ozzk2S7WgPCLmnQv0kaUskxZVeJc
wO5Vb9/U2DCKLFjenbbSerbmKcQurWx0ZiVtF8looHRBh0FhpksxZDP4y/0xnrpV
fdgFHoMOFy7j0jjol8kSfgIeRhcdTGfksScoL9j3t89xFXAmJ4TzGUCuQOu2ltMH
pww1v3fhOHXBtwBP6zYzqnCTaUjrdA0efdeTvYBvUjHtPexJzQ4SZFOUmvhcsfdA
vi8wBQQ5UMj3nFpFNE5Ni2dJyXB19R0bB729oYgXg8F1C/ZKwujZ16nEXludh/HX
jyRqp4Ov5LuSr8I5fc2rVPLFELgStNw7hP8SXP94b5gLh4ZTRKyrmE2laQ2d1AWV
XTa3XbMBXrl+3kMutPZ54kai6obcsC0J+QsmVxaTobZIHLwaW8tAjvIcIqtJMCZu
ceFkOggza3mMJL7ZMjBb5T+0MjhOkyUjl5CEF0PLNltyC7Jkx+06DrI6HvbTUvLt
jC+/VoR8TAIOFNBPFTBP5QQ15H8yhEy8rx9O1HBYVk5xWkyvHx2m9CtouxuRXDCR
UvRRQl89XU9i0vQfMFSUNQKVpS4BW0KCDIyLVnEc/rsg8Z+G3T6QGsJqntJvgP4O
9tkCWcK7qSHCviJLg4eO2FvnhrvbmzySIIthJXhVEhw/YHvUhdW0PyX90CWnJmID
T7rW2OSii1is//7YBzeM/19njLwKOxSwM3H+tVwZT0wb/jfUXO59cKwu+NwU1S7l
r4Ksg+/Nq6AGwKSWEIKakwulGfjxXcYGqH2yS5j8qFjJ3th8meu+LcXrEtCiWiTT
moz9zPkFBBpVqEtKs0ocnVh36pa1CPVggRLvbKUyAE5OE0q3I6RryIjCt29XlF17
yauKi/FudcEWsSGwoSsEHRxvZqRwKilCKZJX//qMz3d5J7i990LQfQbcKDKPBU+t
sqcD0EsyRXuMJwetkS8WFz+wZ1sw42w1J1dGo6iPNQa0HLaaKhTlS1ZugTadkLBU
ng4Zame7fD8a4ILm2Sdf3owSGphg1FjzrYAXmVzxZt7QqFlKwQRT7wN4Fv3MKe8D
fbr57X9nylS3olfATzdYOAGcDtY8gBRmXnYiSF8S8NAPMv7cLOBbZugSdoWaFTsF
FcdZdAgsTDjCBtI5Q+VYvK4yhgANomHmjZx0clgAgJTGxawXrvegUfYAMI06EGnx
7hwCu57R4XEB3I81ehJOBnZ0UHDJs25kYTLlQVnSwVLqRW2wE3ZQ1SnWXqyuQW+1
M4E9qrS/EfMRXo2ms6OYm9C7z3fHw33dEXS+Nix9L3cgUB5M7Dj4P9/G27mjVb2o
Eu6umgMC9336yDqpD70ssfr/P2jpUBwJXZ6LDiB71g5QujFNO6wdnKZrkkZBU76K
bgkWGpTibLfLZp1FHI+AP2UVQOrdsYlDHcwu/VRT3dmOh3mRmBQzAEMRm+kZltdK
BoSUx3/mSooOC2A5gsQlZ1ZY1NBBKeDxVJiX3deP0tsB+vd0Nn2t3xAOXCNmx3I7
FDoPRQOCNSA/VMIIkhKBn9pJUkcP9ewhsPp8lNd6pN//YjUZfG2BXiWL5n379kYD
ixuWo1OTixwmGqDXNxKyW9fHeDsvjvrj9umS0YB0qhKv413x/GuaHfIOmYti7RLY
yVQBREK7qcJ/qylcnAGhYn7Vyz+iXSAEn3w50+VeCYHbtj1Xw0+sMSZRQYOwa/06
QyWIiylV13d/11p6wCRgXQNd/JxmnI2NHlultj8w5wnWHl/HqMyLo2+p2iLP2e7A
o0kys6jzyYGU4nsFDABPs9zRRsI+ZeVvtg/EODH2PMDI9vjlSzpOdmzfAqggoCOE
MDN4bGuCZYsBIn8fEoQWgj21gw/iBzrb9VBZN/XfwN+Yt6VzRMglU3o9BbJeUzj1
rlV+cCaaIdQ9+wbyDTGUeFJkSlSGLd0NhTA0EapOHW19ka1pMZmM5YucfX4PG+Ow
jZmShDTsPCn2Z7Jk7MplGqAOotSXZU7xwvj8vpl+5sSgSh5ArHrdGBqlDtd5E64c
mVwr1LmVFh6/tDWieMeiAThmSeUGVS5cUtdj+9g2wxyo7rwsb09uxnXdstuvNbop
C1lP4yWWfuscsEJUp7ujdc/shRkbN1bTS50BGcOHACMuehRtXivPKwR3NHt9uJz7
PNN7enuAYlTqWGPQgS/Of0VtHzlr5SZCdH3Ip1N77u3G5IBVBgE0zzOElg0bk5I9
a/QqQtC30XO9HWUWI0elnxaQIlGggCTvM5kN0CErElTChdWnJvaVY87KfUbltfNe
F0DGR0sgqzXxzbx6dTYS9Kg6CUFSYp4S0uMxVQZx3EwDQ//PDCtP6qForMpcdGvp
1MHsWjNZhSmk2iDxcVjiUEpEE8LOjw1FhtTjMQbvnFhyoQmBVWjOKIq1Cp8z+Z1H
gppKFNmpuRzmAgpC24Q2Qulw0j8Lq9bPpE+sEKTRgOK4C8+6qzTH0/BP+09fPhB9
IlAL2oi4zX/ArD37RjT6dXIxlOYdPTl2loWPzCMCRRExbrQeX3TFyhMh/LmFp0S7
2iFEkU37to6mHSUozsFxqj4ndjs4b5ME3Aps1m7xGo6rW2VqjjRpy+ldnqC4/sdU
kg6cHBYcYaTUZEXorACeY+1vwYVFDSLtB1uaW9yI1WBV62J6Zgk9McWUwGQ+2i/d
XjHlRQ2gUGXhhojZF6AhHIqRAH6cIP6wa4cTVEGIRB48YmdQxnEMIMCRgFaHghfT
4IEYSaiUZ/xVAsnQQ3Py5r9hk58TZLic5yuPujD2z7HYhC58LuiZ4y1QFH8MbpTg
+DcCCKlDF7nY5HiVEITamRg/audFwMlXKEjesAp7RB4+UCT1QDWDllEl35k2oCA5
f0MXm1TjVdDL3Q6phw+FOcchWHMRMD7wO3q4bnwJBfSFvHRwQwcpvvoLSIxYjYaP
vQiY0nlSa+ndVrUqtVW+pqwiEVDjrZdEx8HP35lphlwFolbR502S/pX0s65uDVAJ
oLUf4LqmmhJvdXwXF8Fdt/iSHCWV1tHYvCvs83M9zgTME1+COF+k1lcZiBHksOZ0
eHfzZ4vQnC4tQiDCngCnRNuJlsz5g/9S6n9+wFY+xfrDn7xI9eMUSgpBDOwPgXSr
jRMUbFTz5qCREdqYCAhJV9eWTsAeVPJ2AGEc9418kD+DlIY+1bkAJFRR9KQLJ0aR
Roch/doZHhhPn4C/jZDggapGJ8QwwIyl1tG1G+8LJNsd2+TkQ7MyXO/wfojK9bj7
AEddOeS+fY55bo3nxW2xtcM2Lb6hvkLPoE+cRcqnFuLcipAdllXiWj+9YwoHF+dj
xGPj2U+JI+MFq1PK/USWiHQI0YdegUSkwUCwtGZdZOQ46+AfxX3JvH5rSQ8xpL+8
QHZ/vrs342Kkw+a5qCCrEiOQUmVpB6HjynpeCssSc7RWCel4rpnq894sYMvsgP+o
BDZpHi/rtPV9JNAmJK7f9APWYaWrpXSvF9EC4GmIMvaQBij58hl9Nzyf8fKR8YlX
modHNFnZNIJOyhnS5EaW8As7WojZ0no0sk9xJI9KJKAgX3VFm9m0VrY56Z1EOH6V
qaCM27rOtigQ/+5/iEIlywqF7ZVS0PkwwqLRNlPO810XxG4pt98Br0wlvcIS3+UZ
2LnxuPTJ9gC/lrmKI5k4i1YWkQu1zpRB80vEClDvm6A+tllvT+3niuz74rWJWoVa
`protect END_PROTECTED
