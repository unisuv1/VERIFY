`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
T9+gahHCjqDvvmlkM8ixD1fqyglxkBRTQTEMTaupc3JpPVTEYvApk9ww0t8n5Cen
pcB2b2I5PJSuEchRnznyH3Dr6hkMIs5z3TVmVwByvilbhGukcC1AVwHt4LwB/OEp
BlfVixrGjr/bjDPFDPWvPG77XwZp9WQSfRPlBtY2bQ9kA8rsbB90M4/j2mGVwyYk
VNoKC8EgVRUQRUWnLJnyKCcR4j5I0q321J9zRBvntW3f73qIk+oU9TsCcfNTxLGz
BTpvr4n0dbDn2zW1p+NBLXxltHVn5SNmbdGA79o2utllLtqMYPMRvO5GK3jfpdgU
Pdcm6q6Ko8d66EfYTTsYjYooqS12Z0ULXJvWY76Xul1Uh7GBKjPyq7eZDsMirh9x
qQCBXuoPT1NPWZy7iWRRtpKVR1rU+Xm3EVLq5y6TFhwj2X9PMmSDF9bXI+Z7k3f7
ezDxEmM0Bw+0hoXGkCOs7TkkBvdk47sVd7uFD2mloRTvXgc7cXV7v/IAfvfN1d7v
O6kcjBw3W9IfnH/iTPIQbxFogbHzYLQ5WwYdrO7vpI76/CPaFe0hnQ/D9evvPeL9
ttuI5B+NjcFbUGEmLoQ1IQA3tY4lave3kgSr+9sBz/V/MjpIwPxiMhyHeqdKWchh
hO28FPYpMm9Emcc0Vfmo5veD5qgKnr0clnmum6L8SDWrkkfJvkoQsYsdSayvNdOO
vqDCVdbMvNYEGPC2p1l63nqhecQnhs4LG6lszPWYgKSL+wZTZLcT93kDW0AGsbOC
QUrkGxqgNuuIXbTWYM3m50EKPQ9d+DjJpspUu0mnZQLEihBvwQQjoe26LSTmWd8f
/CyzZOJ4Tzw84qrsr4H8EKgyHXECCyuTIVlf+49R4WJiGKFj/XKjKMUE6vFDAvSD
lCqqoPMGnaG4OTt6O2oxU0vpfNl2cL3WJ9PchcvJSpNfC6uEMqx5Y+e8fN/06ZXi
R46FxKFrQrdVwOndJfN7PvXlYUslOInNQsCWqaygXJHjORex7+GkKRG5Mlq0a7VV
59b596HJcopQ0TbhINdGay4jGG9iIRwx/NuUFRq3gmrh8EGUOTatoMlw4INL6GE6
SSbTQ/0AH0iiUsm7hxLXJTT5FwBf9LWC0SaSiGRP5SIFgFYTevMEURIQG+Lcj9WX
uis8MscztS03gRI23mhKvnqn+K3MckNFVmxJDbupix8kJWhOyXd783SJRUBtL8Xo
7prcsChZnRQyOi3ZydFSsWNJl/cGVkmBiY2LNcFHnN9/MJrmXnP7AT+pzB9WAwsg
19M99Y5E5VJe8EU1qPC+AZsplnwsAvdWQ/AxkX5yVgiKNsvubSCiew4iPBzjXqEr
H+R1gpRoppSjWwOH1E3iI60Wk2egvJ1IwkdB4W82OpIjKIzV33sBY/+rXLxV2IDa
hMwtFXzetMosswvndgB3YkS4WyowigrETP3depGxulTwJjDvmKzJbA9KyDSVPT9V
8w9t7CVPjat4n0+jKR/CO4w+cUPf8Kxr7QRpjgYaJXSEGXcOICquGi66sZLBtKq1
xMDm5vYd3sBlDUufe7wzld2Bo3TfB7VLOVxRs4X/ZD9I6tuB5rTleAe1T+iEcX4D
Op1VFP68RhDEE3lmTHdcDEoig38oo9v7qUemJKBOOp9+T8zm+hH/KJ+IXw+3Hy3t
ZpZvd3Rh1ttBmHP+4A8WNEyg/jYv5msW3pqsGg9kJTg+2svhvS01R036qHVhs2kt
Y/0HlWPrvogwLq8BT2eb1MOShwOxjE2qTD2k2URJRIIPXlDnHyq0XtKyTw1tXaSm
`protect END_PROTECTED
