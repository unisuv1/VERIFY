`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bMA7NcHKxjhgjaI1iyQSBUkZk+KubWGhvj/6oC4j2V8nqqsvINhstU6Yybft0+Rs
S0noIXTbY0K+SxFU4UtdxBap6rnQPNEIFQJCn9uT2YFrIhijxHUA8CLC35PinW5W
3Gnjf6q57dieQBqVK6ISYxhpeWygCcmJ/bEwbXGzxRpbfvKyjCO6IdPMAabSR3/D
t8h5pUr/aqWguktWIap7u1Hji4sfx3EmF7A7iJrVyof/Svp5ici6L0v+r1CZ6Af6
NoMmZdIwYnObmhP1fL+R7UDgV3ZytDvgEnP0IJIK12DRjKUlpeRU/AC1sO9ngIvx
2jpOw59v9uUTCxN3clWjmDGUGUa6sBatGreinl+M7wY8orKPJLejz7wVc66/cBaq
iF2+Ai/vUjiB4qVteuGlicggrYZce4OPu4zf/ACGA7RoNRpIVtXI5h5cAh06V9pm
7AI4wPjKsyxkICDABiHO8VI03JImvMDZuP3U6d9ptASPlijmZIqjLvIJ/KmMluxR
BYymthyiA6ngaUI5Kor5584SBe+keC8QDO9M121/nL2YfNZH2u8jJwkO/F4w+17Y
iCKzyvoESzdgcpCNOc0S9SZX2U4t3DUghteS4GwoGeu+gCkIcTc45bzqEvO54I9x
mZBQgaIfUad2mNvxwt9zLmYYzLtfXfZcovBM03Xoe2ilDjgqjksxpGvjOJhfww8+
RJrQUla6mMAkgK9XlZZYHyOH2rY5v26sFoR8p6ASuN3VkFYad++kBegFXCmiQ2KO
ViNXwilj9hBNt9p2Vsq5Ys6f8P3Pyuv7wv7fibioLL9YMD0kbGfVugU5fxTIeZCl
zjd2uHD+eaYh1qI3HX7jEQy/tc31hVYVUGUg+7aNBZsyC5ua7m7rF2p5Wp6MCAN6
8Zj/e15yv8KTZMO4Tld+ikL7aoQCV2vXmY2RJagMoYp7j+a28zW+OSUCIHNMLUcX
az/d9O52+QXDVhDpXw5nIXGyvNjLA2ry/JTGVuTHAd6unkKF2fVQ3IJAN28EkUZS
XCXCXjS4Z2FJKy0HYympzH3E0y03Q+HWp16PdJZ0ySVuffTGd24jKLrKEJKCgv9O
giEYMYvJnjQo3vGJ07cVVp4ziiQ0rmjemlXymz/Xcw/yhAjoNlIfnbWSuc4Ou1op
Q+GdfddqDrXE54MKXMmssiaHvzMKFjPNZc/+/UJckUp+R3KBBvyF92PvI0DOEKDE
KGGyWTwPKrLk8EI+Kxicg4IFhxgeLbZvnQndqmqzspsqds4T8cdaeAmrLAKPzLvO
/2Z5IL/JxlcVG6YJu2jYaw1yVYuHeBjPLg9rPBWmEF/LDxA1YeGkHAp7ImO6hsKN
SwA8RE6+mguKpdr5FUau/o+6Q9MyCpsu4LTHfheDoHm8+doWSuSiCcmvZQOeFzFq
kcyywVI6xJ272ogYDHrlawjDSHElR3v2Lz+2qmycq+Q/NAK5HFcPQ1l9uKXOE6O/
F8FX5VurRb1mAdMSoHDWrwo2Ki1dIfXsKnjU2+g3AMMx9OXK+6bY98hCn6eEVqhU
7oA8CjBnDJIj64dkA6MrYoUD2okrHoEIyJQjJMP3c4FemVFVsdYQd6WgysKVl9B1
sdt6Fi+Fg6I2fifsufgJ1Ir52NkE6wW5fXLzrhkx0TIIeL7t4oA8ChwH7d1tDWY4
lEQn21W7ExJejHYvHguCaGoicW0n7MdKXbffP7mNVHT4vn7LDj27j1Takbwg7udV
rhTjtX5Peki0ve8d16pdOspwH8Yk0cTSO6YT2UvMtc6g0Y86/Tl6p/ypV8OtbS5f
dSw+k60s1e+AEIJYaIHAoNwV7KtWAOH2ReChbuGiYyWfOTrQFDqrdG2AXNEFvVy9
6owIukFH1k7jGjQP7BhJ+KVThS3czRA+V/FTeJxd1rZu5OAYn3nu2DiU9MVv3p1g
Rfa5pRM1OFEPT1PFgo6gj5lEUV4LuhzstyHa73cLTLlnSL+uGTnFX5D6ZmFHQDOF
ApTj6nliXPsFJLTdG67n6yFN8Lr2rfffHO7/CrI8ONrOf6rWVmXZC7iLoSbapjWV
dPAL3DGoYtKH15fVqDRVAPFTM3PHcQSU9XL6dFQwATQhTuA9q26mdfUxSq8NZEhg
recvqiyALEgLDfan5DyycyEe2lEPHcJQPT6LGganjyIIJXxeUKBHpYEbJNo44ZKG
/8aicLG/kvBwl41RdUoNVClx9BtsL9Htv9/s9OX0xFJVxB6TLn7A4QyNhaKYadZD
vatOegr5Fpp9X4OkZ/UCdXASkmLLbgtc2K+9uTqas5LBsj5iXHqaPjmdG442jA6D
S2zNlecy59XGy5cN6+JKi3ZAvE7nwz14VN1ydUQyqIFnP9YUWyAN/pJdr2ri4bOh
DXPW4UG0MNfaSabmkFhP03Mbta2K53SXLnZc7Gp2FtMbzh7cbF53oGkP1EsJ0mAb
EHSYgnLqfQg7LLsfWclx3LnA/kD6CJWe5u+jK4k6s4D463L132C0zC6H0hXbgyRU
OK/JC2pUl1hvzwjZeXdjKF9PTfyXo4thcbTIuXIwZu8G3XwrkKUPNK1q8npUpvjA
cEpqAgWTRdT6kv7gLVDL8Tx5AA78ZVMMsnIt9/sv1wF6OMnfUmFuqIQULcjhqR9j
dJI/oHfPK2rwwzwPnUqLrp7MUtvbxOT9cnz6wH6O2vgfzcG2AlNZNP9v15j/jW6Q
9exV87Kz5U4FZeYPVkpiYAgIQvVLY21nN8POwO5jbvkbQKsPySL8Sah9VwLsvPxo
mTY4NSg+X+IgwJEBMDWsKdykc6GV7BBiqHdFccmumZ7N7ZNid+JWjQPCWB1mUB20
JMHCFsyYAIYQzVfAQnuUme/2AZXWlaImfsO+rh9g5gR5B1zwGELxLedChtNNvqzp
yblWfPBJswc61hcMmUp4jiPoP29t4OJG6nMzYFNtV1iqfCzjFy2ugvgnHIPBu+pi
TZXslbWbwGaM/M9I9kxCShezYuguTYncpyaVltha/zzhnd6hdjT6xraYyTUAv6+t
+d/jBNHg2zgntiJF0kJ5xbd9a7JL45dx18B/uK5yDBzAXNubi1dWDS2Kkjet8SbJ
p2xJxJoHZw0gILXt1Rbf7RXS8d1313FElbhEskRGOM2JpNj0z+wW7WS39RluBXBP
uKaduia5evo+2MtJrBq2AfbnbbLFbPUr8n0L5gonNo9o9lzzYZIaw+3ParXO/n34
Pomtd5m9eYxTnxYLmir38e/dHzg8uAtEo9edZJiSOZAceRAXzkfyH6ZX+fWgqtW9
YxUQUTC5hCVvcJMYkeZIlOXkVJSnk8au+3HtEn9sdTUlbpDl55ePY/VETu0J17AL
wmDJdoAUi5ZPGYffLo5U67ratMwv8uQaopbEfb8t7nIMvK9HcCH9T/IP/iWT//N6
msXVNXbyggWrvqQPpyzRh+3G9Jv3huk8PoifXSDbLD3ibN/6Dj9WSBnY1WVbTZG8
qa40dqZCmn94mHrSORDbKxttIT39tqMT/E3lgq5HuYn87z8abQoweHYLPKUDDxSx
w7YRNW9v9stCAo3z7VEDucIPH29GH9myjoK7FieNP1M/+OgPXsghSVoer7TUA3Xs
HYAtWJLr501CEcQD6bSoCLQeeH9XUETIjNMCKoTv895p3w6TugBNcfjTLx20Xc3k
gAShtcELTXVPjNdWTXNnLPC3Z2W/RIoDQ4eXu0oPRsXrhZvfMMO/fQHqPgBRTk2b
qB1aBQ1MQcSnToTIl1aeiM+SR3Ya5fMTfXpfNibkJpz3iRzSRFMxM3Lx1entC2ea
SW0+1fSTzupUy/241CWdcO37KMB1glOIPRIKx0O9BhKL0p07V5qgAs/6GFhI1bdE
CYtLqBszFG6HFntDQr8zFyBbDW0zVyE8FX6sxyqOcjqfdOq+AwqQNKTxUAQ1v1vq
krnrFXIos93qK2hm3QMTNbkpoRXR5P/bNDCgs8yf5TesLoJip1gL7SQrjcvAFRK7
7ePh/7OB8P/YpfvZEaT0XskUkyhsPSGhnJgxqjVS+qTP8gjZOwgMb2G8ka1cjymS
ocUQBzgBq3RTyI53aNvCHM8h1DEN2gVqyoM3PYfeNnNwlCmGSrfepT4mRwio9sS1
+rEj25ZiR6dvN6kHoz38n3/gz2BNy2hbD3Fv2MWonQs3X+NFf7Uvfc8vVETWbGiv
fNUhkkxBxg0JeJhuKM/tm0JOXYz1FVxHTdlpRkXU/19lAXIlHaNCenNPGaTQEZCN
1wwUeRI4i5cZx/CVCsGv4QCF2GRVdA9PwAlEr+IFAjm3bG8HT6NcIWmuqV6+R5Et
GDHC0XvxI3V27Ki8uCXlKAYb0/u12l4vIr8QSKWo+3XyY3b1DiyHKuSp5ik3s4Ts
2o+3eIUtIHtOZMiuDL60MUi1B7n8iKYy4Fj7IdS6ZZ4=
`protect END_PROTECTED
