module	vry_divider(
		input		wire		clk,
		input		wire		rst_n
);





divider_1 divider_1_inst(
	.clock		(),
	.denom		(),
	.numer		(),
	.quotient	(),
	.remain		()
	)


endmodule