`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BTtk1/LNVubuSj/5uNODhXAAXgNuc2UHHXR0EStqJA6BMNoIJ6Jfk0LJ+hTkJxIN
FY4gJ53M2ikRdc37PmcwxYWePRXSKfpysz2SpbiaRSkCItV/TE/ab0Lm/oZbU6c1
iYPwdDdt6M1fmDedsz5cF6zPSnW0njIBWI9tQotC9NTBfk90A21gMwekcF6NQLh5
qQzypJjUvA4OrLbNc+v4fbWmzGs3mmSinjJ5L0zIxuL7tVCdPQxkXTcj+mACLRw0
F3fOPWQgLKPjRm1jLcCXYhPy20X/7Hk/Q7tXg5fnBw0dIpafaNHKskQzyhMKIua4
5PFb4kvuU2qlto5LltAvaiPWvqwH39Be0sm97QwQxqrzRKN+5AO+sWYqfdKhmqO6
61y2G0sf2d7ArqoiL7FBKH5DUppZ89f3NoGbWe4wi3Iax4zgDjaruo3kR/ZNMFCU
T7cK9Up6uWJuq9rVK5aq7br2u9hGO9OXgsM4phMAXH0osn+XfguPvOVoFrDW/72+
td2VFzTFdBoUO7c2SnmPGWPqYMzEkbAzSBO1K4UIJpTDdpF8zBlxnyCmhk7pCo8P
SRx0S/haM4sAK463grb6rvXYflyOGDKETm3EDLgjDah+NPQY0QpuIDWraCc66icA
irnNS4+P7q0PAjvfI565xA4QguJLjDD5LilrvcV/Ook0R543BfIS4iqIwNTM9kac
3oIyFwGMf+mQZmJHYI1bY0cXx10sBwqXoFG4Ryw/Y1V92xJWZDUxDUx+oi1ulGdq
fr8KPQQAm1Ys5umwVSeXfLdj0o168Q0pRGRx6Td4MgTsPG7XmqboGA25igRuOZnI
kw9LeZb09Xe4HGwueW1wJyS/vppd4ReRtsTQdyqDDlfnhf6ZAJWyrXI1bi+1QUjI
HzL8Qcd9L0k+4maeNdy1pGA3u3G3Ty4veOEhAijps94R332BfCcZ7pJlQFFwj0tO
fTk9RVqvd/A0ysRRWEsEbHL0nIDHzLfpCllsay2/q6KjjSP7lq7ITiRji2s64+hJ
DtInS8+eZpz7NTKVhPiV6jxYRWjq/wTGoNCG3p1nXfrtK8crxb5e4xHyURTJYqIP
Gr+wK9ni/0gfkqYOoCQLweturLB5lYTHk10gArQlxiNjjrwOosf+LL4jE4TctiSJ
9tuur/crl4gZoKjxsVBbowEacfHkEok+CrMT9/uZKG1WkY/gE3zUbX61Wi8qZ7RX
lX9Szr4GURz21mVZ89pIdmbCXAOcB/77rThPz0snbZvsCVNlZM0TXshCe9Si7lfV
9L/aJYu4xGUQSNBe7BODY9hUVupBSM6ROHyCEUhsq9OyixwPcDupzA2HDm2uhnzI
QckGKUSd3osl1wo9xXjQubbtumbPuQSWUN/2+aBW42F3+SuUxw3H+PAxssP7Ze6b
YSEzKMVxgzfhAV1/SdkCY54QOppNVOWjMMPLhyIftp4MeNEvUaRCCmjRaLkb002e
mPaLzwg17nTZ3oOUP2yFqCZ8o2oahlaqFqJ3QbNZErnpztltEOkGAR/xCTLn2YeF
dBoIrlj6VYPGX5PaUnCVuWpi2cqf0BCc0Nr183rSi5EDqex9zcZ/qJu3xBrzYIhJ
oSCwcMRkzpq9/F4tNamo4/DFmgJcQYH0ygXbWNMddp50v7Ppghhu4IHnbbjvNVTR
p0DA0sUerGWSKg6ewck3RY9TqcD4DY46KLaxqYlNsADaPaduvUFW7Rk06ny1l7yR
CD/aqm90IB5/CmrsRaIcw//ANNKjHP7mm7wVqw2o0v8gpj84W00qUj2fioqNKRKR
gKDh+vJgU25WhIloVZNqhZs3Gf2DSh7QVivnZJgrK3WYlrltBTGEqt+4ljFsT1P3
jDdafoE2h16z419AHxYoKU5sW4e4/Dm7V0Eo/kfs1PeHLGjtLR5EfrZkIbUk8xfJ
n7jvyUWNN0kSnoG7dDravfWTyrikI7p3fTj+ZyK2nimrDuQFNe/cxsMcOtC1OYai
dsgHMd3otw0m3EOSNju2b3g/xWvZ7/eu8o0eLhXifTW3iZ/jDdQmujHYUcaYsLuL
gDJDoucnwQi23yD/AOFuszQFDm9/UPWHzDJB9mo5sVjsJnEK4yTbWG/y5dEW3Jdu
Ray+zuIqCaEs47hq+m9H1VM9ASPAd8aX3YyfqJyYEnYIS1Xv8tJy8c4tm2iiF3ux
lN8SfGZr8UuLduvKA1aNNBfhPgokN/sF/1dKnS14YGTtDQRTx1+xkYfFn3isXzDp
zLmexD1ivWRGZ1CMH8R1BoaOuWDKgR+n3Rb325FnwedmpDarUZcS2YPx4qJHj3v5
qWbmEtZFRiZ9xDY2gi4C6dMmGFhSKHeN1fjOAlYIzapiFo9i1JMFK4ab6U68vVjY
cLvA50llKGXpVSXD2yb57tQOaT3AU+tHnjqRUIfkpZYI0qtT/a4cUDzAQMOfY7pL
4RZtq9VAmwBj+RCWtWF2MYxmGwy0gtyXSbUrrBxbcBIM21KP6iwU5ihnE2GhgeVm
5tpVLHGcZECUSYO1U98wNAfhIs+S6QBlmt9GYcHBmAKVgu7XpnDnfT6IPDRrfIua
T8keXFB/qEr4GX6jlnbnjaZkjeHpe+XuR+OVmsEH4QKs+ir013rfn/verUFbiWYZ
YbD2b2dy6Xwe2DyqWMDfioGxZEMhxdbaegPWhgqOr9zCJd4IQR4gt4AVy2kvv2+H
x4VLUgEEDnGZ5EBODvZfA+mFX9aAfHEvjK9iap5iA8sv5Uw6DwOpLVJgzGWj9Gzy
MPvhxPB9sLBeCHn5APwvcciHmwKQwRS0bTBVmNZ3Crv5ufkp5kHaaT5N1ege0AP1
5b+Mq0EvUbE+oIl9ESVu2IkHL84fLQClTIB0vUZdDYxM5ZsE2h2fsLMCzxMdmCrC
bT6FQ0f5kNVrg1ldhUOvzulOjs2+j7EkaNwc+sVDBgl+FM1C0ao6D+k7DqPxeuOk
4+vvQZO/dZfz0OCFUbsfqzS6Wt7yFFfN5si1vivf4hBD2AzSilXJ+GG/H3xpGgWB
fOyXCWGq2Fz0aVXEgv0kZuwfboJ6SDpqs/FM5ELJJhjw2fZCMbgMQVaqGutHG5nZ
Bf31w9taNjBsL+2/TILNps3bubuY//Qn17UhlZ+4zrERNP0slshbwmrnsPWB8Hdb
D2rpkmr0y6XiIRL48KVD6+fJfAjH98QoGL15mKhG9rDMdZ3i+zNVhItoq75zvAFa
IWDads7u6feBbUq+LOwEhebx7jUvuU967nXDdFP5xFDf83XzwSA6P8lftjWtPAFK
4E5TAnCww0yovKfQ7RVs+6sPfy44gyFpIo93ipn2v80OXfBcYOBqLCWSiP/rHvZP
ldXZeeSCxYIgO3XqWY2xurDcX5EVdfzSD+L+ynVTzvaKzV+tcIEsurlByTDRNDw/
sqEzri7/NC6s2oFenrbecqh5zVOaEWPels37uP1leuliPExFVsZs/3WoVfHNqHhi
TnvMUhf/5sO3+gEvi4Uq+QGasE4/OTDNATvuwX1gaOWP0I6/3oURJICv22Y3SFHd
zky3DyHyyLWhgp3YlL7Zi9Z40ce8uB/npzWZIyu14ZkHKHvD7Iv2jy+gb+y7sZcT
jNJXjx1SWzFsjpjpl5LGU7igRyeLM3enWop+q1FoFscWtPcK3hud2WRUMGV5Scau
YaJLV5o1Feqsmdnk3i9jDv+mega6askj9dLtafiN1AFX11e9poC9JVsqkzTnwUhg
X3vkv+n+D9okaUlWCIwqfCi768XFof+85sce7pttslHkVBlabkQ/ncEy+5wi1BYM
/JfeIPJNsi0jctmK945IGYLv1RLhVyz386e6VjoWSsXBJfytRbKmcr4R4btdrjWS
yi7r+uLFNmDumObEYBYXPATBFRUfdxyBg5zg24pejO6YfDiya9fy+YcFquW9lRny
0Gt0K5FfJhjDiFB0bjGQe4ogP1ISzL56xnnrx3QIFOh/OUhU/vtFBdAXUBITJQQx
Ak++RD8dbJcPOu6OAUbPIeKS3WJ1O2lE0qMSGfGbN12RbvaQ+xMc5Zl/KLYfrzF/
lFxjiqEMjiWZgQf4zOrEVe1hQx2poFV0T20zk3NMvq3gKjD9VcX/09knX1jX8SEB
p9MonBh9uMtJor43dZ8xCVZtuTAlcF/MijIiqAHFKTVb7dYAdiyFmqL0XZSpQ+7K
H3/NkxTGhjEQscYRbJcSMr/9k3Q/kkLP3c1+OGAvTLJmN/FWcLXXRUk0K1WFk+c4
RgqRWUuQ/rLugKGjPzIjvB+MqZIlAL0lJ6uhbJcz62+nFJTjPMtyGK2XaDr/JpE/
ZqFn7y2J8cmWtCePk4h+2HVblx6x271aTzcLAnd41fdEWeW36ISH17S1KsU4bM5l
sRkYYMMr7ut9Kkrrw8He7dcpXqdEQjfsyo8YA47vNhT8nmqpW26tBWYLeix5q0uO
1qp2PY4ApJEDbgi6xYvaV6GbfQ18SWU3KzDzdAPJe+h+QEyhhgoYTYdzoMYcBJii
asoR0Mn4kkUwjv8qQWiesvP9P97V3WthV92TNe77dc9BKpQyJehyEG59YVhV4HRj
cAA6VvHegIHYrYYNSG0/D0dUgyPju4MR4uf7V1Zv2EeOI24b1YmbIlH3OUyhugjp
0OnBZxGOY/iQUrZri8t43Roml2jxkAPlKkvshqq1mZejxz8dLf3ttjLiT5xQcKyy
GZh6dSnH8vPVR8nTxwYThRd87SdJS4VbK8LHi8lh1Znz5j3qUU+GQb9+iR4/ClsS
2jk1diinaEaKgyBIxxSTBvTnDGEbdJ4hQ0MxXjUEJosHxb3e0g1W8xfhrq24iPHr
7QRqCZvlOoydZQR8aZ8WAZ/OaIMdqCnXP7MOkH0gkzpeDSngkAIVNZk1b0IUQUHh
dljjPg9hsrLBWhdinbIvzZujZxg1kyJIqNd6XfznSzGyhdy/9KSn1DgG+qsfLu6C
Z69s9cZvukSzjDvj8zooUxS7bA9pkEdWPb0lMuvtfTtEi1m9vbzgAYOqGNGZ0l/M
LyCOjXg5gintIuoubNe6ufPaETUg/6xJHR8lItrKWngOIUwsCnukVVhEYPU2TNlg
ugS/N3PrOIN7WFXmPKBnZGkXlsthDG1YI9DGM5fRbJv9vu+kDtOWn8d2GnUbLSvZ
5rmduAVwf/rqgMrXB2LpS6ZjaXI7Z9pgye21NEcLKHYBgGQR27zAGda3ycRykNeS
Hewe6mdWHzQuQvSIt82Qg5dYKMpZkWhG/sur2T1U3YsCmhNKwB2TBlyeU9KvesvC
2wh8D5NcVrzp+olVt1CC1XHhFQ9FETzYVk7PjvnwSrCKOtjtzVB/gTJSbKh+TFc3
hfST9Z+WdZMaZmwhl3oRIfctQ8sYh9IyB1qrA4PRLC1tzmldiRhmWQMZh6JCEO5Z
e0Zcp9JyuqI+flvN08i/7os2FzfIyfBFa73wib/OfFcH59uaHrvdPADcpAkEJh/t
LO8n4qoYCYQQ20sMEyFnU/8NnBO/U3Dv+8himMoXe2Gp4M1nmPQrmSeLjv0x6A6N
NQ9L3pkL2OqkafoU/dfeueq7GSs4n86qXLZkXpGNwuKMWG1uJAaPrjSMuUFjEe0j
15pIKdr4vv7aqGt/PMOuo2gVbQi08uRgAJfr7YKotY/Ga6J4MqjRU5IuTzg2uCeF
20yye5MDNgP4uzozltKEp3vrHpcQ3W0e2ndp+sRw9OB5ysIltoGgMl9qmPxwbSMi
oUjALLOZspkF3v48eW7Rjrl5TkWOe+1xmRRP8nTMjvVMncK6y4kQVpzctcWZvXAo
ZorDePwBy8V7a4z52GUfGTqePsli9WHY9Xq7Oqma6RWf9cuNV+MqwffB1Grv+hAb
ypQpVGP/a61Yoq4hFcBIQ/u7qEP3azIeyBwulBkW8nB6bWFbaYJUMuGCo/dtsZHv
MDl6PtzLNwv7V1PMGeu9Qte8b+CldhgT7mZncMNEoj+D5DUrlMkQrezVBAZjwlAH
dkN46oTSweAeqIYUQSwqj5R/upeq7O5RxH3b63SSg1wRix3NYspgKvnaDThaxcMU
1DrpPnr6pjem8dX5yYvjPrdbbnFTde+aju+kkZqICZO0OPe1k5KgKvGHT1eO0fZ8
Wp1hRdqdOTH5PZvkT9gmJAwPYoyv2bmjltlywEUGuJHFM2jEQtVAhtPWhJGrcP2W
qcnw8t8qGfe/9MURN8e0OB2GMd5WpUpYjyDF6L3TwpKVTR+IJLC94d57UECOwipj
oMF18JwH+wc7mzf90D0Fjlzg2T2IVIAcF2TII9+hVieQ/YzPv6+JyeOsrHikqHiy
SqKHckdPjQUJ31tEcnGjCMI2JcBBzHqcygnqe9Th4FdVzjmP4mqL8jETdv+vNARs
dHONb24nMkt3hCFOmLz+oL1pdkS9j3CkGsX+gfc0PPgi3MNFS/cw5UWN0d6IoTbE
rZEeBLiOuy7NkRRNYVfhuzhTz7tYzLMyCaqdtxRxP3s+Mqem7qIls9WO7yy+jiK4
mTwB2tWsSVa/1YHd7OBf3iNs5KMNIQVtal8SAya2hpjfkcEgHLgCTwmmEUDXOOjc
T/DdbeQa3k06OvMpgXqJFO2wgimOJ9vfDUWBU8oAkDs8sLncJGl6ObxIpxKBMl6x
G/1qoWkLgSN0y1xz5Abc0nyY4DDHSDDoNLjnznOz9ri7wQOtHfK0RW2D89tBjy3J
ODsVhXx59ePytLyAnwFfVcg1Rd77Xwd+zDcUA8IGAgFS5C0tdH4Y7TjWhjGFHgC0
4XUWuyiqVY5ZHD0rIJDqrsCi9WAsZdcuoe1edHmdyV537R5qMRDtpNaHmX8/sez6
qlgDDN10o0TUKTaumMeWg6RLQJza7Il7FmcVDsApx/GVUzAP8/t2odg/hcbKM3dy
1r94JjzlMydskFrmAEDrDguugSA3v6cG56tDOSLu6dH21LIBYx25Fv7SJlLRJDWv
KbsxSAeLOMKVNVaIkFqq7IYlCY5XRaEnJlhyjNYAB9QMiQ9+2JnzQDYUPquImJOI
erdSBHHYJPbFVCkrKa+MQ9x2X0ounPW4hO3FXrj2jH41qa+zAJYLNbDdV+cQ9qf6
kyXmC6GxL0CRUM6I0YEYG12+q3NZwGI3ndwF1eLL+JDgmMK7mKDyeGTFsxKYazom
lthIZpwqBdTCkeDvplPRwzhpJvC7Gi7fu7txcBw/yVUqMp1dF1KGcCmvRc5qveHC
+fuu7H3+XNofpl9vXiSgZh5U5nkiE+ZE+MhoMoDTf93+fQBo/UxVfS9lQ07/7aeS
znTwyETK1xxzg2i9pJMQPMmIP3Y7P/rik77gI/BMHZBHoYlgft2tY1XflFcZrOv0
UA9xIUZ9Z11FxGA5kE83i38xNkJ8xFXk+FDybIMDyYpucc6vQJbsS9Ro1a414a9h
69wxV9nq+hv0YR41vD7i6zIffbbMVmpVKGg84WsQl2tnCAg5n/zJ40BWkIbGM4Cr
HQmUudvTACE5ZrcpJT6KvlNby1nLVzLZ4q1UeURghOkKaorTQpD3sPJ2YCAIl6nc
g0Rp+EnhLWh1D+PHNOaSOsJJEG5lGX/9HBbbv82WRfCrUxzzfsCtC6buqQnATnGT
iHLyP9k5VenEZ1pqmOFf0Pz0FTp/9kB6Vuk5+967cVlTPe1eD/uScfpdLibJwxG3
Se/nPoZPjLS0+allicdpcCQmAu1McMWk9A8uPkYx4pv0PvNtN+xyjnkBMqwJHfKE
tSUzoDYX2Anbw/EiEhBoXB5LYhfg8xtmB1jdMqmjIGiW+2w+sSiA3LwwVZB1fjcC
dTW8szO2xrxXrfzwEJuC2FnNp0vRWJSpmiFa6zP7JfGRV6qDEjbGUEYYAjMkhXYG
OTqpR2P3keRXvJCIA2McCXEpPYt27BNhtHjULcCDxxohGAHaaSZwgHZ6wve6SgcC
ecFxn6fX7yVA+Tn3brVw0t87z4RiaCSxVJEP1R00/tLXpecerEGRBoKcP3slLtiw
a+93eIEa6qRzldHmX9kZSJhI4U9jBhs9atCPmHAHzlSCXjJ/CAcx2wl3qx4qZaz2
/mjOBlY46Pbhd5tzASv2bq2QWeMb3nVRkyhEnGniMMTxC0Am2qvZ8oHwM7AD60Z+
niAAv11vF3QZaaLB9s30K9YD6ezb/7V3nRZpZkpa9bEdLbbig8zOgQcw0rBu5qpZ
8b8kG1/nOZeetMkPjqtE6punds6GbNY1UNo7SPajJ60dcCzQ/VppHfxT/1TeN6uS
NYpZmS06Xfva9xITYEIYefDx3vrHBMdxQwZPCLfYLxyoqxnCjAnnDciop4OgQqEh
M/Xqr0TC839Wl/7TPkdQ7HMUzRLdKqRLkfYT96SmzQT9UQP/E077zSUMJJ+EUu9k
JkQ2DQ7iqnnzkCuEDK6HVLIhrIKBVxTIyHocJI4MMc8NDr+UkIqmEb93Gqnr27jV
hH0+mx6x4jtO8EuHFjNyWowIOZCmRKbzJ0x8ZosiyBaFpQEfKVB/B9sy7StyE2fh
erQMrkBtBeOmnp/QrNt44HArojsj5FoEV35X6LoYuZqQXeStajFoRVGYxEcsRrpO
sYv49IZB1reSL9qtedek+nyVb7V+JY/MElOdJxHNV7xe/U3HhWeSeupek4jpSOha
cXjLaiPAi7Huqulyng9txNJksmIdx1UEvYOT6yZ1o1hR+Ya4+7a5LhXsVNNPGB0D
zTeCEG6MkM7kESfAUXqtCS9p9w6uWkEB6aOpU1gisOIKXTS0JZPea5JjFk2AakS3
dkUWksXyTK+MnHpkDO9O35cNtOc+03eGZ3AA47Solh8HGJtJdlakhyiLHjVQrd/k
YEvtuX/3x6MM8wlE4DTXSqCdIRwvlTXhV8XmiBzGA8P3hBubGNSruoKkDglr2eSU
FrzRQlDepohHD3t5FMMJM5CfnFyVyh01cxDrOebD8pQcMxZc+xEjaYu/tsch5OOn
JOPc0fP+m7lCUFTLGAQuMKkhOHOE8xY6HB17SR5YBn6dJKyPaXDpJsVqEUA7tWx0
v3HRHu5nn4TQzyNE2yA1TUMgFoKg9IDQa594seqBgcQ+eY8xaFjSF12lEvT9egG3
7CY+AZw6FeY7xbiwCkvFzhcFxDpTutmWV9Y9/RpwVa6ubRx07Wg/vDQi6GfrwX3o
n9bk5EGcJ6gvzouJaVHDfm1N3bdkx/bz+4li0xa3GmJMwWxpK5YNendo1fWSUGzp
uP6jiGXLQiKVDi58aOVG+LRR3+/L0ctEG8U+beSTb527i63fFBCGCuQAjWBprkCR
JlVkRZi7z5vPGxXuR+ZN+FdA6WZmEP1kOEiVGRAxlmYkg6aRERYRxxV40M50bNfu
peiseP9DGZ4sIsLspwDnCCjQqUKSJQdEdS9S1zGqZCiBjcloYE1khb7wKwkc3Lv/
i2fVjOCQuRFvdHAbRylhXPZRIeLYteNe0UdZ/NoTEMfoTKHs1mV89gQXGdSZFthe
N8S++w9C2NbhkPem9xZRd1dn1mHsJfdFNuPvow98xc1ASDu6HKHl3erwc8AyZ2rd
xsq0551mwmKG1TT2WfLc2RAtWjFyYXYoHjDflTNO5s/MpBeL9AjJexuJB96QnWxe
gige9CUTMeWiWr3NkkO9WYIUsEPMYFEtMZHd4FX81WXeHwPIkLWpqWod6pdr2IpJ
lzaPY7w6lVAqrgmJfvej2nhAyhiy96oeBFve0+TfhJZcOSQThva8gLAHlOMsADLO
/BgZDrCnd6jzSReVNkNkgAXI8dL3/PcQT2QPj7E5sJRL8V+Ascu3KXhYvWaj6kcw
aK5yk32c04YIx0hx18Xs6auPVk8kVP7TcCtN6uZLk+GiCGSIcD69SfdM4kZZxCJj
/6BaI3hOsNKKU0zK/pdaCfTVA1RsC22C7zDhWp+HiuUNQCsI2wok1JUM1kG1r3JO
6rCvhu5KnMAeMZkKZzccMiRgjtJKdDnVU1iIkVdPBu2fW1yZNkxfzynQ7JLeOnR2
lx8t56/lbq3LKokl6BC+0IdxAlKLesssMs+QmV6jf4y7XWQOepk2poU1G27OdOPp
/p5ugXbaGeFD3ZrVRwNIoscfvdDns6faxGfG3pXWmvj163YG9A34wojN4kQh5Plw
EsFRwJ2GWhfjINrmhp7nNXOFvD1YhHMpEc81SKz+J+HxpbhcHoUwEuNit67RIAgE
Ey/FuTAttSrNxzA7vRYvCD3hFE1SkWEoztdiEyM9oGc9z6WfgLsrq3wNBH0tMyVS
SNaIwSwtLYp3gy8jxxwWDmWiFY+QuChaskfd+1vMlHpXVdg1omSxsHSfb6P+7QZM
VbaRWfo4gVADEvpSFnv1UQa8kHyaOejGenSV/WpUGrLzGXdaxAZsE25Nm7Dh06Kn
bawpUQxQuRxP7uXj0+6h5/0wY3UqBk3r1ph/egq6sSbpzs1rtmC/6HbqUl+0GPeD
o2JegcW0NMj9mWl8uD0bR332mhadTsmu5Mn/6VM6XhdO1aL5EO6x1cflWjw+NJyp
1kuBFnaXyBxkZhliZhFzGwvVJgaN/in8hDszjTK8ybjOoQGaQcgMZHVkWB6lcEff
XHFkHjXqeryI/If8PTHhAxk2mDFaxbx9qA8g6nYjF8sEDh2SV5kGl5pBwr6UtTeV
CmplrwMxHRv06nqbSb0xMSDJxDcH1fYM86Zb/wrm/eNa0/api4dFhR0VyNoiINda
F8t+eIjZ9dpVNPUOt0nWubYe7fzpRgIUcmt9hT3t4H+/gjiDCybGFPzOygju8duK
oJMHsiwbjYx3GsQbhMlQZXgAeuHH09h2aaBz1z4suHb2yM5Yhl58gsxW/zLYM3FI
BIyh1ZN9aR0sXS7IOaE7g2t9q2kFjSn0y4QRYY4ZigQOsNZLiQ4K9Q60AlaCOKU9
JROXSE7GIKucrPIJaK+3yIWKRsZhP6jpuot1/rBLxxuhCQuUU4XsKID618YKd4UK
FC55dapKPf1oTXvCgvJ+q9rKjg7nU9elTxLaKOMIc25pXBgqUylAv7m8il8gCPYn
ZFcWHx/+8DbpSvIe9RkY09PzvKxn+2qVnk5s1W/Ap211UveNvO1GhTRVneNJpKkI
lDITke4cKvxKRrGao8MyBEMSzKPJNwFVw6dPJupn/Xi1m8nXaZmOGjqcheurSfm6
P9g2864jWmDALI2XwEqrWr4Ll1wI0aqX+idTmnpwCK8KOZn0S+PEcs07jVgUwNNX
wceHs3Ld5NBdTdOEuXQrC1KRWdHyWErI1e5jVAkuKez9vlK/QVcLDuO+yoW4RjKI
SPIKGmM+XygAvoSTbIQNhI/TGGoahskr7ITqr2EDIg+ZpAGgbPux9eGgkpTDYpt1
MEs7JTD4aYKUUi+VDz6hIhESAknLxkmfOSx038hW41iTdgmqw4WVf8LZHB6v+hx7
6YbEBzpAtAvPvB0vsGL4i3E4aM19OBa/hXangWuWDbSRHHx1is4AaHrwld7ONtEj
4G3BxDKWrmJZrHo6CR+P6m5PCQcrEtRCzpW/a9vtos05gk40MLR+03a006Ls7/T/
VJ35e8qd/uMYqhj404NOX5mJ416yHSR8qKjuYeL/mVaqr5LfALpeSnMztoHsQv3F
I97WghlLHiPQWAe0TxPI9AEpf4ySDPF+Hr7qA32bAXCx1b4NApV9g1xWPWzxp/s9
2EzJDS5ervthRMSNZYvAgflCpkRQDa/pdd7jZTUj4lHwIlgaZB9cDlM1hD93ayDw
G+XXoaoAYEPF4zpg4XLDoWsRGbFizvly+bNa3jBSArHTjx7N1yQkLMFcsDuptpjw
MLfqnLnQovW4kJBc7avp3aAu4eHX9er953VffV/5SSNlXwEnoph3ncIgiwnle3FB
gcnH5D+FPR8pra69ZkcLkRwhCuZionCBE79cvwbLH3pUu9ZDeyIUpx4c8i0xutmM
sqxchkpuZ8frda9SBrJM/CmVjvOHza9h5dHlwsyIpQnPYk5I+CRPDDJhnz3bTFaT
QROyWfXSpqyFxSNOsNZ41O66Qe1GRMiEo0BEUERVPZNhVgjsi+F/plIItAXKqkSe
4tRYHja6UpZCDYB494wbaMHetSxQddeFyhIWu8Na+F2SdLIk7TgbsypzgDvNYibK
66RXtukL1YOFd0KW4SxGwZDkf6I5GStaRyh1uIPo+jNfgkINIREJcGwkJHpV26/R
AHplAh4QPmgGHHB/huOI4ch2Etjd24wS64rxAxzTVH+Ieoh/YkAgeQsx+KrapeNQ
PA75FwLu7r+ugVMafMmX/xrnynthlmrtw97270HhiDtievfYqU5m1mkV5yTThNUa
xa4ifFOjBVnNBnnPFI3L/HbmQqgnAewgwAeeLT1l8j/D4KuTz5dGggM88D77fWHM
7uJPTojH5J0jl9QcRVfHrmA0EqsWoCYrIbmNBDGGV4bU0Ja7bMbJ7wzUuGckidk6
0c2THXayyIDnMcC6BxmWIMeo9wEqx9KIHfJg/xvEFVEBkt59ydZnTQpad+HtmDQZ
6PwB10bOzA0yeES+LMg88nkqhgHbDv3rbgJY5epVdrVKrdLQRNawYWbIvGRcZMOP
YbInHfg6GG1Vlt/dQ9GtEzXqSJVWs37WjDz5msT+YuY/YQZnfyXc9Onp0ZqYQ7Tm
cTPRseC85a5BbsJ0boRIcAor5z41UXAlcpwTFP39nGoD79woqXgL9vAVAzaGQpbw
P0xdOY2aQ8JV4I/WVNt2cnZb207Q4mp2m/CsEuwWcWrTFp75FpR7tzMQxQ7i8QXF
ly7hRSeOEYGouCspNK/WTevNskqMU6IE2jV7Wg2/4JwLNbmw/JS4qAYqa/nWM9+W
tiPhpGWRiI7f2o6rRe7ngF91Pgk6vqW0IjzBJgucyN0oUvcKHbVCIyFkOVQOSrX5
6SiWRZvMiYff9/hGPDcbtLTAtjkClShhYS2K8HpVBbX5HDk9DcFhjrwnJUqf3t16
2P+WJW5Vr01F5WU9aVtMJmb94iSbTTSfPk4a+dUntYca9+IdJ70/CtfnUSYu55GY
jQRptaadvrnxVvOIXNpvG/rMY8mHzATjDCpSEj3KFBNUaIw1XC57lEpehwbYxVOw
emenWHwEaBvyEzuvVNLeh5SFmHTy4ZrpxL721kO1VEvTqGCt+xNi7xYBUd0JOj27
MkJ6TviOFVtJ5HC79+uVe9m12+A9sjK3SSi6YsuIIzWx4o2LJ7beNHcL3fQ9JFlv
9FXax1F8WbGeSH6peYVmvMGb8xaHSoEluNbZdJhBvZ5NKnOr9y+otk2tcDsnwdOd
3uiXe4KaErL+8Mtc5PqE0w/JxGM2jsCmby90xP8fUfYnLyXxVwPZfGmpX0w8dbdU
`protect END_PROTECTED
