`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tNHrVaknvPKI9FQAB7o3WqRZQ2Ck/V5O36d9Skuc0IsVk0FqIvOpinpdUgCvIIx/
hD+3u9XLvMKy2pOQ8JHJwsiD6pZAmHQveFm+Uu9b1vclVYy0z4QtiBwbU8FmoqJs
qwNvI47G83o2TkZK0SSERkRGiHLsVRFb+BA2CMBfzdtybtQtTnz4RQwKuDgfkZyd
KKpdjGg4iaJhWqVzVFdhHDR8y0vP03RyjLbKzWen3YYmIkLWBscQ4IPUiv0U00Rk
IO1/Tf6VxTY02patfFrjK7iCB3esEEss6f8ItaupBLtP0H6SB/U1JxtWDY2EyMAe
RryG4ZYk2RIURhBGdSDGrQSQP1W2aBS4P6aa5unprcwjVWm5vSNvgAluTR8e1YKM
9sntBP8hnI4bCI6/G+OQk+VMtLQFDpox5uQnFck2cQvcePXg0LIPeNQ1GDgdJSZg
NIqkbr9wUMyEC5tH8fWhtQnTC/lA0PVtVn7zILN+Y1rYEv6kGzDNkWQwiqo+LfYY
bzfaf3Oxk9lJ7RJWvaUEcH7cEXKEirtVUmMCvJfskcZ7WTgLxqZRDrFJG18ERtpv
BU4AndDGOR9MIQLtlgDEBUK3MqMYH1sIYVgf+DjcTkhScVuZI7mthTi59E+ox9hU
FmUVEt3KzL6PXHLDBaXZPToxMYVSd20rwnRa1tYI4YibiEtMI2PidAwRhKQdYldR
i2LZ8kV9d1OBWQRNbYTRlTX08fe/amKKGD/UvzGqjBnqtJRpE1EoshJaur9Hsfp1
63/gn4NFoh4WkAzqfyR1voHHY836RoYqF2nrmWCj5CmJWd4a6EuqrQyn1QF4SjHS
Oj9rTdDhPsTaKocNotWJW8ldWWAvgnN5LTqDe4M9PIQ8AAjGTiRj4NSwzrSPf5m2
cVltFXzHB5vJKKUOWtmveEPDJRn00X9vWrn3os5rgNNPDfmu/OK+Rm4DVpw5I9Ww
RnaJnbCR4vAVu6sgzjfqjqVNU0VCY/sDFmyAn6ti6nmQqTgr/lYjX7agmbted7Or
ScRMQ4EcJuwJOwpYU0kPdbU7uW7xtornypKNSm/gbQ8/NPkLYtAp9yBqBr+Q6IQw
wcq2nKDVSC3ZGLYAcSpgsrFE3P8rQa5wzmbXuCBaQme1wVIvY7zXTK+MSp5t4/kt
Tz0z+/sENQsO+ddGKaadF3A73MRd3FgS+1+fx8ZJswM5ya2to6WUfotmWEqv9fWl
Oy0Q9ati2ky4VHKvF/LoTJw7b0OurrK1t4gHpnVc6mD4KgIjP4S6+60IplwIHfd5
DL1B2B0uuy38PyVu0nQaQuigutuSeFQQMRLQEodMjRTcdQcpJRq/GLJHdUvGPLYS
YIrkibl3Q9agmMYkQPg1i3NYSJ3MIMgrfo6to6OPUA2c96I0Se+6OfUq1fECpOqK
sbqTi2imB6OuTCoHDw9U0b3spItTOR44+7X7VnTAPBy5iyKyQqeapadu7DCxSOOR
o+KtTmjuSVqiDAJzUX/1tPfejQnHX4z4zLyrygaMtbSF/04mHFJIsX5bX6qhQTyP
PMTKV+VguLphy79A8YgJjQhGL/AGYHLpwxhwoC6a0sBmZ6RWE7tAYdxQSSvDvWbq
FBTZUcfxu2iJ1CnZybgecIwAl+ZGbTzQeOGC3T63d2xyMkJizDyPHhcf76Cs1+UP
om01FhFeUlqOroQc4jreKCAQTh3u9vGHt9jKY3sg7CtGvmRYBy2HBCGGQ2LQRfCc
m2N53fzY8bKZ0afIy0IdTaxUUEU1kE09Jc72VV2+FFXDHN53QH4BLkEmxB0sir9Q
qq8xYE2LYC2xBB4mwM9EOA2b4GUDKfuGcYXeFgCTZIv2ejttOSQZYvkXUJx294X3
ijVRrpULo7uthqEVCCtywVSuFEZxNDLMQhiT2zTCly5jxq0Ho2wvFYAgM+gF1k6V
xx44B4aL645FRwNJpgXqB4vwkUYYEbHBxE2t5eFEEt+LcQ65QLxop4OMxIm27Ava
0oebg9w/UecGdFiZrbXu+X2wbFfoVye/boLW7m6SXOBJWylgkFiV6ZnjwKu9V/Np
itXq07o1zdFI4Db9h95LSOzaGZNDua+zKOR1myEPaiSj4bssh+TUUxrzZ0O9zI4Y
jqZEQcpyp94XlM+1WZ7QGYvNcCIWW8sLdPTdtRDoz8KToK0Z+uGAoCDlExKEkbyp
Kvc5mZkkSswOMbxwYXkL7Woqd+Um4WKSbDfZnbl2q5FuTGOTBAnWha+MEogzrBc/
GcX/rf4pJXCwBr/IQeniM3fRyhDN9VisP8kaWlOadaxAHZy7AgiG8394RTtwW/bP
ls9p7YuU0anVVV2WXfhzDIGq/jg/9VRHdT+0PPiOrekwR56RVQZg398mkgFujevo
c8ZkwJw/SQtP+UJBW/AqiOeTYKGLidjxisW6swfp6AKkXO0A5GgUNxkX2sYBLvxS
tN9IXLlq7U4kMRjAjfyS03NCmWbEPjthi5H9Pqh8VOWtsvFET4w3918VBYmfA7dh
bkTM1Qh1azhAd6gCGt4DYuJZXfPhuJMho3do/U8giZ2cg1ItysAmWLdq+ceqkRvH
Oc7s4zO0tXixj4ySdXt+RKpYYgLop5gLbYtq4MHBy18BMyDyzczCTrZ6+t3XnqX5
uj0VdcxpuutjCbCg15hsSa5w3W4wlo2Xbevo1OHReVIyC7XNBPvn8ojRLYTpFMJd
MbJTMX2G/quP49GH8cMQp4+sLiDkxzYCMLiInjzyHkVnjYZrP7uXa8s7gqVsSy3l
mxe/DnPQ36I/AGpm9788wVgcTMXtV4+X9x/joiyK6qS4A5z130knS9/h0ReH6BvG
nNEzC4BRmwqo5/tsma+9vUb2BLvEHqMnUS8qprTqsm8qrjeoDfsXM+HVppFyBzXi
8b7PLR38Rp+Kk26Gjcx0wQyZcs2mhUMCRDgMVF03zEE77OgMRwBryi4lIrLfe9E3
6WNT7znmOUspBnG0f1+gz9EsZ8ysqS27v/ZP24bmKbjrYzHHH7XIsoJ319QzlKOz
h+DxGQ2lb+DScBHRpyA+4EfNmwHlxmYyKGbiC814lBw5zEFIJM9QivzWEtbFe2T8
M3f4vt9CLPjzthh+fZuD4KWkI+gDLjIemR2GTABZK6VpsMA063BUn+ul/eFQPGOU
t/e+d1wp0JzDJ6ovdAQCga9W3sMGmSnQ0h1BHa5l2HdoZ/9rW0uAIoKKrpromZwO
gd/5N0E5s9juAnmF+v78Bj7No4xaWA+rzjpZc255t2ls7pFmezX4fMOJqXeKYkPX
KA/Da8jy5U43V4yadTRlbQrmykHAC+g34T3s0wjNS9wdGTDh7MHLuIJh2VKdk6QQ
lTYRHL//Atk+pS1v4KQFUidKDhW+x4z1kRsxPEWVkWtzDDoJndjGF4JkyoeUOVLM
kjG58qQ2FvONCxPOCvjJGYbRZnVr0FYL7v8VRRcioKf0R9wpuGXszMr8RBU0WY8/
v2EMiiSpSAfXqIeaE2FfSeN5ay/7baCKmd9CgMUy53SqXIi1ZfPw0TzN0M0n2qyX
4oh9RAXfPmYYMhYY0sWw7WiZLlCOoJSonEZCHJbfOYD9UiBGKoeEj3MJDnpjW5Ks
BCJMwd3s3vYaqrkOhAWfeenKu1FLAaH8Dwaf1vPwjgMKxlDNaLd6IvNLEEbzhZnp
CfYgSC9l4KQEJ+lot49Ims8EeXrtLzpAMKUVC1gJFyxvzlI3G4PsAnUEj0T0KSOH
/Doc3D0Kl/3sbmSflE07AIK5OkZJXm95N13R7zIIUfNNMQL8CAO0a2ZH6i/b+2Tk
iwMQn5lTgSOZeHdGLbqDkUdOd0fu/DpOVPnOj1Bpfdk/7czrDuQD1HPrT+1IbcuA
3hAleSxZ/L5n0NBWFN+5DcnKz+4dRCkuoJS6uaxKvq89f96cz4qPf6TR8EJokWLu
vdUKpjV2WJxBDQj4jfWKm8X80WzrYPMWrosWTfQtizRVOEzpTMRHPpTGAsUYsK5T
pyKwiTZN5K4/Itl/0ibjj2qVN+aI6Umh9FUGg8GpP5iZ+yuePrNqrfWC6l5FasnG
1fmtF1Q9q4/LYSsob9vgNLqXZran4zDQE64ZWkBU799AXddfOjKSEn6ptfSnjke7
argaakaGrEUmkgA9Oa2UMZxRxgrTCoO9S59Zt0PridNNivI09yOjRa36yQH15gL/
BY93O76Z5yVBijbD0z3eVbCFtNmu4pM0LOWa7rfNpoumQJHAN9ZttkWdqKGFAYCp
suuIJ7/GkZz45crXPqjScrxV09TVsUzLaRHdoq/sT8tn3eiFgeqx9N7BWEHLWIuy
a9uB1lQLxxr1kS2FGbxGbuTlb4QyzyedA25Elr8IKAzaTfFsORvV1UdZ9oF0uYjs
CcDM3JPPZigpjCAgv8AZrg3J/+EVCBhrgzwCmJUD9j919RxQ7vZ0tqy1o4dL6kgu
1YE8Zcz/gvmhXTP6Q78bsEZJHMNotda6/iro5QUSsoEUhi4ZCwkrpiotqjBHzU72
V5Y8ZxDJiqIlNDRTlR4di9yO/o1HmA/oilrEOVD2im0YT4ivfjpswVQy2mMlXzVl
XltsnWg+VUp6lYeRDxz7Xu7ngYJAARvc7DXV9CyEkIoPNd3wWi9OEsubvqRbFB53
bn5T+UhpoOc6GuX8OlhscElysjHuWmLE+fvoulIE/N6o7tvMR0skdSaPp1UFTSy8
HoHNfMRydCUx2i1kUv00nST0JxSFftSCBElOSmBD3uD3o6c+L1myO7R8hJ/8srIm
M7D3Y3gF24v1zxfQw1d7y6uTcrs7sORsBUs+x+1xW9vFA7e4wqVtLC0jumTYZyH/
umstYukjAUIRALaG44hZAhxHNESwcAyynFRylkPTHyUzdd8zwUn/RVmiaPp+H06u
ooSzWVgRSDMhao5JCL4IDdHeKyKW8cimc9nD0ovwFOCSECS69T/9ga+wJvV3WkeF
53SGhgQeb78eDH5wY4uDzlzny6V5pqF8/ZdtE47/XT++5izT1l8z5WTpm2OkAj2o
fxZoZYeTzpiR+GPCUZ7GYuP4AqlJ3pdsu4ao3NxX8JiE0deLIyuOY13huw3Dd5Xe
YDhzojhrsH/frTilUYe/ePFV6pknozGsc0CvSsUrC8MNf+i9/lig16xHZbNWF3jK
ZDWNgC92S4g5fDlAYT2uqdMB14Dkx6mPHU54oWSu76SNoxAMpIXtBHmmnjdeu713
8uCa9LjWyYtv0EFwniLfUHgS88go/husMN8R06vmAWHt002vERfU0Dr1jmkHzzVD
KVu2ptnbdtCCYlTE+o8qSbEWSzXmxmNt7pQtVUY4EIeY8jGnadHEc7vQyG8X/Q/6
Ocam1xeMHk3e4WKe1/u8EBikehEqWMozYb1dAAOYdgia32Sts9keDaYY7ZAuh0n5
Vef29rolzWGWFyr1yL9Q97/s/FbG2w6D23FGcdrBxs/aIAtHIER2ZAcnwxHKpg9o
Q0n5M64koCUENNijxutbZlilBAPPYBDm3NHjHEIuqNyIJBJE27UobV/N+xfc6IaM
Y6wi3eXGwF2F09VFB9qoYocihp8BW0LC9pv0U2soSixgowS+k2UnUbTH7YxEONq7
+T7O6f3m5UMuozXU0cOn59SRmgZH7u9NCa7Ty/eQjLqpzgAKZAafzyQEXGfPmi/j
tUxkRuvicu9Ux/P+aYRb2k21teNr6GZPELMEfyEEB24Cmgflo03f/vv0Hi8ClQDu
IEj5SKl4BLL/wql723n3taQhHQujRqNtzHokNFdUi6CvUcaON2A4BrWEIe0jzfM1
w2+CWENLiSZdAzWcS7bYWWvU2DyS0QfRxVpq3U3bbF5yhVxgromriiOEt2B3Qs8H
bXII41j/O2boMrb2u3M+7UdixCrFK/nGoIifE797WxirJlUYIufqzaSrjr62PMuW
vg0+ul3/ld6QfsHRus6JZdPGBB+z4LeVHwvvJfik1TX+O4EoXVseli2Q05qzCCU6
LY2lQA0o0Q1zaR+JtkLwug==
`protect END_PROTECTED
