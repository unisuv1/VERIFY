`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GgdWu8kVLBoAjQlD654njrMXziLbbgS8cVZopBVQZj15nc7qsw1mYn97OzJfdBn2
QdEGDmeJewJSE679/MKFazG4TeNKqSAT0ybqKQGc3ll6r9KQgTKeFM5VvN7XlvY5
n2vF7Fx9C8PUxvvyj4xoKbYtlsBLJcKEk9RvWeQygPii+H5jWnSfPUB6IMsafZbX
Klik+L0S9D4v35lrUtvSDEV4AUk4kzgsm8vYTharkgKIFHCdnSpA6gSymbWK7J2g
tEBFfarpiTHNQrC8+wKYjC4jOLllX+rlRKjC74NfYsOfUJbS1XiHq7j+uVYs3tK7
gKm40EnERhBlOmWGLlUf/SDe6gFHct5ATLwtDcJkT7MUNHSJNsF3Y0JJr7+EnqOD
6KG/biFlIuZtv8cOtdy8h2mr8n3xUgJI/QnArA+EnTySIDfOfN3niv3VJXNLN91j
v3qLS5qU64FwX7iVg1Cg47OvWatzXHkTbQpviy6eorW7czdYB8AOJYXU8YoHtSW0
xjbEmNrXLSq95HIBSGn+ucxy3nraKfKIQHBuvvuhSHVEbTodPKyrAxD16A7/uoqh
gb5Ope2UcCk4gurMpgpG5yRWANgxloYqqGE9GjyaspmCucSttmsJVeYHX7gdlaUF
xBohaY798NqHadeFVHxrsl89LVJzioVIR0IU5aJBBgqSk9sd3vFBfG404NfbZojV
2B/z4gf71Pt+exqsxPfAdT9VssWlB5nhrZ5oSgWzYUOLTAFb2xg2uD7DZ1Iyrt0T
cjJTG6Fe38krEP5Yc+AgDFE0FmzGahjoZMKKQWUNaML2fX7vy3DR7+JwUlJ9w399
zzXI29Vys2ZWm+aK9/08vixl8dsGDzYMXx1yZKQTw+7FzzSvjAgkuTU/LDbjfjIa
m7LTLwDmb7sCBHk3wf6/yKHym6z2/hzC4AM555+V+apYo1eDlzeXRlrB5ase49mB
xZAaG0Vu8hc1VVJeG/EtX2aM3ugOxJNvPv5oxNKlEMWlvLaUCSOca2TeTq1zhfJd
LeetEMY52agvIjIBWE67dKCWoJOkJT7IzTPRpUZNM56UgDAT+8vZqM+M1T2Lp/GF
P3VtfBcG/7LBMex5DOnppFVX5Y/JqoAESeDTGUmrdgHUxjRGM48of/k6qOxp0G8o
zRpXYB382LtqgpzWyUIbXuL2ErXt3sZGq/d7bIKqfvkO+o2s43X/ct0RgOhAcuUL
dBGv1o+sSTHIaz15D2yU4hn1Za49TgPdXrG1qXN36hjX3OPwYy+BainJmTXpEZfW
SQpWC0hbvbO6CProNwjR2z5SgR0wmB2hEssDfEyiSQxK+5ay2+oZZT+bCPD4I20e
2paGNxTAcN0krszEo195vlnB916jlMCZ1KsreUmE4YA1RwjP3H8gIOGg9iJiV0Vb
FSA39t2O1OOqQpz+vZx6p/DshEu67tQGif5kfwF25vfx5AEKj3TYEspnHg1TwAmp
/2NNItQgrulmIGALC316FY8dfjTdNClXl3seI3EtL+7FiCgdwen5Qk7nS8SQVE6h
MlXkwdE7fJOvyGUe6BDeIXSHLzLJYst5gNcV7OO+FtrP0hC7SfKbsg1F5ZKDeJwW
s75R4iuwWPZ9dlAquq7JFayPk7iVBtGL7vpbBoKfwTefD1dQ2U59RFb7a63wir5K
WELYvJUtbBhFZwz0BKVET9o/enq+uAWT5Q7BRBv+J+F88kyZkSI912n6DNVVR37i
uhYf/okcKb2LQvqFqrJ8x5q7gJ5wilAcApsRz1bVJbTkG1sHg23AQzJP1uY65Y9a
rBsxUbhDLsRxPTr/O9Eu8pkv1G8QILonaViFNb4eyuGsCAAFP/cQ/XDxOql2Itc5
yLjGiQEhN+a0MpMzwRP3PSVp0TVC9zuPVyXipvMwk7LV/FshviMgMir/q6PzJW7I
pMoaivQAVwvlnn905xsiNk2wzxiMOI/TamrxPUHYXu5cmccAHoDS/rst9XRrnF+K
YHE9F0/4Qlz1nWb1HBl8em4lThHc1ZKGR2wX++fglxLOgKM2g5+WWlCulvL0ozjd
OUCEVg0vdRBu8i66RGGE3Mixen5mop27Rcp7s0SbQQkSwiFeWbszSG0Hp395MR2m
R8pdoTY2mhlQ3j1zV4zi7YMCU17Jes6do7gsq8WPcRNZifB/qQZtQuuhxox2a/8R
1Cfo7v4eW7f2uHf991/OMuNK4O0JP3EjOUpQazb/+ouhO8GbvDAooVRyGOrCQY6U
vrjbTNGVIa5iJ1j9ZT1Qw0AXIpCjH9yNBYNTRnaeGqbrw6XKlNeTHjTC1fqCA3W1
hfiZsSOt2qGanIxCWbexIw91LGelh8gYLTSEOTlfrVz7WX+MfYRPJsvFO3QJNbYY
MNEnlYMsU+6HajBLig+cSGVN1k/u+40ffPcMK4w5BkObfk+G++c6y3RiTmC2FHQA
WQzPTaPI2J5bwVFIyxucFjUCzV1bAPQ/L1pDzN80BneCjtQYONH2m5WGkTOaBNoU
6c0y1KyLqEPxBoD0O23Yo7pDPtSBfTGuQhe56uq3Q/2YsW9BmZzgLZBzH+nPnDsS
8/vYtIufweVzyYku1pTxFwk6rLqASa0E5lzFYERhToJihaWYqHyL0VpDC1jFsKyC
AukblhPBOAr0JupeebikeTRcGwlyFBmEgjsE14p1Ggprm0olAo1ONDn2Z1h0cWab
uwib9kwgUiHReaFPFh6qSDMoRLa1A0670PcuuboNfuoLRcI+XR4XpCaRzkTaOntj
akvBynnyNunwag2qim0sydIW46aJBMWRbAJkKkesIZHYEmkNXgEWCk+4203nkPgi
dPP0JO0pXiz9Ov5HvCjvxfrmEedySucEBW/tvhuKWAkVJZ5v8FQKJWzc4l3UubvX
OoMJbA2bU+xgYc6lC7kN9zhXAyiEyQxpoV4fJTCcEflzfhCqwUbqbRUmfAvTNugM
qPHAJFTC1nZv/TUS395uUC3aq1nY/PghiSOlM69LJShApjATEcH9+XVlNu3tJC5E
ReUwbRjsomFEGBaKXmZOhKzL2t4v9mh6JOJbGo6QN3YTsjp84kCCzfQfj25l2wFy
zxwsG13B4U59zLZT7xddaKnikmNHY94e/8iZlIKhnjPO5y2Go/05891apZSK+qtF
kDFocVWSunes1lCWFVB8CFkrZsGSjntsShLkHJVZr1avXSUZKwV9NsWs/BWoBK7O
LoNESP4myf1RNnhiKXyreqgnmNELJ1lDcXg87jPQAnrTQHFN/f0ucT5B6R//H921
2+eOSebv3Ab3FwFNN32rEv2mrgi4lHJpYSpZaTqDq4ZIsMOX2hyll2rb7B2SpjCu
bengje4jBjaakS1tZ3ISax9owWvuDI5dpEHJpWFER/oFRauWAwfdH2RxBAdtIQ2A
5ZpF1VfT1U9q2NUGWLX5DqHRReXU4BZNBmL+byW369STjjJukEJL4hjWCSSWD/Il
df8lQBb+woB5P0QSZkky/jrv9/c+uJo3xeJn55jrs3ufehFGSqySYoNSJsZMewEn
QUV+s+pTJfVAOHj+X2gXIAD+S87U9hdc7x+uWJmvazsFlTCRefKpojIvqgI7goGX
jQq4tVEAMihvRb3H5GhgT9ayhJG5ikNB/Q2l2l7QmwT7yZpQBevnN0K4zW6tqeZ4
mLjplD6WjIw5m2ZQ4xl5rX/ysd7BEzGnJ3CsjJvL+0bmK+x2ycspYgCZDO1XBHJd
sI2pffA10lTzoQZ01pTVI39i7lIBs7nkTgQ1eWyq25XlME+0zxh9MZqdUGioqS3W
z/zQ3Qum4quCCSbGt1qL/25nLq/F3+8GIQyv5M073hmDLEjgyZUCvs37ZRio1gzQ
erYdEwyvgkeDCWnbNsy4cpce65N4bTy9NW1vfr5TAVeUq1Jxo43fJqx57ztajXQu
UsYDNN1u5DnEKDyypnDblmVDM8zHZWFOxeZZzP+OyOSKJf8cjKfKue9PgoV8wWAC
XyluRgkio/GSkzHZ7re93lHepI0Up14I7GZKf4a0AKwlHkLcYq2MHFrUOcJl0MCK
60rlVzHPSIn71Tt+42VM61lRj0wZea6Sdzh9kovI7WYyxQOmnjlDZO20T0dSAKTB
i8iHRnDgvxA5qiH3orvbmGN7Brv9pb9Mm7bkWklk3nvA6f4uPT7YOh0POLnJF8rO
ChRDBBkG+crn5bwbsxgkLf+33+Cd3rIMQ00s50ZykWiOmm5nxycTk0HhxNVZ9jnY
5PI3DHPmhJzkKX3OHf36egUTKwCKuoKvHopkjNhqgzDXcY3cuqloHBXInkRsS3Cl
mp7Mk5mCGEy3OlH+C0MqQl7NVk0ckBfY92XVnoPYK7vV8R3+wKfqrlgqAsXOIWvw
97ugliY736rQLJyfYIzz8vOFBuYAyFj6zZOwyo4J1gX0lXpUBfNVU9eDft5ALT+e
jGjPt/hwm54WHzcNPXO4JYbZ/k69O0QS0b43N+Towo2fQEfXV3j75vPIR3lqUJ9m
FcBBQFGRHvk6aSIQ36JV/4KSryJw3zzDogXJ1YJSCCRhmiUvms2CMpwFAoEUBhpG
j8nh6eq6nXsD4dtpOuKLlqVRWOIWcnQGBKPq3MliPJhWDnFCphbyRP0JmMkAcZQ5
Re1d4T5EfaCenBC11BPUTi2TZCGa4x3ZlvsxwrZf2ogXqF/COCLroyB35Q26mxkP
FGxgrfn7rGr83VsMJh+/72dZXKyVRe4qppNuSeimC6kyxvbiao/7vYH9LtSZC9yn
tgRYyh9rm3Cq8qF/v7j+kV4yjfHvKlLKXXKRuNmw8jQuhErV7FRulokPjRgK4qob
EqKWTh/QnnpW4dgPPy5X1KrGvctzkt26dIEA+FwSJFm5FacGvsTSd7X43SwfE7UC
9+dYZqnEDtpe2+kc5hLEwB392/+oIJjRX308Ixa8MVlrC1XWJ1u5bXeGA/EE17DG
rvqktA9Dlxh8+OyqqzBEiR3MdIEfBTgwQyK13Tw2VJ3zn0F30DBOu9DfUM9KO1g1
fRD9PDhRD56jsg6rO1jKIZreu0YHnpfYKL3vfXvR3ZQaq5/JF0wFZ1l7JKUs/T2h
3TT8CbRnLZAi5Vt2dNUCS2dZ08n0S9HIMDlEFmidu5LfVxeb/1ATwzhL7gcV+B/B
e5rVE521S4+ATfrdgIwvGeqUiiyBNgpyfRC03CeS3mhcn3gwRDddgOkZEKbFTOjV
0HPDSPIJ3rbWaCECT/LSzQn+RvWdjYzSZmN9+Y25I4pmrkB12NJTHD16msPLuQJw
RVDYb+W60EHS+su0VaVo9t4yCaD7AJgMVyeAieD3KXKjGpuLAAZNHAfOees4vch/
OnHF1MjuKCCyK27lsLPZPnMQYw5VQ89VLyLz7eh34DsMu4KQPExOuR5y1zN7oIWu
S8GMWWVOCE/hpKBrPKxW0coCFtfHhuuGDhZyA4T5oFi87cMYFrXSnNd6xzLswNxJ
uW8e1VzXtb5fWcEIfNuz+AhWDH1A/KhvDKc4sOsWycNY6RpjFqYTFBHzldknobw9
dd6L8k6QLT+X8IgLoLT3n0gm09qf3gI306+nt1VFWiwRAa6O/bBnu+RypZAlxz6I
uGjWyXvby5R0sbXFsiUoKdh3wQjmM+yuxhi2y4vzjZJXi9sR1a0akcY2G6/4/M3i
APkTHIYk6UFx+ftWcqytsQihjnlcYidWudvokc0BFByvl/fNObtSAb+4mDp6p6Rr
U0mQDiLRJEZ8HoHFat9PrLEXwIQN420EVOwoEvf+AHQvucgLR5NGgLZN5hn2SDhk
u2BCUjf3b9uQvbEFH3eCwUe8GgEdO40kyk7FPUfjOzy4p7AfRTxoS9en/nZEswRO
IKYmAeWFtu76En9lrAzTkSj16MYSCmSo6duCyCYdK9JEMPRG1BMw7omUiPIG4vto
pXxBSEFGCtFKuJfkqrLIbG659JBE2V5UGrkl14QbXJ/htrn+CbFRbexAb/+/mZFB
2ytNvM2Nl2RRpi0qAvqDVc57HUQruP6fUMMJ+GUyGrjpC4zvbQ4txiUrNgKX3hI+
Q2UwpWNf6SD4np8oP78nftKMA4wvovaXWwriBnsA6X3ByKTVg14J0fmzPAWvBWot
+rgEn2HoKIz0aM2LfqZJ5FrLzYSPb9dmUjc/1dHBATsAOkm5QBpMvrTeygw/0Owp
IrEL7kzRjKPKYIS9CwbfZnqtOo+3z9ECdybjzRiDE9erNfFp38k6PnRaqwEfIepC
gCl1xeBfNDpQuoQhWtDTvMQ6FAnHSN+Ei28JKnF2pWEvc0+ntz+Npox45aPNjPPF
z2FgCFqHnywHJpZxzrtMK+PCEkzYXuTN/dN82+xLgWPtgE3qwHJ/oL8bwrZVMQ/r
/P8zVFXXeXHsZwd0eC4BgU/kzrQYm6Bw5es5yU8fyss7u7Vb7ma7N/kjF8tzfWiR
TthYKCtmCbPofKAw9uj89IL9CALX1CJQrPT0H6e8XY2IZQ9B9RvjgXm6yhLNaLrP
3r3Uj2iiketmUbEsUMPR0bQSxL3nawLEK6ifZXySYvhYvm3Hy2d/wmznwky8zV3t
OxcGoHY7YDe9Z7NwDL/KqPFb6KOj5A/vzjly3VDvGaNDsdesRkoQ632qVq4hfWe7
JfomKHhJxGfBTi1iCmANc8bKHfUN0gulHtM80EdZH+B2VmAQ8Qw2EimRQZQDPYZM
f3vOWdF3YwT1TE2uhZmqTw5lQOlvvRtFMtgTehCD+alAztt9HrnutrK2pF75ddtj
ZCZIdp70h8CxUH6DvXkyiVyr4q4az0Au2q2MZNSkeQkyPv4b820Wbn+YTamRtEDZ
BOiw9i7sevdk2BuGTCGqwkbmjdDaoOwiPqnWhsgkT0Km1dCok+1rUG8J6Ty6eTiN
nV+R4lh+sE0l3rcFdgxZ7eghfo1j8c3e4wWh0/cxxg8zvji+vvasfJAVjjyCsxpw
Q0P/6NbSA+ztpcNss139B9vERhXsOc/Tger9gTu2wuQhuHyl0pYk8EVtQI3RF7vG
N2KelCAqly/ZbSIXdiG07R537Br3FoojrOLE57906ya0teoFs0TFqOrQA+sDn1I0
VIYo/SME/5+f4GhfNxrbIoGr7qggI0w9AtIOa80UapMrPqvEmwXP998GE2UIqTuz
wXp6fIvkGtUnDXFNG0jH+vI4i1ALvYKeQhK5sh+lgJOaPA7AKcboFyQw1ZK4u7R3
CsUQdJFIWxdyYIRizaloTi9zs8sOuX8zE898Um8HlWZA+4sOx4b8b9OMgbxftOAX
oDIUunk429PMGlcYpjWJWEhuFZofuhSSvKK2tvWrM2tfrSU7m+RyWR13pV1xJzZV
pDiOrdKFgIoTuPyqQzcYjH4C6zcZfdL7WmkNLW27YbBCfXnEv+snFzHBIIHSQvMO
0nn5k8gbZbU4vU0e/KBXKqYbFYHRXz0qAYXwjFDDpi2TcrqEkUhzCOgisg/UpKT6
kfLquaJQ5qR3R7JKngZkR84BArqUaNXuXb+T2GZ6Um6FlwlHTypaWe0pM0ELtRAd
QP8RdzgWNIZUU2z+GpYkX+W196A3miyIhNCsKc7VxQJoEgY85j6wieKZIJzu7w44
/nDrCYODXK/XLUQsjKYNd/AnNEwsGqK8kKRiMISbMoo8porZ0Euo1C1hYzkSjetZ
4jQYxLZ+5wJetuDQ1PumtfdqDOmrgJg3HW61pP+Y8bQZeJnU71WCQ8+aYjFA2+m1
9mKJ2t4ezxu6qqm/fwsHOCHuDbb5R4iOProq7VjgPnPIHnVcDhPZ9grKbBMt5Yzv
7jhW7yAuNQINh4my0vtXv1OpXINUfbBw8ptQwGntFMsHaDIiAju3WYaDQGkOF7Wg
Hfkg9LNEPHrKb8pygSkO8+Q9V0oGGNUipfiMjRIXOQSG+BiK3WymYuh+ki4NnWwp
C0Xr7ozDtVDpIa8dXOuCHr6RYY2xvdrPZHy+Z3Tq/cRYhNb0Ojcl82mwMHuePOhV
YrQ0CJdh1fVKmeygdZqYlJNU0SMC6zfw10/Yqrj88jdEQ6NhxqCHzZ/m8hlrZ37U
djTx9bNT8sdvgnfnQoQB05LQLQuXAuBvvkicnvcmmP8xBNVlNdm0YfHmdE/eErWp
sUvH3qIAnolMfm6CZKILjfYejnzwf3Odr0W3kHs0kzoU8E92XBwOgdjY8yBFLrrN
8pDN3wloulYCWb7gu6j1m6fuuFDtLRvzaN1aOigGqoYRrNZQ9Lbq0Xmjzjk34SVP
+QrDg+rhgmTSCG5BaKCDZRXXXdARsJOiJ5XmvEKfWV0T3CQwNtyj6UUy2271dDSZ
TrjGBzCFhnIa5ghT0mkO8yE3IfeenadFmlSR/S/JIcj+2FfnVbETUPLXm/fDFpMb
dihnBk12zBhpT61WiWgwdsOTnkG/qwaUBIq5XiyuCf1E4u6k/2pWtVxYhgSRL+5Q
uoFAz1j7K8y62KsYGO+9uN/BsHQ73BmLnbJmEOUQCtzKWMeaVst6J8Co3x9cNxew
dp1gVU7f1nmp9hz/6Nnq/P8guHJZQ5wh9bMov0Bm2yaTqdgBJJqO2R0bVQrkAdfi
XYhWkH1CyFJQZCbJh4q4RxTbD6DMCpLiEWbqC+ckIEkEXY3ukBbu1hvwGhh3W6+1
sEP10ntoP/Jh8hbjuqJ0SMf8Aw3JO5JlnWxgPI2kninMO0lvMMFv/pfck4C7AOXy
A1MN5jHtAzcNK8IsLARu/irgkQzjIw+DeGqoCnyjtxmed1Svp8LKg/G3q2sQx0jG
LKMhSFqpTfJ+0TaYpKukB5imzfye4wGvdk9tBOMn6gnM/RegRI0sfLdX79Xg0MS6
zAO3hDLORBGTCITgiUBNQyWd9R6h5EuQrUYBSZOisPDpGifbqw9BQkLfetcXZnpd
2Y4CAblgCYdIyxrmd5i0PnSBVA59lrXgsUFMV2ZcFLkhlQHOUl5Nkzd9503o7s9t
3HM1Sf0hz90jxxFzYXhj+WlISl1+P7R+cqk3j+QUv8Lv/vS9KQ0KNzpfKnwm+HR1
Pg9opLyO9PA4FtYSJ2WXAGvYl11sGlQ72At1IzHPY3oiENYwQNVG6nZyzkGIaKqg
UO+tdeI2GkxiqWyRubUTJ3OlY+VKGlKp17u2jhpmy7bzzp6wvlwgwZFHwM6PsU5O
IX+0cCOmr7DHXxY3jIHIVpQqSimQ5pJ/48ptORBK6eB4RerAKXiX52M46IKIXarV
dMDBE1bVPhTMneQl4ckQkDwKuP/Syo/84cVh6/vlnARP9ABd9L21kAKZUYGdWL+7
NhWgXfHgD/8Bp6tgIUV+LxatyqmJj6/upiZvtdaLQrWrV0YILdZHp+M0vvIdrxHI
jOVSpIUA+QfvDfdrBvvdL98MpItptbQFMq7Sta4TwlWr60SbBDZcJ2A+JyZX1kEu
9jqQxjB8NPLBE3GRsg9DjmZ7uGXBsijqEVwmtfUVAN8kpMFBFyqQozBernWs8eG3
hLactP4rJErzvmstT248co6OkymwbViTY+AgB/1KV6btN8ZHQXv9oz96VHJfejWv
CNFnSDflUmRlyxTEZ5snUoBSPNoT+XwFv8jVce2j5MYOhAx15kJgifIzjRfiw/oO
3vHUKJtWfKW/8udq5E75Q6mcQxro2gbX2qtp8AXPV+Zeujejd/zeyLRpXOG6dCiP
MUd4PsFYsYKBTGnIYi/mx2LCOYPc8CUaEazt9wH6X5k8crhDZdJXOz/IHidsf+sn
AeZ989DxtsD8zNYiPFXx3i6NxMeHYdnMoVAO7GJYV6TEmV7qu/LRjo7KA5ZM73uC
tf25vUP4A7r/18MLDuPbDaVgdp1YUL7J/C6iR2svSY7FR7t7Z/qTh99xpY26CECR
hBeMs4AbVrEFyS2MVbV1EvtxiAILEu/2T5gsGttGSAz0gqxSwdKH42wPOo32hFrN
fvH/GqHgf2OtW0L0zjGbCUGLWv/bmXQmjm/aWGon+Au2gGV6jdfN0iuhLWwFv9F0
yFoMLfUi6GQs6AA612vis9lXV7XLqGRqmO0nWJ8y7P4MjMzbGh5s61v2t2D5LOW7
kwbqTk0R/+HKpkzzZdFtnCsb48PkxwELTVleXlosY8Jjqb6mlRjMqkwvZd2OtDjQ
8gVSGTD9GdL4dYvvCeX7bKSO89PpMw3Le8P3jHe9IWiqyNphZ9R83NqRB9ZowxsM
iTU5Kqmyd/fV5kJaomx2o+9mimMb7DjC2EQIFfsDYm7ANpRaORdw0RyH8YeX7tVf
K4OXaLD5CixK5s7MEdMioIi924A0lIknpjr7clPlmG23zRYKJCPG1ke+5oT88igN
xopmJaY81B8gXNXz8xSv0oaqogmQN1WcHDuag1ON09+euoI43UEncRG+C9J9EWBd
wsVoxlGE1m92eIYaCIKd4GcomIeNEhNWdEXT4E4xAzCb6XCPYXkwaPP43jLZiiIo
Cuk/WVSLHpYbq3aVIUCOIzwpRL8eciJAOaWY5XQQ8NhjwWVogzTL/KsIi0et8RQT
nZXpKod1i9fvroh/CLhOQdrCMGjdxIuCa6wt8B5itOLeVBFhV32KsSbEuYjYu0sf
Z2SvcnWa4YE13dSP6+mXYNRX6FloZL0YfcPXVDCb+5wMFZntOP1uBqgCUFqK/Fjj
3CfjnT8fge5CWf6i/GfyuoGDY1VSqJ18Wu2KrB1Xl9Egjl1xD2FOq8OtsjbD1qog
9Tti77nvkXAFNcqyLzyQEi1qvrNCC5lXBlnzXUbNSuweIn9wi8LsE8KthEel03+z
zFVxKXZx4Khh1C9pUqbTkwGEZy4jxWDOfbbZiuq9LQfX6tIkMdjvZGmShzX3eftj
RndJmebB61DtU5l2VTfr7CZQsQakx2BGBd13uDiuuxthitcjXGFLAsa8ZD8IWEZV
CDkq/lu8gBLLKdmSPjaIqeSGzHLKN+b/6r14G+LskS8aCZzfvRAAqfIszkxepJUG
B/AXh+OsSYWJ/5GYDxUf4KGyOizkOCkqdbwDtf6Sr694f6IXFrzfY9PNWhtos+l5
yZdcWtNvQ4K7d+gdDltqQLr3aMxXtlW7/7B6wxtOSLx39gnn0kqgtvudkp/oY58s
P13FphEPCMUE0srKvLqbzJF2tfK8vRdFuVe6yNf7cJrkOdHX4CFopcOsQkHNrcoL
+tFVYP5CDHYpuEl7vjVPrFcaDPMzmMkBvYCg3BOggswaQPXMurFuH9HLFgxNIhdt
cmIDgvuSPBx7GpFKBzEh8M0xhp3qe6A7Vf2cQev4hmFV1Db9IvhGmOxxbE2w7bXv
WbqOlMZlcoLzThlPsrCjh3qxVPE2zhTj2IvPtfw8fuFFOo4mA4k5RnGcb+UM8KrB
sC70s0+VEm9V4dOlkOm0nZkQBMZrSWR6cYf7bRs0kzLUFkObdye7SS8FYIb/EogO
j6Fi4XKijMq1+Kh9bxhV/vwx/vMDliLIg+nXpQSwMDU5Yeiq9WQ3ZPUth2A85ZST
Lv+sgVoCqew0Ad9KFYYiE5ut4Fu1NwULjqCqIyiCdOnO/deKpqjaKWxZaQaWnhes
S7qBBH4MKpJhGyqOrfyzx2SQr6R2mFk1FapK2z7esnk82SOQ1W6P2q2kpW7DFfU2
QdVwf6D+YbJcSX/jyFq2YKlJxylUZliScELnreW7lslMNmxRkwreuOVidbffDuLA
ow5yzbfEdfCVMCA1Bc52LTjEukfYvR1juFAndKpuxv3/+Loe0Mox09Pl8BpnHeWJ
ILSLTkrQj85PtirEMAZxmXKlLfBkZ02/nTYUu3vICz92+eQFJwJS1l+Y0eiC74i+
lV+01nvL0yNooYJebNBJhRPzw49RTnqRQ2c7k0MtYOId+KTKz7ssVQM+yYFuebOH
I6MKVA+Bq2as4Me/3TKGL+scxtQKoVZ8L6jAfXsoMFfhulFPCjO+LJy48hOojPYE
lHGFp/uiD6bTQAYluXPhezFRnPSnSPmKo0YWWK516EYDmOxW/afE9AO8feGW8LpI
zbGPOf+pDnLom6M7dXpNnojQw3qwaACfv+OF0pvk1XJBk0kdULx3H6B6I8S5BtXS
Gcj/glHOk8nxhSXk2jkJqoEmMCSzDtL94KdM4okVh04MXrejf0JOSNCe6hF2gje5
/Q+AJ9dsR756weiCRMAFE4pmK1lazUKj0t00sqU229SzwJFaoyJ51XnAQPYLKuMW
PKBuRSOkL+1qsou0tNCtNF4GDrAsABJZR9beoV9qUHg2a6L+Cp207fM0Y8uIpvly
P2k613W5IIvlykrWW8C+xOmkTpkrSIcIvPqr9DQe23z07uJcvI65k2GLHuq9+4km
HytsDBjFk24HzCoF43QYUqNbCccctxHrY/VvpivVTxmR3lHerJqG9k+Oqcjj5cGX
WlH0DSlSGCwpbt6qENsOVNg4lO3sW0i96QFghQ3ls9mgz5acyLq+7Qb7zzmPmK9O
m5xtMA0e9lUsRjNs1bEYyy8Y/BhJYZo72QyRu3wr0zH1xB1z/zsrxJsIXLlhGoL4
jliLWiRAcbL7egmVXdl6uePuXqufk6xwN27aYqWo6vl8YOMA7kkUBf3xojUvRJDV
V/7QCruUIXnB+RUTGk/fF3MTG/KyUdXQwW7Dnes1pm72JcHd58yvisKnvYT658hz
5gzD4g4Il+Nm+MFPWOk5YXmXkVIjnpcHW1JUcsTVPqygolBKgvQxzfQvM0aIMy5A
0T9jBLm2NMqy99JJKdMtka51Q0DkOhO/86XwySx8nQyVNwZx37nZewa2pADexPAk
8uVgAKz1pU3OTjY/BaP61gARaHUTbJPS9IqE6KcGLAXDpZHDd+Ll0vALFaDnEbsm
qG/c1XkId5KPcRS7xyLYfKyuhYosvrEWaMTb+yp5sMVSRyaHoe1N5i/iZ4gjeh1E
ZWYu6fR2sGoXfK4RI1FahXBEEL095xL3PRhz8FJFzFCLgkCRDVmQ9kUt5d1LFO1Y
E2rXmCfkTyNl0lAXFM0KIPi29FK322Nknc1RcUfEm+vRkmQn2mol2hOMph+lgNZE
Oue9kKP/pNQwzi9vALjmMm4Kyo4aBRhM+RdxehFjnQH/LlPuTnLQLYZrlG7mf9m3
DNGBHdA3OTeaAjO8RD2Vi9+aut+5RgLmKe2xCZAvfM2XNLGA8VF3CvyJjNRlCbJO
gvgxdtF3yWLbL0dZQAD0yNyQ99RjT1KtO0ZtR9w4JN94rdI/ZY/bL/nOD9D3PTPO
+BXDVt/S04tpWhQVv3Xiaau3n5jAWAivwT7lqYrFIOYB7Ln9soDVyfadQlsGGdAy
dUBURvRrGcmiN2IU/YPflHoxUjwUZuqzzJjKzOY9w8Bev+mwCjdUdKHBkT85ws0p
nxoE/WpIzPcJCECwndNjzVsQgGIXhmJaIYyxN5jYHGc1K8gVvbg3gprr44p+sS75
hSMS9wkEhMWqAOeWDicneen2KHEo3tiTTJbRUrDztBOFK1Jw1h1tRyaoK+7HAp5Z
8/CyB+TMybYSRFQvkpkqyAxhdWIZSiNnfg2Adwh4Y+BHnDmUEb1GFNyC1GB6rhUC
l0s3u1TDWY5xjhOzt5H20aVLyIdlUw1cBgbfJjhbxGFJqVnd8VBIfjrOaZ52DTo1
vMxCJkINe7H5LC5xSm7xDBlRc4+L7wkUcJEB/OYy6hlCO6UoCoKCwe8VrbaX90qZ
gKB87vQjXYe+AdIJCwjjC93u3vIPm9ncpKtouXAYXjVwvSZ632VTyibHWepWjqSk
wb6lIADaY78kcfRn8jfhMO11SvbF+tTAOtRKX3uPu0ywr9Z/tO5Kt8h/DXhj7BlW
fWVLcLWRS5r4jYZh6ht1E1uI7yTgRM5K7aZQuoAig0QXkges0eEexBQqo8s1I6yX
D6dQGCsBO8P7H1CvW4YqXXdUjl9SmPTtpkPQNYe4mwLtW73Ho9C5INipRQNavdfr
KnILhrJX6/cT70u6AJCLNANxkGbmfgMl+i1uD68XJvmXxwcggtnhxf68xwd7O4Jl
eo/vN/eMqWtnJViGBBjaz9yxK4NXkUpNj5rd/+xiDSOdIs2AEam0FzrHej/mtRJF
Z3H1R4IQG8JYqtmN6/hCBr31kQMVFEGnS/qa6gmcr+eqnmY6yJkDX0cMzCJDtJ4d
tlck+cI3BFsTqC9nS46IFXGkWwkmPvuYhqUwjOn6FFlc74dLi6b+FMwTnq4TI0LX
6WRIz3nvumqzDgnqmdGNYvR9PAKV3g+wyMeNpwaa7qPyoIXAF9Ofb5JsOm4n46iZ
yPr4725uQu3fI4SX+G5KxaZFbk1EbM/sPjDcC5Hn4ohTRW56gxMiYP8+Hj7TSYrT
dkYKA/LF9T1fuio/GkuI19Dt+k48HXM7svyBaSKpx6JcrZWVKepvo6yLORU/oX1t
HRGAgl87q3b8DQvZJ77HJprMwff5kaI6b2Y6Ph2ieI797iLr/mYECiK8caNmqylq
tW8DtfuLpZmifqRS7Z4S8BRCEsTrT+/FtsETXO0bOgcoKvOapRdqccautNEyQGwA
5ED+IthR2B/X0UzSquQouDWSnS3Fz1LCD6RhUF+tlhxlo1b/vn5tn8pU57Y3vQNt
sp/w/e+S6yWEgXRnGag9GwpvDckWOqvj4RsfJ1HIz1XzvlTu36DMOQZe8eL+SVMM
3+UDQZGBe6R6uR1FwX7GnxXlrB9u27c/iPXoIyGrEQijdwXnaqmNhWMUcE6h9TOD
9c9sS2hG/idM6cicf9WjS+5ag02pTK6oCOyD9oN4TzZDbJ1MGm7j21wLq0nCsk/T
XhWKvgCDLQsKq2TIecknjbgcsuhUDA9B4m6SsM1anS4wJYqXjcSipc8k95St9szK
Is0xMwZ1o+ESfVEyrMw4Z6vYCi3c7Prum5TkPZOyfNaRkEUUD4KWoWRBo0V1rBwS
LpR8MEh5iUbs8HCVRA311DB/b/ClPxkBt6AofdT8GzBE0djJFZKgfHVbhbgedk00
Jna6fnERStPYxa4wDjkDBJEq/hhHK9MxbTiSp0svAjM4/vanbdL4wQSxSbsd8COp
L4XHOaqrVE8SCvrdbEH2wo18M/Symof2hgsC2qd62PRRNuEHwlYZl64M/p2t25zL
/x0om007h2gAJy2YVxVf3s8e8JR17qr6WdHnZEeZx9cbpb/JM3bOsVAn4DTL4TS/
h+bmCoD59qXqwhcgZV20ObLKw7NSfIGIdnsp65ZjxQ6+VmOR0vIHwFdVkxD5c/nn
Xisdeo8s1L4Cm2GRiI7NTPH6elLdgO9wyJh+hdVa8IUR95smfe7S9xBAB1IlzFRn
a7aYOmivOPs4GdzzV1wmuQp+FNz3OPy/j4D6APYHCOJlasHnWo0xxXf2w7n1lmD7
/TsIQqnBH1h77/yp884jcJ0Hw6T+lPD6v5TT1GTqE73fA03kqYCbInnt2IR9GKoK
z1mQcdFGrLe36/mzpowh4t29VHzloQ5pIFLHMh6hfyski0zlJHN1CuryVSSVgLUl
deLCMQ8lFBcNKr6TEu0v2o9oOmGTEeZWHj3xgSf7AW0LD79wA8Tw3JV32OsLg/4H
WkiiK73oOxF4yO2tX+0a/4mkqd6QKgC2Eq5m2wPHtAlVFwHFP9ax5cQjUCRfXRct
KjSKiSjv6gCGHYoRB6ZsBvH3p0+X72VoLbyVeDviEa+qCxQldPnO/L312X0dO9MK
LrnlXHrID5yiiHyPb4KhRu1xeOfTjF1TNAxrdui/1uKMJqe2D2cQLPr3g4v13S7l
tAFX8347zbFN5Bsoj21oL2xh16B2akEHEzz/G9AdPK65PVV4D4Dm9xG6xHfqdfPX
tx0wQCxcctSLwBmUVIao1cmh/TUHAWvbPKC73AgPiTPsNy94bZcicinizyP8leTG
45x0CIdFTsbMUW+fJBB9RuzTl1exW5jR7Q965ZnyzbdETL3IY3m2cdZB8FMTtaVk
XgxJzEkgk4ZbHQV4i9VpUUl206StsI/OYEB9syxoWyEBbZiGfQXR0IybaYRiveKQ
v2bx2ow7Hvjt4k+Kp/aLCQdlHVSovaME3ejkLCpxCXlQc2JDzroRosN1nV2PYRbi
VnMyBm8FemaJ8+iy4ux9/84ue9SMp/MNpyEjdunxNt4moMQmSrKldRPQyxdaxug/
uY9K7MRrk+P6ZSd7spOSODqSDzn3IR/dzFRD8RXY5uGwIuD+iVGyJfWUt8Kv8GvY
t/WUHZXbAbtvjUn8aPX/x3jDE/uDnQ3jGSnKqQoxrw9zSUcuC3ONNyUxT5gDeF2N
o3CJP8Pvwx9ThOlFFCJFq6Cj19+bxt+2hLjD1uE4sXEVsfcW2+Co6oKzl04VE3qi
4iFdFj4jfLR4c9ZWysGRUU+UZDGXnxLcX9YE+ZuBxJJkC8yjQ7UwZL08IPMBGhQX
oSGPOEtbXe16PnG5++fXwYSZOUt7fLyC5frRG0v3Y2tlUTyRmumfzDMirFObdtxt
dxEN8jcfYsY5bai0AxmQl1b3izrJnXL8Reys78202fJtIuz6jwTkaUV6E3I9Vw7z
2dLZDsKTuF9mphjbOtqILcCwzZCTVu+1XlRMRF051AV1Sk6emRFgG/qpQ1h28+Fb
TMcBy+16V8T/ok5tlVuthzqON9HpGTRlcAPv9OaF66HrlL+9Nwe45wNoH0+CaTo4
zc82Pde1eRI0lXYh3vdVv3Q0aJ7AKoMzh+sRCMp5eHSbSm88lG3RI5EAgS2NLbbw
QyPftqYGUrmAnsV6FPFli13Api+dbIriroJrlVtPVmgk6apZ0jD8m+OtSmDdvSqB
t0xkNqa3U6TT/225Q3gOCHeYuuoiooLDjSvQvd5FuOHPXFOC1E7X0407O71tJiHL
7W1n+SnBCmWfgpZKdH0i2LctrTQevYCejJc8hnsJKgrsnBLJNT6sEjlClNLca8yo
lMoK8/L3gka1OxZFO2Q4MErTMB18DCE806wlOiW5Xf7BUUHN5oOHq8hBg7OIstIY
ThdTnhiLIVTEA4ju0uoKcO/FMmTV/UrZ4sGpEMOuS3ppHuEKGNGvjQb2nHyHPIHN
wa6WTYlzDGzMpbxbBCYriRYFQX4lasXOTO86bKOxJLTaqUJliLZ3wGk10wFdoqzY
mX4jznFFH80tBGXpbfYdk0FM/FbD1sLOBhnuvGC9qtam8NXIUQGHARtyoD69ft5q
m7qQ0fQ1DGFAx/LWhp2ixi1C98zH2ftQ53bRfGFnDJEo1fGj6HF4RezQw2/dkMQE
VAZk71b8tGigFm4W2g0iDTl1hexjnPtxChqBk/bbVEa57szYLJazo66HIF/zLowR
GlejezSjhkePN/cMf3rdDngecyGTOL8A0fo/CQrSWFCGSNFQf5vF9lXnztJBPo0N
Ysjv1uhCML2ziRyMzKcyld8CvERTnSQDKXVU+HoJL9VFPkZgFm1eoTaIryZ0pTA2
cx4Tx6SJWdcYOqJp1Bt1kGKKHtV2ITtE/EcXnQ5KSW98I84jn5omX3zFMFrLL6YB
nbqMqAe5VYICxR8Zy14bzvh/AE50NQ8WoqbIgQYRzGzOW3+QjZz6k0G2NpGu6oD0
hJH/Nlk4VPSv8NAGStQrfjP6FnnAc37Oej4ECAC+7y7F34YVHRZ3NiiKUFwgKsKX
KGRkoV9S3xee5fsoK+qtBhMtrGd5zDMkOwSCdBh4/vW18KZ9/mVhd061qMWzBbKw
BcUds5MJCCSqoE3pkb9FBPtx5bi31s32e+0qJSN/ETb65JHN92GmGCZQYjgtw3YT
93XTaj5oVnY52tO0fzIzXQ+lWIUMLvzThuX7vxBYQVxY0p7SNB2Xeh8OL5pMG6yC
Lgu4KeKTOlpOdUb2wedSyhY1d/v+6bv/oyyAP94KDESWUcaujQIEFUDKMkOmsVDu
Uu2M1Z0aIq71yZuPUs4Yua8jP/ky7Dn3gWhukMi+G1JsuwfVQoKtn6Cd4+fCL4iI
VhGkr+a4IZ/L3lEu8qYxRXnpcAflufBVde2e+arPSAZ45If8o1BKQMSj7/mhmZzB
Uq/PI0V028Ad+wZBMp3XZE2utMOUPdeGqHtuLvH7iHXQjB4+0Uk8mPXFNoIpKtqs
9ejnVNAO/5sfD4QIOmAt3bSzFsNseutbWCLJa/UpfFazW4lcXJpSJRlAKXqvXZtf
zKJixwq9SOdNwzjGyScQgPQkCNvQbYx4l7nIkLqpCqDNfGEybuXmUqzH3uvVnyqA
xh2IDr+ml0duPAkIPymfw4dwd048cPrgrRbgKL+i0UwsI8CaJlDK1zfhiELRoaiy
r8An0maXiTbNa7CTeAug3nYWvghtysG+eLDUTJGeDHqWnCEJj06vsbJMnLhlQhUc
q3cDvhFUyExPK8QEoUSbDiJyIxZcOB7GVMxWkOYTxahVx77kyZlbWWDg+50UZWnH
lOxxrRblNs2Dzf50QNUYKcPaPKI9xwhgSpGyW1E1ionzkxhteYSLER8ji7zcMRCz
INpNjWGJXBi9LmVYBG1e3GtY66Zt+nMTDFx49v+tZcsD1ah8BwnGBMYO4YPZy8eB
tSZ0GoVYPCh4Bj+aXxE1LOquiU2FE1Wxvbdg9zm/dH2spIXZQvD820eMm9j26JoE
GRNDFpYSofcUXYLOMeKpHCQw5Qnc136yOnHp5CYSpvr63h7L0Ze5TEXPHNYaLvnQ
ay/9m756RusLYIg6/uheAClIGwtHJ1fJ3eB5wX6+suOi8CG6rMOkenfvC64OjXAA
Q+Q380aRCyzdJztaHE+Ow1M4sjv55Omj0UVtWyxQ0rqJbqsWfM0qRsJqZiUt3qmo
AE99BRmrXRqOLK2NI5BRr+hCqRLEvSAgEZc1zVWYJubbh156lXsKYBSLNL/XR5Po
OqFFLzAPe7U9nDfWFaR6KNXUhsVUwAl053dp2C6kKJFXjQTM1VyfE6kafzHuLFX/
ziXBuAnXHqF2jqidJPdWDFRwbmWrnc35B+AINUwapBSMwD40SKAvk20k4cGsVYqQ
BHsJRIB6KR7wD+dIhomRiuUdEvqDn53N8aEzkgH2k/MBHDrS04SBvZvC1/DoT1j9
PbVR3H1ziUg33WJF1+tI8vzMPOePnZnIROjZDhorc2q0z1B5uO0tMv2yHp6wad2g
QfnaVKKp9wO0oyQ7Idg3ClEe2Ahst5mpJeFP53DTv64CHopNgnQJWL6BTkEK6yLN
VqURgBTGUdylsaOuX15EhS/Ix10ckyWkaPMppRNH9Vom6zdIN049vFs1FP8GCb5x
Sa/L36LcOWrdGlazwMTWeQz2u2WHkvjpyri+aBNQnDI3faXX/JNCf5bX2Vkjhv8m
Dgu+wlxoRqpB2vgNJuPeEspJ1Qu+QDptI18Ro7PdufKUmS8/YHK/N0Yl4+atXJ1t
TrdRrov0NO/UtobfC1ykyoiw4C8oUZtKJqqNkcPAWUJD8Yz4GSlVJ5+e6q41GXUL
nMRv/tZP6rM0TeQcisDJ3R0X1MUmLcq0LzcGI0EwCGTN8VwXZsruQKhqmylahriV
FWU4td1PgyFhAlt6b2vJyte9TKPdYZWUIfG/FJC3EjIvWe+yzBqm6lhlg5XZpbI/
QDZnk2M9ErNN5EmLk9xWvZst5n+pk6XDE/iCKLLkk6k5gqrU2JtHOe/13oms4M/P
B7JOB4ntp3+w1Owrtn/CCMcf4eFxDvevN6ck+L1eCBRQ0ZzHCOK0lkEu6YE6ozII
6BgSWBfnS/Rel8WVpKLkUYCnz0hkV8Xxq8Hl4AbyMcAVN/xVy3YPyNQ1YFC73nct
ALASg7+iEJB8dswpd1qnIxl8fIFElNJRq9QVLwGzZIquwsKtuG6LoYhq3QOLOxDQ
s9eDLV6AQr20gv+huVXMa23MzRYbepxrArpF0eRUnPVaU0SDO/+T/Hnqbmq4IWe1
yM+9tZ9jPf9YSrjyyZYFYHlzeTwqSE3LscNshHR8Uv9HGaswxkKxRn+apSNCuv6D
vFy44bDh6qW2TFIF1mfKVzG7pFG+D24UDzH90eXDIwzr5JzgJe6LXVC7cvIQEALO
/x+i5DYN1GApHi2gTQaJ6GV1Wy27vpGw5QF4laZhZ0BqPBXV2XNxnTHQHcagLJs4
+G9Nl7xjm0Zqicv1tmuV86IEVTZS3htw8XphQ85ey02dToUjalsyaMBm4aYBytgU
6tzRaWWFNUKTRR40R4krV1moMm4I8I88oSRznRYkEU/W5205lb4h5nsjN+nBiLdd
G6003iil611nPI0BVt6/qrpIZITrA6yscWNYobt/jLQZd7FEDyFU3vyZdpD5CASd
1WkgtquQ7dWpZBXdbWuW6f29c/TLQJ8VKMH2NAC4hk3VlGoU4w6iO850LsL67S2/
1hpquSIsyaVc8nqknye38TYnAj/fdtep6hkT33may1pKQBe/D0+PuzMTyLoKlgZf
aB+km32ySkJ7DgmJM60gMnesXOT59prAfgKAtZM2H8dFLiwByY3QGrii8LBniz4s
sHengs+OW/pQxAFFBZVvKLt9ykyQziq4xQ2eXeLllxKignfT01MTDYJyR06ArbRo
V16OJ/0IzNbdLmTX/dOmUirKOq2wqWsAGO3RXCRvYBpLNXOt/j2qd0kqMbRcNKWV
+NWyWBkGKqGoTxSVuguK9G3FuHBlVkM1Bq/2DrJ8ApLNb0s6furV/joR+ioebIXo
p0yhc7Awog414YTcC2FGMMlZI8WO+YJL2V8B7ArvEkxDG6ClJ9ecb3k2o0zGsldP
FpeZIEdx5ml0UN9cqwfL/LSerVDE3zaExcEIFCe2/xMtBmknhjltwUNvDZ45VFiM
wZQuI/yBMkeFiEUL4YCffv2l3CmmHNAhUJCbIGna2vyIiL8ACBDVbIqywNDCWNTy
tMp6EHaTUzQNSJAFCFq/8MH91re3rOmY/DPse9RVzcatay+x/G5dvMVpruGD96Y8
LVf1dI0ElODAMCY7pycfgoGAB6YiFDGVq3OKxkEfIICBp985iX8NIWJ8PKfEoDT3
8itU3zCDSBxsn1mlVWRNsuFOcxJ0Pp2l56hWrpbDtqPUUh+B/0MZUkhE2satzKLm
OEhTxoa9naq9ypa3R/2Q1Acq1aurt1eqjrl/Rv7HV0bRcTzLKvMrclPNeR1RX9Nx
zFjCEEtM88V+U6OHJxSVbvnEsR3nxv77v++DHh07mXyZiWBywmOahTC/jKxrgRV6
21vZgjWztCFLngsZNK+mUcrs410wRXFTQpl/GtzXVQIBGYdJETjBkzrMSkcmrdOR
wujVVmEprk/CSUK7VmjlxSRwT+4ftwyPgwNvkd0369UVEI4XFjM9uGDrgu1Yy2Wj
ibu+6cSle/7uHij3OKE4Wx/jeNzMAU+id8Rqemevn+bLZPf3wa5EDIEszEJYfiOQ
Y8mjQgSH6R8xnDJOXjfEKWv4WMP7uISroIajiFdMOEVvVDVTgYxVUMU5pKCPdczR
+n+ZsxVCG8BsDGbRSAUgaQgEcH6y9yYyzOX5j85ppHFM/Gd0svPknn89yCbxCPog
Pq7bY60xKJuhs9gDiHDb6+u2qlc321+qVqEdzBTP32314Hp4sjBRv3vzGUJQJSnp
MekJm0o5J4Ik39NVQ0Vdn5bMsMAIQBf9i0c5lyAlKH58IA0gM2YQt/l3lVwffifN
CureVSyxQM9A5guMWzmwOelkUU9eGuAfzwGsY1fJ4DWJ3pwHijiX/rh3kIYvbGn0
lP7cI9xZ7S0BrILT2EeZuqPZbuewVeVzaOADG/xYmq5nJDvPQQV2x1I0YW9VdnMT
GvQI1hYK3lTse62fHWGRi0lXEL30pcX31rwAceRqzL/lCIa2DzYOdb7AuOpyJN8A
1eEWHgATEpDEXI3tKX8hmwIEPt4ME7GnLxRQvlYAh6afCS0zYf+a+iCgfXebwTpm
H9SzzIX/qNtbvEN91xmKjW3aVnYCRiLrqcs/Be0pwrSNA5uMsaRmShnECMP8iaIA
T0frgbNSWJ+T7mP1VQ9O1sJrx6c2h2c60eAuUnUptMgO/n3WruOvZWYxSbaoCtN4
bweATvcnyh+uaXlYU6IfcVc7QiTe4aOaYxp+M0u6FUjXv7qBSXkHzN8aLMrqdh+D
MHzs5WqYZQsbZnqpNvwAU8wLwDpkiN5foxpE2dTJ4zEQAK4LFDNGYahTHRIN+OH2
2VU8LlErcw/8i4ts9RKJoy7KGiu65To8NEgwKEX5itI723r99b1uhkxa6DXFsL2v
/YMi1scHcJUydGakuahSsNOjvDRNo/oWJAJeII5yBg+xEKFKivmbhE+dYY29QfnP
oJQdL2T/cSysr3SlJmRk66MBy/YiKZCeJ04VHXkrU6kwZiir434tiGwcCytKnyFu
tLKOg21zWdjQGVLP5TYqrjVWhXK4JmJQlwGKP0os+qjGG7m1+MNcKoJg77pmOJlB
iZTZuxGJWiKnoLLoPaQ8g86LOsbigiPtdi5gir6QmdAZY4dwtT6zAV9voG/RYJMI
LS9pBykKAR7k0VK/kGFaZhrxe9D2rYI2txJ8gdRqHpTWgCc7DhJvVPm17910omGS
rP/GPPZkAFgl7Heqbl64X1YkmxcelE4svTn1Ra7DtqjpKOgX6Hs37EvB0eDD/NPM
qd1gBJ96F8093iFP5HumevT4+RJ7ex2PMMqh5zM2ICjo5Nruri5IOnpEtHKlJGum
SppTkySi40glcSejUiq8zJH2sLOKSA91L2eNo9vcy+Edcq71ocs3gav8I3U5ICI+
BZH/Kne8ZRJ23i7jNLB/BgkYzoiye8RLSpCT8WNRgDm5Ujx5FhzfhwnuNG+6KORN
kX0iMl7wiN3lSMMdnVSwhrbJAp+AEEfzBb6b/bP7OeGkKtzsobZPcii47+q8wPsk
sInr2jrZU1BbwLepg9u5IdMssKvJ/EXesKWd8nksPscHXc4sI14qL3Zu78r7vzQh
XjSuvVQSjv0QSyquRr1o4r6f3Uazu8OODmU3lfRkfcIiNwALCIPNZj6lVey6lQit
U6yUzX+esADyqPz3omBxxzqyAGuhGEvsqGHQg+VHKW+YrzlPqASui881dVWpS5Md
DYIthkqIKTqkr5Cq0t4grNjtaJEXqgP9kCpZkOcoPHtgmQMsLby/hyShksyi8CFL
EfcmYw/2cINpRTNkWanSPbEmLEtVMCXSo5wXfh+/VCXM/b/nG2Q0S6oLeiOnKox8
ycR6pQYKKkiWnWWbX7zGcmBrnRYdiEsyXMPtn0h5ugON/4GtlEVmOJnWoqBoF0Fu
w3ANKIzVX6vi5jONfIDgGBYyBWnGn+XaPP855efYLVCNFOZf4GWCK8FAgPiTfDRD
REXh+FqahOjaEs48BSneo6bw0SxrqHhgt0OI2Rp46dJ4Chr4fycHjiYGicRcaCZJ
GAPip6QcODrnXUkgJfl+yHmZbBpeeiU4l8oSAoLpcWeLs0c7T9AX7w2o3Q1uTTh6
mnoAgGRNfAjW+bmsyK1Jk97/MjJrcqpiB4ga2FvgNGzebxGi6OTc3yc3jzxJOdmA
2Vlg41Aio+M4fzKRQA8k2cbYkE0DdWPJxNlXu3qtbNky+cLvnBVNtLj/5RtFELau
4P8LiQlvrPkL3KqOyz7oBusz5Bq5mv7D5qDN8PnGZmjLTsxWHQZo+1eReiH5wf/E
FJ0LGqQBDo1Eipo6U9zfkjNjVeP0JToRjemDINI2qz/UqpFRxFzNpwVRcEwzj2Vj
TUakwbCuHb5pIfzkKV/eXiES3P38IBSG0hvescn5mgBFqGh+6og+BmWTPAp9LMQ7
6HftBB7UW0ce6xugE7ll5bNsLvP+HEfBEBZwbLgM/b4o0NpL+qB0/Ch+QNmMQSBu
ZaD4ddYDQWDUDnMh3I9bygGVNMNEIupQkaTNLF/YvmA3p3w4C02MefQQ1+FekFk0
uKJD8GrFbcU7JZOK7+A0xlwDJL9olkoX4+JR9oS1BwoC3Rq0uVPzr+4NiXXa4zq6
JUj3eRz/0F9nlgaqx+sEnqoRidUSJNIMPSBe+c1HiKBdKBHLHTtZ+lp2u4jE3Nby
+V3WI/6d8xvzsnJ+5J6gZBiYCLbe825OotwB2F2Qvl/Nt5ey9PRNMjXOip1XtOyS
GYHqx1tsOIG6YmKuxuaO58weDktPBndYpcM8k7etutffjYjUWWiXxIOMYw0Uk+I0
g4bK/W5/3skerzhMCfyZly4o/KAGhA2cs7YvQWD/2PYHBJ3XpUgCiJ2uziRKcnKn
95bkfBakBsIL2JCahLVKni7LzIjrVMO5txdPH+u4cyWoTyfy6fuEmryx08acfW6N
wk0Rj1+KeBZtU7BN8bzbMilQ+mvYMclPp6NC3kLTCJtBFg3ggzKY72Ofvfq6uoyy
u3AqB9B9HNnDqoqJEMd0RgnqgnO6MSgLHyyy2D7645baCla3dw3KOSfGM+G3zJKD
MBNL2sD7jLBxZtMLoYN1YCZPkH6V41F0D/UMIfNK+Ccfmr2OrrAoQ3mEwyaZFTmT
bNc3JXdVgR/Py95cxZSkRKGGCZZeSgwcpKNulREMmgaPsuX01rII/w1x1APoEokc
CtyvXLupSf0GGuIA0Q+SKP++H+tbmhlR+KbLLoIKRNzMS0FzdGHPsN1eWREZXTLd
7LOzoQ1D4tq1ZZWAIrqyUzJqXeqCEdbeL4wqoR9WTXxCEnzu9yz6DPKVb9oeUspN
6sY6UwunDrAhYAEGaBuGZBYcub9pQhKIvIcvPPs+8lYUfs4iNXn/EQndJXJp/4/r
LpgWg0ZQZ2uZILCUzGQwgZlU83pvIutUDmC5GgQRPwvUIodldfil0ZXWdGRzfDwM
7hnpJnKJzA7qkHieD5NQhEv7riXh3UGwziA9wsnILC/FErreOaUs6Yqp0lIvC4Sq
PiQqllMQp+jwsw8zxMo80F675gLTKt7V9/YAM7+DKnwaFicSyq6VnHcmS1kjSfrA
rUOXHrQCrtfr5opwN1vpcLat3npP84rO64/+X2KG8KL4w/LxCLxREcTKhoZxX41l
xkhOHy/v7uzoZ3lvpnzHsdwNEiX8jSBPMIu6NZdaSJVUm46HqjsCfpe945RSNCl8
OQbr5PGiSj2OFEeVZ2WPkcqMdfrwCh/veBmquq6Bk8RPPmZqtiGM86gqOBIuNcd2
sudkVI00lveWWqIxaywX9EMxm5Gx9wGHUN0M7pz/gy9B4Q9cbBYQhZX1hUjvmcGF
TQkTJrUxojdiTq4ITq11Ob8RkedON/JMSW9bt88kXXEBP9t273Zkkrv1wZQXV5aU
6997YYVF7HQtpO8dQ7luyUmFHi51RCs4H/TgoSsQapKhemgD7Ed3tsoTdSYIiOos
Aj5e6FLiQRdSfhGp4CtnKRlPbjAkqVoEyFR5yKSaKV4Ep/DJ9KSw6udChm/+hP8N
GTH85O7fLpNj6Z61slU60kVxSquWsEaFEQdrTFD0/V6D2uf7gpFHUP2PiZK/wSoq
QYpCQk7g30gi/ZWkxSMoU1zJsv0iaouPruoyGHLSti72r0yo5QlC7AaKAlpmeKW2
5aFXO283poWAKrKNk6O9SucwiZGm/7J9iqS+q/5I8YgEPZ0IU1Jp91UiiqXRmuUF
0xUofMAV4//2pTjlB1JiHo3au0huk7S6srJvGEUJZlUAoR/QqpxRV43xWQnZBuE/
bDH9mIp26dHH3N2HAD2H0MaxNCjWY6hwFY9kcr8MBU++1iKUrwXRUzFXD08yzfdN
hyImLdWYT9/B3UTTaL10cuwhVJZl0Wi7anN5t1WDY6HdP77znW7Z1tvjgtMZfYmR
3mdD8X4TJSn51FKD2z3VvMJ9pKfwG//D+mJOOLDndNjlvP4g+Hnvq9XHvJSIuzLl
TN5gdUvt/HEZsktnno9ALKGM4zZj+tm0UzQ69wYFIO4ac+mbypVI57RxeSgv1c9Y
xFz0jxcnYiRn2FFbz3tpFFEHF35yRckIDbW37re/aarKeP0STomIh4+t4S4f+rpC
gC33UtgkbMI2MvGfHze8V05ILafZyONeB5vGe65iKK+6OP8t8Vx3C07JczDW65rv
Yo1PwNYs+2HIbLPcowgfK7T7UwsM6YVONwR8OdI5DTxBDg8M0uRCdhA3wgrDEKx3
LJLx3WIROlVOy78+/VNP5Ea7HgO90qCnv1gwBJkYF9LfubjkDSrNU7/4Tpfsr90A
+4lTGFPxlK8rUSiZmz+scN+ZZWLQZ68TLdMBM1usvwYXGjErrGNbTCiPE89vYt/m
XiBxYhw0BThE+v7F4lejQPgKJ2HJSBQhhYssCawvslodz6vVVCRYD+nQ4uf/18E4
jZ7gSXakMkl9H3vxqc7Fql+A3Yw8ZaMu2Itgihr7Wbsqbdi5VMuoP6Ec8H9IiRaY
DDA7WYvmsH42uA6Zkm8rI+J6jr/x0VWU51hDIyecWH/ykywsJjxtRHBjINztroUW
nfcQzdGZyOuOhL00G2MmpujiXm12CcLusYcXjKfrAxvC/Ex7Q0Yy2q456XhOujn4
LZcR/IWLJrF/Ay612xmDaHEQKhnhcqS9KrOfo8puZw8YtsOozC4FXlU6OZH4a8TJ
2fb8pTRtTsUe0CdsAQk+5vq5uzgM5A/d3Aa+F/FWOJQLxEgQ4xMFRML8htQ9X+op
dqEIfzQUN7lBs5Ervq7GV4B9s/lCzunO5scuL8e0MMOxGvgKVAMzfly2JfckdJW4
S9CFc18XHKJCK4kfu5KOkEfPJFE6aQ6kAJ23nUtmqk8AfjouUIU2en9GjOCcN/4d
8Kj+ylCJIXvoLz/2podrvAjHhahun8Hs8jxXShdFggxFUN8p+pH3EtCnurvLNdjo
iX1oi9qTJGLMq8YgzRYaUBCcslp/xruOh/wOOxuI7hfnD1h+Hw/LBlsWDVc6AXcw
g9dooNd/60mkdnv3u3su4gUzmS2sFK3PeU5mc450OBtsvKCaEQ9lUF+pKCWzclRP
aJvDA6fQTUUTJ7A5/wwK8TkfLEVZq/X5S6ZrNtbk2CC3ASRcu0/EXVt3MagbOKcf
raxVqa+3fP4+Ygugid2APvraYmAANjiP5JALVPUiQfwpN3lD+NE/YNAjAzt1s2bn
A/4LdMOUTTFDgiEWxxuv57tze+dvVGypuaG4KzTlJkgbcWH9Sz6brjyJFhXLRvDg
7n6w2J3vwFkGreqMWP5vVYHfw0vur827P4UtYkMSCpq0cpcm5Aj4BTg5DZyfA1qH
4BqhkbCIhzXe7Rdx+T3GVOmcVqtmR2iCsM2mRhwrGiBKbu/SmOrpcnoHMzPtnprT
XPp3sNiDSt+Cu209lt4H3lvToYqVaQJSc5wAUjnMEThhKTJznEPW+9UHXa/1APMi
chNK5rqwqyKgpQYO1QbPvUjn5Y/O+gS/yTdNEs973aNvJUZ8cp3l4hEZEq091LGf
Hm3L5cM3aV4Y0VX87gQnuEixmB2+E2Yi2RM1WnHAhFdBI9UMRML0XmQksH9EFmLL
rQqadq2rMvKawDA1RKfllCBmZlxgKg91exl2CBbIAjgBxKtUxI6koyrPmhOi2OWl
/oTqvqldjtz4YlEDtSxYcMDoER+eUs1ByBP28H0ImgneG07jqnImGyCTgeFQJGwB
HEieZEL+GTTj8ZEcH0OyA6Lcoa0ZH/X9C7brIBVocZKtFWFjQv1kWvsxGZ/6xdno
oNQSNLOocA5IAmzSfQdFP1Wk3XwTO+jEKQMml/ttqFLVXs/mO/Q5EwhcvlPoIdvt
kN0wp8O6yFmTwvYJducYz/TCTRAORX8CC0FqnL3dBcgAtdKuhX9Z6VSNQEsy3JwY
j/qGEK2VvkpJQo4L9IHzhCjJxCYff/BbABc66aXOqrQTzmLvoZ+OJJj/LXdKBPUU
JVdef0duBXpweaLZgqh0FpYWglwY/zypaN7rjooRY0+fD76aKzgilXBP53TvI4gd
O9Hsu5eG02Jy6e6OtRPbsKy3abU9OEl0En1U0W6He0jWE3pjSRy0ic+n4OTpIY+T
Uae7iiW0YI3a5cNsKQmTG5vK6G6IIiAEG3zFrhDapFOyCVDO+wGrFwixGNUCtQUK
ddZRMAoH77BwrxDfYyR2YgK3uGCc8uMQV8TeHwKkF2mYpOFYdKrKGEX58jtnW9fX
e8ZIYLQUAXZhzDc8IIW/t66qRcMlYZFig4wn3F/v0GN3M/8uwDpl3UXrmdRFPzo2
7eLL8ZgtPl0COy67O9fJZmHBwt7sTEMG/QUlJ75KDFMllctjkvKI8txrO9FMGTQ0
zuZHNxuGJOq3rAbxZxEaVndvH1gz7yMYfLzsX1rHQSrqf9JkwTHRTBIf4DwXxCnD
yrtLc8h/YtpAfJZ7N2XZM9GVPKIqAbkMDS1BhFVKfZIIKlqdlXbsN6KoR9gLfaIP
M/d9ysIee4zItVurHA4Gq+p92W8f1e6Zkm3cEtpF/q+PXEzh5V/FQD1OLgBbZLj2
EljLQXGyWTgKigDGiuhdeR2Mn1vM8+6PAeW/4npViFyeNXWVIqrcDi5IdwiwExhO
3PvZ+M1B3UxKhCZc/iUpOdEd5rGI22SLjFPEtF48tsB/DXEhCUY4VOmFaAGqlIKV
2F8q//Y383EDLBUgm6ba41TN46lXeS9zFYF3AnYPRsS8/N2xL0FQEnICv/9/XArx
UmJSQQAdzT8c2eo28jB14VizGb86Z4uKoYruBcGnxU/z4ZxmwAmudfQujKdZorIs
93TtkRhDx18pj8KImsy1jpBROCPyG4lW4UiI4/61MDNw+y1sQvmAn8tU3irYfwe7
ILsoO8qNVpLIuguUZbVjb25MvOUd01fMR5b6R7/GT1tfEp3g5/0lqeFawBcxq7FM
ZkKAukdqfL7vVbHbvhEN5dgf3HcZM7PR0dc7/Yoznydm2srMaI58jffbeV8GymT1
vofkac3Q5LPVZyqJ2i8XzYK5SInnHXTh4zUgNvAeBFCq/2Nr1yXHlZ1T9t7E3+uu
LGZjhd54h+lq3pceshbsBNsgP13n868oDY23IjV42rPtlbXLmRhWnvExS0IE3akN
fT2Z8m/brBZrwj1RrEss1Mu8LWMbz7dkRiGilbkMnKHDj06I3ju6gbBDy6VQJYji
DegybBqnK7Hs7WyF56WXHtUSm/hK8K+U98aeDrqFJUNAMutk56BaYiTY6DtkjkOF
LkY7qofmHWf/s6+WOe6bZhZb7suwyATkqsArLk+K4ZJ3ZjWaRV81tPE8GDTPKKIi
DMay+w99E+m7IEIh6BPX84/IxNzfTaGWqDq8nyCwPMbhIQ1G1ZEYzpTMFnXKYfId
fX9ZsXo6tzUTQLDgY/LJu8TxU+ywm06Jl+YxRHXwvQh1ttTeJUzikuB9NKX9l/uB
WwhbzFQ7q/eOnFktuQIReLlhVZbTTiZo+ZkHLJMvecDyojxnR9Ryp8qYlVo5RLwR
FTowr+zY4i751bsdLoUfwWOah/gYgNn9HFNtH9FCseIj0Kx/Hd2X1ZVsXG5k5rfl
VzkgbEngBJfc/OES/5yTvzMBAEwak0DggG8XilcQ6y7t0ZlcaFGDDchYgeHSkNmG
OYQo3z2rEI6dzIJDeqg9TdWnXwcq7j9Y+6dtVlC1Ukse8CooKEwHBZR8mzMoHPdj
D6Bpi1GIZLBItZSnkTZDgbQH6KmOoABrZ752PKTApcwO2lwg4r29MEbNNQYs+ODk
5j7HVNPFKuJRU7tVtErD5c+9WVGRV4q9dpRl8+ieK2Vm3lgtOK6z75KjK/lsL0Be
2Aqy/uHFqAHWC629pxy9DO+ZWziX6uHPfjaKYKJSARwyzzYn9Xf3Tf2sby0Glzmb
EGHyp3g0ZORe7rfGn8aL1xc2upIPSPpjSzLqCpRuMO5k/VFD+R9IJ9x3bC85bFWS
Y+icnjS7X7aaPx68mIVsMBYRHFtTToPf3OG04ZR/jGsSr0SPNTFaraukdrSLy478
QNZi0hsyCXpQ//juLecPnOkJ8JjSC3fv5rinKhdogfnZMFV111fmIOk8prUAoFpC
rYYxPuINM4rrfYEsUAfLB9n0Kv7VxvwctqdC7/2AUVGmSDK+dAyPXKqN12UDFfXD
TMsI95jiIDx+FK9lMgmB7JMi+cTCT4xiEzsP0PxT7ZibVEjEOE4LS5z0Zq/E7whB
8QCsX6WNQr5HfMvS5BNWjzRd1M5jxPnLljiM1+lTc0SgEwr63NUlmRxmIcNO8nz3
CQ7j+CwO7+DA1yDQh9jurOzTd8firwrBMXVZP3awp64TxVsDzC1921ZMfLCUxSPM
g4FgMA9Jeyv3WWgjaAEWCuPDNx+tgnXpgN62oOeSP4FEq+C8Yw1csrJc2SBoqeZm
snPKOmxfKgPNktgi6xfMkGr5lqyG8ydEyFgutVts6zRKgg+L23k2+0QQhvYBQ6Ss
KV9vcuBRicn8JGBg68ed2wARodosxpgNrNWKvpjB82Kqo5m9YS4dJW7n+3OBs7oL
IbFqxxHdVdVgESBOIBKe8DT0RyeMP/9+R6JlJ4dgOw/KTZ6FwAN5gMgh6H/KObWL
k5AK1Fwxgl9nufYd7XTv42q990WhyOCXJ0bvtD7UXr0tbk1WMkSoUV1LT623ajXV
Y+FmAuoDn8L4DFcDOMnpNTiIKZPC+2LEeoyyUM3ZEdOuWu+C0IJEoHr+lxgSUr5R
t/nEhVVuIhb+Hz+pIKRp+auWhLGAdN5nVsbD77VdXCHTIGYvHKMDDUyN2nSGoTPM
OQtgki6FvxUwIOFD620CjAP7TBOV4m8tsmm6UiAHfYayARBuWSs4L41K+w8xf3eJ
7ajMkSSAdcBZei5wVGXXFHrXLeAmKQzxC+2IV2z/kayFOw2i9CRl4mF1aBqtdVJ8
67QV2SijtN1Ae1ClVgsKY2V2GO38U1y3hc4Vd2qUIUv1gHUjsBjpbmzBg5ygHwrA
FFG3Hlc9Q18fdFmdEWqefd1zS0VpB9ckSQHYnPk+K67QejZEnKRFkMbIjE9hDzCE
91OL/MFhRs6BcraOvBdmpKfkFqonDzXUNF7EzuuNrmYx8U8EkY49u9npYKGWKOFg
IjNJ4iPBG2QAg3kckquYjC/BHXCSNmKQ8LL/bk2L+JXLGS2tD5NR/RXAhi8Pdu0d
XhQRgdQ0mrKW0zQJ4kj+eCePaAAmQUkP3sqmUCsNXWc0+tMx7oVE9k//hY63ipWh
qu3FoZhbg8mKD/zFUO4kNs1JI/d4dO8a/mj4y3hw0isVrM2QeAvLZPEgi09ApWxU
KuRC4yjCPvjXPjgFcb/W8jTVXmsb+wKGL+WWd9lrzFWtYe3GOaXIj2Huc7O1+pmg
qsAPqIiMjSiNpSXiFywWzJt3YlnT0YBTBQBk1xijKQBBG+5CZAlRRnZGJDpDbKeV
QxJfAlDlRLRW/54cnFsqFjPRHAggD1U9DNBF/OT5K4b1FnufpNH1gcU4/qKRRjoC
8rakQtTyiS/UJCp1d9LMlU1S6wCswclspIrT0r2q8pRCkg6fT1IJglkBP9mWrrGV
28/AbDZBsIrFF40yCQWozrHxkx8RD5JzSKHP05i1MAKNei8iuqYrgAM1amM/l+tY
zvMORW61GROHh4H6BkMptgQEL/totxSUbx57HtWnUqLm8EUV8nt7YA/m8QaBTpuu
8RpQgMDhWaFtuT7TTLoc7Qy3CQpO8arDx22fsQV2BpG6NeZYD64uTgJrzq0vX3Qf
I3CAbevYo8cyXnO6eI+340LFoQORU4ZYb8FY7oKCB3AA7M5M1vx0NM1UJaPWJR8i
YckHI+ejsMVbXfUbeOaLPZK5zp45IPpXuGuOX1+KNJsDkJIAOWkI+gS+9yjA+goQ
y/kYy1v2glWkfMqpe44ymGQnVCBW/X6VnIAIU3EXDaOW5VxTCcEu8gNyYmjHhcsP
JLUeYx6DM9oezQcISkQPq6AygTcqqMkjX3E/eonC/taZYb8uCGw6AjeXTFRI75q2
rRw/IPiyPn8wltEbR5SmBFYLXe4HLBJWyZ24qH7gixoWtokBOj+ekdrOWV3x58LC
HV2qpQzmuQqGo9bHfv9mZgmmukukSfDHRHLphBj+S4M9w9xUl4/zokataQw+H5O0
CsNd7VRHuZT8fJuSgtE30SOnK4EfSNwTeMVdeYF6TULzJ0Y4FGrJMrYWQd6GR9xW
8fcmQBEfvv/nOGuheRjiQ4oQUdvHsqrOezMMSe7K+tIHBP2wNdspIGBJvZDSLD7T
QIdXggZ/bu6snWhL2GT8y/6XT4MU3u+hSMkOOGYQMuN+4BhfPPByMtmVSa+SdUco
QCE050BBNKvnr9BlpG0w1oQa5/wdbdxw4NO4aNM0SN6zUt2nqp3a7+gqhCQHZhx7
B/vnQmVRbAWrqQPqL45dnW98906oewAU947SGvjZdDi13MKKDEuDYNYCCC2Zg69N
yucEKGOq+fI3HkG5ifLTHtOm+KccNpH0th6zubthL4ZVBKqeEbE/7LES+c++Gtkh
YyNTq9+ExX3faScirgCjGpyiljKFAh+4d/YXOdxZojJwlqd2EAuaQsepg1uE7aKz
0NckByyHEsRCO3Ag7/ZKgdR98vK7+IFtVuwqRXnBdZBLWt1BaEm+JC9B4di1Ajgf
JjWgFVfMMwZqYkxtXT80CM7qja/dOIEjCCWj4xOftGDBQV7D690aVHAsptW4gIUc
GBR1JsbpG+PMtbjwAEjrX02ERucHwt3GFQIAvlTlj5LdI1u9BBfT22TvYLnUfI9V
K/3SDT70ofQRhl2TKBEAKbZr3GnEECLaQc6Z2jQuJeeG284vyEf09JufCPG6ID0x
AuxOA31veM1bBQb/a3GqX9jX9Rh8lSGyRPXpPf7dDepQrFRlQYNMaimWvk+v0MZJ
5NqEtNDKn8O/plBV6Q8KrVzqYctW4wducDiTf7HxXeJ549/wVRdXpVITMXBEuVBh
iCp/LYf3PQydB8G0UrJBfF2MmWTBbPTO4Yu7lZ7NeRTO6IdO+w8wh+qtTGLeyNMR
SJTtDx5u7owaK9wQi6lPw0CSHwY6cc2irlzBuypUKCRQ5b1TDNdvZc8Yjzcd2a/3
ZAgud8Vg2PTYZbU7g0xQGSSYO8h2ef1WZHHow7U86aLJczEq5br2ZFzD1CsmOUoJ
sk85lPAkKFq5wDU4WJdEuoGdXquAZ8Yjoe2gu6xKqBSO9zlBxilEg7SQm4jlKqcD
90IYA9zw22hN3GDBbKSRQckg4Ne+/h3EpUSUyAABwb8hc3Vvm0sn0uiokVMAdb9U
iptY1y/NXOEvjnP26glFKFNWAM7AMb31/RZmVKIzZhQAUzcYSECZ4z8+fcPeYYj5
jgGtt2emxMxT7sgCzF84tI/lJpDpnoEAhfM6b52nywIBur5gUzYQf8jNqAS2bjRy
lYEnE90ShauZz/qtkMmSZmJD1r/tzssaslqR0ItS1XcDdRpP1DgYRMcTHknjpC96
O17B/eWUCr2jua3PKJaaG2/wPHZYy2V9JXgq2svxE2pv8B/dVwJsIHVyU9WZFDns
T169e3FcFmg14NdWhJ9mycoHxv18WtpOSvHLBptEazQglOMEhRwvUg9geb55l6SG
6b49t2lxu+z3bUAL63hTTzTL6kCzDGGH5tbIm8Lq9+Cv75s9ozPe0Hon9hffO23l
YNHoZJ2YMs0bOCggr/Q4DxZsq/ex7atEaq36/J3Di4FMtVTL/62fPN+EdrxH4xCl
x1QBn+3SBOh072yH2yr3y9B4VFpsnaLi+5+koHAFOhD8Q7uWc1GiFYPuTXofcW6P
bwaLszMOPJG1KGqAMOUo0bmbQhZA1JihZEx69iXddALQ2nKJ2L9SL+tzueosPw00
ky93UbYsQopBOVptCAD8Sibg0vrz2rYZwEty0KZGyi2RpYcf0Tb580Tr607od0zo
ZNKCMtW2RcT1i3U/FC6OhDenSWgiS9TUXE0v046mZh4OdpVxbVmrmBzUQcg4FCnW
EmQXSON9/nvS1IG5Uh5zbr+PN2W2Px7/Qo3AyQqte5faSfcXiA3uCVatEP1RBnwu
87BHmM8YC7fYw2uCqDaLq494BqhQFBLvFj3KGOBj2HARWNcUX1AMGFEY45dBZnsh
Gn/PMxhGBrDoBxN7tfkyuVwOUxIsd2JjFld3mJIF2Cp7gejIOIgP1552Q+WSJQAB
31iRP5i9+AHwUanO2c3wo8+Fm7Via+uBle+VHljF9NLxcOnuk7dGkYcl7NqKHeTk
oFeCvBXg9SBQAaQWhATjf6q/999D1FJzk+nRPiiPzj1gdvqT1ndEsjk+0e3hJjKe
1h5WhRDIXNh6hjNvvgML7jgpJ6VqBPRVFRBPOrvjaepiO1En6uIAl62W453hpoNB
mIzspgeoCU9Dx01YUljBB/O6fHIXHLlswwREBjjwSczD9YVcCD+OG/BufN485S8J
TFurIg1QiFXf6y5apXghIvjvpc/JKq9gakEvXLlkTwusPRjKQtYVFrmyc21eHcLb
qedC6aj99rRceqe6r7SVeSDuhxh7R139ZEf+syGTXNdXOvdou+JAuYjEHZgnr8ha
VVl5L6C+8+Y5FRVZcEjqmIz0gb2WESB1WnkDo0RGVTJPbjNuLqoW1j15dO4P3o2o
lKtFuKk10wFL0VcLigq0z0MKw0zMDhNiJazOM+/SEK76/RULWndVFWVeJMFu680e
OXq9gCXAAfcBmEyrbfk+dvMz5g2T2JOeF+hpQB5DvvON+OodUgKYovfxA8vQjpaL
vr2eqnYDmK7kKRvPJWiUMuQHg6WLr20TMTD/wOhe2TP08if7w7B7/buUqipOVBDT
EhtUcajR9xwS6LBhSYWy3SjhTU/b06YcmLuh3J/bvMvKQu31t090V48K1Mu/0tfP
PS61n3D12Sw6x6ykXW1SQdxiJ8g/4pWfJAejbrMUZdytwg1MjCy9jjrtNlGEXkET
K/vU26ENoV4cwTtEWZwhjHXT4e8PQTe640G1TYIqAF7ZMSbTwYgSPNI0GUjJ3VBu
k/qi4/Z6OzxnlisUXWK5aqdqGV7Qw9rKZmplyP6D6q11GnZYIhqrumLiNbq+XQWO
A3M5sEYOTS/c2OrUqMvBsP9GHlZZ/36B+fLCF7TpR6qg4zaKLu5SHUjFN9m9fgSD
9mT7G8/bcazrVQNUkfRC+VAbHGYeFx1c+y3jK4pSkiUH0oDmXQdJ36ciTsrgTPws
Rc01jiv3OeXEKTwTvxR3R9u90tufkP0nOFCLZLpNtDXbllelNcEX95yFEd0/9+JQ
YRh5IJQILspLZkM1ZIOs4ZcNpZoOJo5CyAR8Hk8RwI5thlRgaezvSlsOu9D3tzUS
LpEyGwvNayK4DALDhSSTQUBjnoSGHyi+5uMwF+0kGnoUla6wVZ0laupDMo0SpLME
LY91Qu53K2VyTy5pXVrMq0dwQfDPxdrCJ5kro4n23q3hZDl1IDOyvMDAPCZ5cD3u
YbXC8Uhzvn7je++D9/JRfa7g4Fanwi2+us38T1TAKaACLPN1MWHHixo2IVq9aXJ5
63h4peQslBbsAFHAMw1bkrRBQvU3pwwF7nuebrE9BpWLTwcn+jyQJOZqXfeTpYlN
y0Djq7jMI2vbP/8a3ZPkb+NdNhb/cfEngHrHaobfdD+R9v7CDwLld3t/ZcTbgqPm
mRiFMktxHEzeUgK8t3+S4msr5WkrPa7mR9sLMXXOAshm00LA1PL7sTTQy6NKASSN
RZqtexS9trQo0JaGcU06sE+Uh5G1sU9DlRkk1kZZiazBDFCO3ievmn6f22/ibhos
RF7bN4pAQloOrCEGEtDEc7qdZd4iIIpyTg3BdDqhTaRAKOBUTlQzGsxAvZM0KTzv
QINGlBdxp5V4TOC5hDfR6HMoN+DSOVoUbPWtnruGTzW0uF3fiONNNHoqe2TnSiFQ
xEXSjOZ3EmYpKtonZKN6PIUu2oJOvx7dqDTGqhabVAOWiH/dlIW5weA63lRbvF5R
SpI3dnZFETFuImMx5Pky6DD8/awabaDYFFeQ/iwqcxRXbHfuUSAim3KVICaY2cZe
KTtxWMft6ykCdE67N4+gxMp8uICJmjVT04S43UD3VUIaqLo5YkGCDLLWLJdDjYcY
q8G710Oz3M1QAiBhOznrdg/7IY5ptxvBAmmQYaBGuQVLF4oSqBxgVFzj1yC08uvj
lqpMOLJcUjOh4g3Hu7LblMk/YlHkvd0iHNVAZa0snGjwKJlGDlikSoV/wRq79GKG
SKAwETKLHOGakIIwZ4OEOS2tGtjfhVR8Vg7W2MW5Doo2+As38x7do8BI/yLni9Hy
9j8bL6RcNuRPIqS+0J80ql7/16TbrAcRQ4VSge5+c0mvVa1i6tjZ9SusZINspRAU
3BtmDsmoRQZaH0gLBkswyPp8k5+i3f0dgmr45B9oFyvwPUVsXiAq7aaW5ThT9oJe
GFTlqqnhYm5sA1PQl+RFOtT36ih9Tk4z841b8X6LDGu4sWqs1k6eq1NKKSWMloei
pf9PIXMUNbipYpBeC5Wu5bp7mucO5380B3fZ8IydMPbTLcQLDjqkJ5putMWlVu2H
WuSnudAzeRvPcb2PlMQ3+f2OqTuy+q+gFz5g2aEbWacGe9RWjTYX2SrbbVMlwUX+
QeUtcq+VxluJ+OWEWydbwWfWL+MnvGkHL6Xm8T3Kytgt6QLimhekVboE0oJ6bq0+
DE9FTsmscrn+k4hMEpfoOt65cUbcWgSkaZhgVHrxMR9KDCnZJ18lYjmtUQKYj4Zs
pimsL2Twdw++cMR6IZXT00ELNrAkmD57LbC3aANxiWb8F+1bctC9uT+HijwOtFw7
0hMWe4nsVZuw7lVXYquGiStdATAFk+xOAwkqf+DxgqQiCaVTxsmOIIJ0cDRqlE9q
4zCk7EJNaT90yH6k2GR0P/pzy0pWur6CHbURgydMuDrS+Ir3g6zlSOm4RHNYazlI
1ua9mwxq6pqwiWDuHKbg9W40DBW8R8+oX+bH6jEQJAxQObvZRM+InY3g3mwgUhl3
4LNkytmzdWz22qrUmoC6IInlZih04BISM0v+IPg+FV363kZvnJ3DnPmnqyWLBpt8
I+BeItQFWCZjFgBbqLcskHsOG7LHwFqh5N8gA7xLSrtHnraKLx42p3FbKNT9QIXi
XUHxRhkNZsdxOHf6jmrKho/0dJW1HtZqkrhMACydSnPnevPRMWGSTOsY3rITpw/u
kNqNZKUXxXKnJo7kMrsxZU0Q1aCNCxFOQjvEOoky/dXx1GGZVdCdY+x0+vCIz3Ke
thZWg67piHiybMBzDvuUSTpWKTAnJnZ/ucmwsLctaQCbwf9HV5I24232uI7ZT592
IX/6y5Tymy+lYcAUzj+1HCWKLI/zVip1Qnn7ysz+MfhGFVLgSX3uMllCChVufQIj
DfQJIxDXAdMxjW3heI4Z8yn9aWkT8rEDNKCulOO5nNUHkLh1D248r9ATAkB9SthO
3aZN9ZFCbmKmCGm9tUNfDb0ARau/8+Hjsh6GhfMj/Ir3fnhfWBYTBcEe7FD4XQ4m
u1Sjy+yctOvYUtZgeEn9CE+V4kpvipV/Jtlxj9kZQHhyGvzU2gxJ4oFAuGxlyJdd
kPVqnoNJlf9W1jMQJ/jTdOtuAsQDhGsn+6aPI3Kr+fyra9vqnACrnk9iNFqscke8
oX77e0y3Xhse/scd9R/IebCQvOxDShFkxdKB8QSM+QVuHtAizIPIXgiCkWC1WvKv
3CdMPsRnnijLDWWXkAMPuE7duwWOIKBUXa6Bo3v33I3RomY8uiPBpmG7ToysJthp
1IPkqARcpLMKTOIxEfp4IJrQ8tr9yAvtbekZrH+OmtUG86T+Ow1U73Ao4hGDiR7l
OA6K/B1v/fIwOTshtnC7jlOH0Lxq8HeLOgyYPp+QeFpJBU+D6p+DLXN5M7vDgKCO
DQ81x5FJhL5TpqH2mnzXBCoXXeHWcEMf76xtc8PX1js2C5MS4uaSTWzhfOaYU7UH
Hl6VTomA3sqXlnWwr3hP8TZ9kpQkuqEyaVzYky4WxpxJNxf+lUDdZL3GL7vs5RzL
xBrMG8ZZsIXJag2lHG3+RSBy8vjs6bxWEoXXR6VmMofdiPviO/k4IMjcJMnQApd5
vSFR/X/JDdi1J7fh/yDgDc0c5p4Krnp5ikfPud40cNYnzMZleHsVuUtNqQKQDZjo
eB8wnnfGiV2AbuhF6yhjWZ99KwBemdhqgnzCDC6UiC2bSby5yke8xp4kJ/mVWtzK
MQCsQWCwXiEOqiG924pgVtWqoulLPWiNeYXZ7KejdAcBdfj5dNweC1ninx9rRz4a
wyWjQ8epp3UNkpuLovzm3uMpbVa4P7X22qd61qjzErYUgmDBzlnY4RkR7oYELVgQ
oKWe1VQMdIshNKx0W4vFd/utpq0miyar1rA5Ztrd5I8xWOpSfBE/DLsAKH7IiapU
Fb+pdGSsTKAzG0Ry7zl435Kd+uVqVFCfGr9cakT04JEyFv5EXmhndVet00DY5vXE
dgpFpJZdQcMmCKFX9Z6b33jpI7uOBN//VioYYjH9SFxhBpetAa+r1+sKaQHeQAVr
Oi+8iEwTEYnYMYFHttfEP8tRNw1zhIot+GHMlGDDlA9F0M3JlV9xLJ6y00xcmQAR
KHmk/gEAGDkiCBRy9jV2tnKzz/6Mn4iU6tzI0eFg8EMhwmzl16jCylb51y63MrFb
sU23XhWJMr8iXYkGwNP7HaRHN2L44gnRqDd7s20LwQoHFZuzJ+PBPaqguFnF21E8
Q/md/iL7oI5zawYEfE+HyJaI30TgSvLxWC77yBo3J4FMh2Ee9cQ6GDnQ4aSJ8sO9
6Ir94J6jnJO8d2u9jyYyuzMP3qcTMHWxl2mBjI7743I3SOz0ArZKIJ9TcuyRgUH0
uYphfp0BuMCdOmY6zIZOwDGgxPCoAfM/VpgJx2XSAIu5V5TXU+FSntDwhEnBST5i
oiPg/NfiDthXYLZlOHN8+XdDgjF6fVzcMUuIWMX5m4Ny6YB+eLiAroTBmpQ7au2q
eaOUj4ajVsuhrXjdinHVvEE+j1N+2rmokSf8vXgLvnDaUsUEeciHSTfPkBCxc9jO
yibvoM98sZW24Bb7OX/2oQtzLgiG31C5autqV1iiN3wEujEm3sxDDXlCIpnj+ak2
Z+rfcw3I1YkUuv3Z3mJkCF/579Cuz87tnQkCONkqbBvtSthyrzxSKNd4uYfGCUMp
xO0Fy77dGlNoRdlMyAzIOcl3ByknJtqp1ISfTNuZDEhIst0KY9VmnZdlTVpme3KS
jIbXa3HD1E41x9garilAlmpXASMYCOU5aGwptte3KUhkPDcdHgy4TyggHojGfSLf
iY+D2t9H8VO7fSiFWGcMm/1hWd8f7nz5cFxQsvB1cn4EuWdwJTmkb+YwmB4LHmcs
fJP75BYWSq5q+nLoR8nhwhBIM/jwXiKtqSf0Vp3tdH5RZlVJm/6LHRwqsEu9nSWZ
K+aETux0ZBE+1oCk/maWi+CX5TI0/mKXVxfHCYs9P7P49ECTZ6AGf60E9+TVQZk7
r5AZdIeWAvV6p8ahNV6NyQcsv2Hyh57WaD/TUxj69x8x1ZHVX4ceyhELTRKPjkpp
R3fcBa54/+BCoLsKBD8VY/LD5gfqerFs8IgXFzMtsxHum1OaP26fvosCbk0cgO2V
4Y0Wm98/ZVFMQdFEjoCplLNIxEhaXlDRFhMI3z2X91bXYs1S2+W9tZWDQgeVOsnY
CqcoUwvJpa06SATfLweQbxsZrq+RJ2mi1/tmLe/z5/pf3q8VSmPREA1aYMdURFI3
Cj2NzADu7VUPF+0T0hpSCkcf7SVq7v0mUXe8sVvEmuPpMk5P3p21ds9BdhceS8Ai
PZKMNz+Ma7DVZs4To6Qc7Lj6XUHyddfSv5SOPSSgh31jpUnNn8XnUZH/D+FzoIfi
4HCh5woxNQvXQypoxxntNdLSt8WTs7DPE1HKaZbo5u9DJMmBeS3gJL5/CzI0GwDe
+mfVS8topo0a07toGNzxmSsagzY8DnUAhEDVMC/7J1mJ+W5o0ptKxk2PNh7rCxSq
KMD1n0ldUUO5fFDRYak4eB3MqKDRVQQ0NQ3+lNDa47bIKe4cFSnDTW2g8L4yxWN6
aid5rX+v3xS00f9rZ+JHFJV1kjpSrgGrY2279MaByjhZyj7hCdVdXm7mgSPXU8sS
ywAfBGN2gy1qaUcMsoNLGTitSGZ3W6B/tQvbLYdz8l9LNT9CtCG5NMihOo0BThWE
Hmv1ATIAax5HDgHgN8SOB9k7Nd3gZAFdk/HNgR3IKOXgBLGjxzjiuQc6LIzOgkK5
n0VUicAwlfA1s726FFeS52MLFeFAbV6QhKVSdy2DLh4+DrQfGCXfJlBt69qmeHxV
/Hv8qJbcw7kH8agBDiFC7xqjyU/ykTJiVWUETXczQcyB00IH04sxXPPJI1+gCQec
cvRbFz82TesM4aAYMdafpD0f61aFMiYMLuqNy854pqsLegKvXr12qLGli8iRYlA+
0aCkelK8Yga8p5ZeALcp6fperJRuavdWEV4gFvCUsK+9ibOrVuKuYrw2yotXKn+A
txydNNK83iFn6APt85OjpCGO4INEoXoMTp/FHUj1865PahbRh3m173f6+PUnYbNZ
i51D1XTgZRZchSTLUIDJTtqZRAJqpBRvfuJ8ry78uqhOIxQ/CujWqdsSsk1KJ0Mq
hyGjRnWDvvTy7BwQmhhSE8lmyr3dvbwE6Bowi0yqOud5C/C5W2hCo582OTDt8Ui0
nGAZlRZDHO4sahRFs3qmFtcK1nUljMavovGWesrwPLtm0+knQMCWnB1TjBJeZ3sI
1oz7H4E4eUmSQZgBfK+aANDl4ES26ZQ3iwndP9ln+mAxK4O7m3dnr6q+JMSImD0D
4xCMhFdy07+RO012SLIoJ0u9YLh6Z50+AWW8AJ1t5mltBKBWKGPNK2W/LPSlosGm
RcciVScPaNz+JXthlZEwYiSITAfATTDmoIjxno0nJ2bV5nvsuXEwB/o1K8SEtwEd
VI5Mh5V0AeRC+jKE+CgtzJLSyZ6bLbF5DrcfoRkmMP8nfcb2PyLgRhuBRkW6lFYP
DahQCCgSlylQEh/zIzseqXjC74ahNsJru6A67Rt0DqfU7TJ/GFbcsixMJB4HseG2
WkwKEBlewNRWGwRq1ML+s8Y+jSwuiclxwN63V5PECNV/p2Md0pJyPHRnBWcBdNI3
aTpeZg8a/JnvmWzIy/Bo2wVPJmw5ZrQb0heOR4VY3AkrAWDSpBCzWkC7xw8PRg2I
6DoKatyPineXS99p6v8Q8b3jXde8XE1jrQo3f3DkKVrSUwsPdKb2W4lfSe/nc7kD
S/zIBEWsvaOBL+HIkdF6C15bdJsWjSwJNG7XBavcTSydBc6wAnLx6RD2dTsL9e+N
JeL7aVds8OuwNTcZFT0aV97nGpt9Nb+Sn4RGknrO21jBJb+MaRlMbghQSDEMVlyb
rYP/OOaj+VDl2GlcTBU+/PZPqcoJMBKmcGLCtmnj96JRqNGPDua666oT9JlyS/km
iXDegcvTFgJDzsKrG+qbIluqACwE6bWFrDQTgwqk9lt3Jc+o1uQKyEMOecIMB8VH
9JlY24iXaOWzQyn4SEsiUJYS4wY3fghPaMhoFm3++qkCA14krDfCcASlKNiQsXYE
B5+lko7N6KxPGX/ka3UnvtrzAxJQkUg9XKqzjwGESzk+s09Ud6K8Ym/PjpM0k3OY
FoTMmrkw672OPnPCVVqkiMLE1ScLOcdF41OCpy/D8jKqR7k7NprU61E7abT6juHK
tUpnn1CfX9QysVTMq6JOeXjy3IKbph1aGm5tryFni7LaqMAyYdp1+Kb17l+7h4BN
O5iqRRwxeuf3sIEcyTvwMoJxencgUXr1YrVdj0dIHulA+WAI1Lp3GkqX/rc16fF3
6CArU+nIR5sTnSnNXHNv0t1YQm3aarWrD3iEuWUx3ne/8a+lJmGb4hI157Zx5+1O
cWHvOLR0IyiGdQBUSn4jv37vtAJWyUAJgIfvaeLXnOSaI153Z++HWg5CSlHq8lS5
R+1B7YZ0MbqqF5laM3B7PEA4ZgSurdkkDWNW2SvRnPM1V7Uw6+QaRKdQfdA+zyKZ
YfN1R5yCezPOtWBh7B6L9YoILPuTfhT5IyLvJxcL9x//03zzsvB5QKZNpyl9Xnnq
Tu9VgvmcHA74d770nfF4PDyOzOYSVr+yTkMj7RolB/O7QhoRukV5BnuK+44di7Xt
puW+otMr7Ay8pIgTL8I14AMYOYYDId/K7Bz+Y1cJfl5DDvmIUsyxss5RD9Cf5lCy
wThgFrpWbV6zu7lDaB2AC994y6RLXBvBDDFONzUy261aTa9kpjOX7jEhQCyaTacI
V2/No/CWPZB7ikTJH9eTaJz2clsevQyXeM6KdoQ7tTJx/i+imgFvhGdHCygTTm1K
+BPoxytsKAv0yYdHTP9Pshr6Q2JPkBMJTtRQYAmAlsaB+BBof7sppuLEJBKgVUVV
nVjIsB6RWP6tYA54qRXW6HUQRCMAIg6jujvBAuvHGOkA1fv5kOcKUOdTLkPbEa7e
VM6+gcenSfbdPp3qBggh2Zx4q1wifyihkZgBf04/YIfuev92McCicExpzq5XotLc
LccOfG2Og2CjkDO6jFhjMM8pSr/Bi/PYTenoTAidfcMeZXNw5uWXJAmXjCnSzUrG
gvR3/0oGi2n5KekI1wws3L0q50a+sMgsEIRBGW4AUYOb9Dnj/W5qGhxZyVCge8n4
YoCk2VsI7gjbZDwUSTtc8eZE8AX88nkNdPUg9XOk/JD9c8uHNV6PI5u8C6XG6Gld
3HjOXbnTkSdCKHOEPX2ioKLA/XVRkwngc5K8yAdgybcCSwf3rnLIi8osM3PZ/ntV
f/7EWbdcaf1KfQaZ/yhrkZGkm+nLL/UuNyh8Xioce8J0NzCa9Vnb0LX9L9v83lyw
shv7yhHsCvsPtd61UIeCSu2E8FvqWHh4uZqC6WqYp+lELULR3rrm3qPICQtGJ1qv
Uc0gZ41yEdkXrWUXADlI+V4t5/NjQeUSeM5fjkguIu5bdMSpA8mqrMA268fgAX2P
IrnDMpORodsZR1Z85ffrAEOdMTHpwBewsPMdhdA8xN7Z0hDf0pwzJ536gsEsrMbi
I7Go+dRA044og/yfpNON08F6OoIhUYak7vZdll89r/PrHx6RgVeh58Gy54N2TzoR
9A8aYjbJ/cIu8vSfrnDZNMCQan/sH8Wiycl7ZVWScgePUyCojOuZIIVEBt9G/yFG
G72dVX50NyEEACrg/FPtgvacEI5K0jlzJIZWzipSGWY1gZZyqdoiaZZsLzbac3+4
yQLsBtMDU2cA/zCHaEEcqFzJykDjyv0/JHZpYSOxFe2LNk2kNKlgKDmanadDThET
GS1hAc9NwclMx7+D8Y4J2KDN2KHpSZtgFN6YOevh1P83h1C2KmT1HoWyBLd7lWeB
vGvTkxdzfQjQ2BE/jiQ+Sn79wWUjFnYuPrXFgNlvENiVi0ksqFxZ1g1+EV0v/RLe
jpemHJh7r7OH+TCXIWFeMuXHpE1YjrbKtL+R83u+ZXXHlo2xw4FE53deuRpRgxNa
3P2mBhBBsVZ9cnLLmsD0se5lc9jU9nns072nIBU0toWkst3SV0pmpsN28K6HHAd8
9HrC/BnYfKf9miFBQf3OfWFYbbLlTxg4kzakI15uLsayDcossV+hlRcLFsacyl33
I7OjMl0S1dhJZCir2YNZJs7Gac0C/kas7JFHNdSfpJaXzOB6KAWEk/rNcU/20eUS
PCzbinRMf3yutyUFOU25zho21yaop3pT3xI5LKbJkmnyFf3t0SFIHnzh/Fb0wHrE
JLkgToZxgu+dXkT50ClCiH0Nj+2ku1eG0VmLwENd1RDfmpyYO6xhLwSlVok4Sx2P
3lFVcseX5niW+P5qZXwVw/GgFzcS8/7ZTZh5jLPZbWgdKA+mqQnLdbSUmR6bFj0o
0uGWr/SANc0s2rLqwkctSnW+k5sOu0nmnTft5UM8rOx8y7Fa9Mr1HmFDL3Q63gRL
a6dCJxWvdVcDk7ThxXRebZipK3riPZIamVppRUkrCDCOWvKTl6WDYveP3HUnbXFn
5h2sLl6mrZYxjEGGE6qrdyk+CA5PIDRJuh0s8pu3NI/F0qL2dS8yB9D/98Xsm+9z
Vat+3nNoALOJLJCiUnlAerblr8lSM0AVTFRUeYzKVoxOXW6MSEwDH2Iw9OXutHNF
2RjixTGgmTIhumn1KfyvRW+6LEWsHZ/1Ttn7pYQgcnM7KWCy/ZsG9sH1s/NZKPeP
0rC46JlpFadEc97ZRFlbdHdkfrtEcvGyr1vXSdbgspXm6hMXIVaXpfgg9/Bk2ux3
qL3whZ6Ngsn81vgi3EHt4jq+VyYnrGi3VOf6Y5hkSiBzRDK89AtywEiz3Vbn+YHb
CM1dzw5bRk0xFJdu69jbciM5iQ1lN/iIneT+o1d95PoVyFMJIt/9ozdWLodE8IFM
KnoAhRIrwQpPs9m4r7L1KGfAV3RLW1zhMvqDtqrIWgj9wVhijxzk1E9RHhI6+bXS
uq7dNeZgRJ3+C8wObgQdp4XUeZ+Ptpv3D657AZdvd7gU1oaqsAPMbqSYwdo2pIKT
u0+aw/GmSzH3INAPxR7Ee2PPU8EXvsYK6s4evVCYxQlNH9tv76D4tJuPbjc7iejH
yOfdLokQ38PE1B6BQpATLqdif83yXkI6grlerbcKUnd+Klq9t2RRCsFGshz6vYzg
w/tQRyq4i6iRG2esG72I7aoCcJxFzlV/AZZ6ov5VFk6R+nEKp88rCrNge/zIAVJ2
9EWA+jwiZ7taZ8xTe7Ss7xUOsG2oUd81ZMcb4uQaa6FFvvBGxSBZjj75PMqqI8f7
eVaovkwwxkZeY8Ex+2uZNWvl1HYcYyBWBQLzJs2c4aBO221ywCSUo4mkH2aAAixC
XT3IvC0OsK2GlMOnc0HzX4kQCoMJzrJIosKtWcKxa06INXX4QUgeaifsuiW19I8x
7QmlgdpTIx2quvLaPUrhhRnegCODz+YgyLKzqyP73yA6F9bKf5+S+s+qZfDcpu+k
yt7hwciLzDvFd855O/rpN127xPFgbq1V1JQQljtjS9W8e77N5W57Fb/59+3EcQTi
jFSBRNamWUVe4AdI2daYgKQWY4pABrPuZHNFUOuCqKK/6jFOnaaBZI7qWNusZRKg
4gXukQdTAbPWpvY6+eTsgS3Siymdv1NL08NEc+WGv2Vdv5cEF4FjFIP6l5aJS95G
tG0MTeePeWBriUpejb620i9QGOGvuEQpmndJSBiMsOsho5OM+qZNQFNcx4ea92vC
zqwiadEFFiXkDNHaa0bYBYvIeCU1TqXd2E7qmusQjgUM25wJGnhSRlapp8eKDdgQ
alr0NDNxakyG0nY7caDRJhtmcvpyFgXPwfN33OLhAu4A4tKaeYma/VyjHyMZiOVu
bOBtmBPUMFbYwBh6C16XpXqFv3ICZJUMxTwoGHYlPkunecnT7H7SbSleiN2ezyv1
hnWZREIhLzOJ5yVvbQYCL87J7Zwz5Ck2IHmtrHu8zXPBzVYSVyQDGCLHoIpDgP4v
jaE5YrpXC0/Q+ZcziJTvrrRB0pVExjqiv6GtW5Q3pYBKkud6HT+XyjKKNoo2rAA8
k7zqLWdOiKAB8j3oopg2/wig/nZcmZ/nlxh1IfYmH3As3xAYMHq/AdfVKScpV+BP
z496Q9BUEJtOE9iNQTn8/aHBj0io81sS5gTSH1TXOB2TVJ4kgNWU58NuU9bdSWZI
JrCGh1BsnSRb/W7tcsSFDQjQDos2kv3WApKLZ3rZ3ZmAcuJFPlhEPRslMWwyTGCP
wuzi/r75acnBylVJZ3zs45YCnx70AHjiRtzQqEaqr5AlYwDRR/0VX4PEWMgU0Csf
FNacN7aOFohAv7Sy+ObQk1piT/hs3jASkWfmelV3ZpinJ0DgYp3fXD14Wsoy7Rq/
AguJTlWx77xSMLVk9AcwDmLJlcFPFc+ecVVERVeHHR4VOY9TQGMx3v6FarFssrUu
ft19a7Wx0y+RQUS9SYtKMrCaDMLRlv/qW+GWAT0VEtVlNJRaAcfYhF6Gw5G8+K68
K6M+TbGPfNWV/NHb+EA1oWLePfVpYlE998EwrwwIbZsEh7nTy9UHIDhkNLPmkxxk
xPXrQIfaOcTUm3YNXCIaA5JqpQij/Pdcyj04qMYBrdEIe2FyYA6a6wuYFY1ljwu7
+JBSzGXza5gssFalAsUFiaVMRGlqvqADPmOxqzvgYCTbynJdUQBiVhyf3TxYzWMP
GoXS4/8RXcIyr/ks6HROdE0a77iKSoCENjPe1en1iaoUh8zBqj866RXVMr0sZhd3
lb7BNcMcssdLz3kxl72kzDJEYx6u7WlqeT9rvEtZgZLk+O8HJY6zjRIw6CipnPdz
uFvdIgJSQa1cX7eOaQ3tkIPXIF8tCjleD4p/Or8fWrwxYxiz+P6nkkYWf/nY2QIE
4W2pFz/tGusD4i0rKy5Wcx5AYVsrK6W2dHkDM/v13XQW5KNKk6oHLKwQ1Ch82HBR
0W6TDqLVDRo6LwSEovOp4kUR5MtiNH6FHZJDFCYLHPnXcG2OJLOE4OCR1OXHlD5P
dM+uyu28g1LpqUkzk4Mfn38NX6mMMyRZ/ckobOGuKYHfSzzu8H/mc/4iuTUPBe3E
D8s/dbaM3iHczM2JYAWhdPAEe8T9tTQsHvuQjj9aiMvrYj2Gxg7FM+OguPPLRqpd
nA4pfy3V4SHC3bFFUJ3Cn12xOrGbM0EYNireA7yyF/ip9ain852FS5Ub2wbFnDHy
OYqGneben2xLU8qB014MLoAPdDf8dwk176pXRScqCgNfRS3/S6xvM9fskjf3/Lg9
Mj6WwVAcWBfKUBwfvBuJTIMQM9iRFP/OsoHx+jqqe7wdoQ9bRhKtIXM3JgUVR4WG
cN4LvXM/G+zR7AlE+MimdmjXyU+NThtf9Jmhbv4ReHuzu3PWE4zU69B+g+7i5Hk3
Qnh9Oi8RsjDzaeUJsmDwNEBPmDCqwScGFyHDlZdXc9kdKegbCfwhNC3KhEkBUljI
7iLXBm580SAK2bChBJBKE+XIpRIsNn7vhhK+xP3lzTRS+dEKeWebyCHHNWKiOVH4
+WAyrQOclpqJGpma2l0tbd+FIgNqJxgdx5J9I/U9iqw3g0DBg3URxLeZ46jgThKz
eWiN5gS0wYC3qAn6yS7RNB7Ym2D/oyaLmHipvGDLqZaLA5xJCkUsdwAMHYg4nE09
Y1WXGmLCBAo4j/lIreDGqWRFyHwHtRw5fRMhB9szNkMZc9yV9PySU2rqfqiYNzwa
fGMfVOu/EGuhRoruDnQCoYGSpmTAl/m3JHLsJSpF21hgAfHfAnqEA9Rp8vSSQWd+
XJOW9VmyC6/f5kOSs+pFcd14Q7c/qkZq8L/A4hvYFEo+Vp9Xp8FuOY8kZILOVBAn
ACLDIwnugcjQc8ZwURTMo5W7J6v4s6LZWY9MjIjLZ0h01Xuub1cCS+eYVsYMHi2D
J/WWqd+tl5RPlvVqc3QIp1B1piVaFCb15yvKXCp541RFtx2QiQRa8PtSFx8qS4i2
xoNPs2sX5Pz5U/tAEWfAGmK/MU1j07yUwZsel5NqAw0a8tie8Vysz1VGAB9rYc6o
iRNmmw3tdTwQ3d8EY4p9SAM4quNEHJu64AG6fktVMX2y7tq3vRZ4pK8I8a5IDL/+
kNOkkDMLuNEQ9WSOyZmY+ykicuKBnepsHTyx+t5t7gdrn/pKv91HRI+1IhsrDiwO
UVq22iiX811Ipdi3kEe9s2UOoF7hrKld2ySrQ0+hMj91ED9WvmcmU4W8gki+U3FY
BVIklyA29yEyygQ8I4N2ado4hSLwAgXmI9Uc7mc82OEtD5o+6ttLjnP4vtwyUq5t
w3HD7feWj1U878oRCyUBfrMvizkH9gwYuvg7AJrsnFCpV/Q7uAEXLslbU1Z3uyyh
ZNngV8UnUk/MtbegOadkn4Rk8e/vpW4kUFo5VIN5OtVbYFcHT10Xicz1abD44/QJ
9GFXiJknl6GIrM0kENUsj2QXui5/SXu/ILL+awlqnRPrl3xTIROPNTaYFYKC+7H6
v517gBYHoY6dXdkm3hpvlbXAG9W3jEYPUCw+C4uAwxN61j5Vlu0FbhGxr2lDa5bf
csi5oJ/tPeCU53UylFy83WpJ0TnSy5RXQCpI7dLzjk+q0S/soDgjkq21pRSZXlDq
VFI82BKuxM1Q/y0u1j8ZWgg1vEcywhoXOUpPEhtRL+HUS8x+DBaLq3YrJN211j31
pVazm6Dn3KlepCm7gq7rcCgiEHpqUduCJrngO2X4SQPNHAtc7XBBAG+Z3ibqqtRV
Qh1qIn34pEnwUXkCSNny5MeVGlif1hmpV4iip3dcFniBq1MUHi58JxESezwmIzPm
bWzA4Eq3bgbGUZIowiJk/aj1hzSe/GE50MvABeWepqIGjSQrxXdeAqKRuXW8EXXl
ul1hdLBRz1+mmkyZwKOWd0t1XOsO2f48fL8smqrGyGFogJGx2SoG23RFZUH/y5NA
wsmzc17rAE368s/NoAQg/VxrQ1S6zSQOYuBMlTPtSm1uL04sryDtr8JZjbXxB9KJ
4BtOgv3xcGKmQ1fdX0G7XmJRVT8in5PePq9O7wDf2laP1AMZI5lFNHphXjAhrwHb
X98cQLgPyCeKkwHRv9Ye7y3fLMGYDPm3Exkjl5C5h0RooJmCQGkyTZn4JM92FJBj
lufpUJmEd8rPjfSg33lgfWqj6QWeEVw4dfRAILXfUUlWt8BZDOE1ldXUBWdTL9mc
uqHsnu8xtbm/RIpqMLFS5TrjsgfmfHUaaTYSvP/UG9ZKi6VMuHgGu2WDfR0+jTzA
xzmxVtFwEZDjLmpug4tiW3q/zI9P3XCoyo5uPlks/Hupu9lMJok+kqLFcWlBjMF3
BOJwNLyzmUJ07yQ7H38k5JPQPpjuEBoJImbdC733p+caJyaeYTMwa312Hc1DRLKs
9K62MbG17oHQtyHZs9N5dFu+luEVwFuAJ3eUH8XhhkS8pUR0mzhsMXeEPqy9oUw5
banzCDs5aS8SOXXgEtqqcqiOrEAsLKeEPvMbNWg+FNMEcjh6C9Un7yQGNwSsb9SV
84Wmgw++rCGCFwCNWz969t6s5Fj/nH0+ynOyadEZKcObgAH7ba0fV24pk1dmKmHi
1azliVV/gWtQZW8rw+Ed7lJZv9Pjrb11zUmHc0Zwd0THoA418lV57kimmVf7KM1K
B3cjiRNb4SHcsFynJgOCu3ATsLpWRaa4MFD2Lq8jTo8ydcBNXKYiC0wW22pRwI9Q
DIf/RigMV6191ZSQmYhzFJRcCdHQhUy7isRwqh4psoto/DgpkY3f4WPUiTICJXif
kYDjU6LcyGnchKs2fTnHQTD8Cgq9X46yXG/3hpeyT335UJT8k+WNnql99PkhzehH
jrj2zf+nLYxJy3qsA4jUrovAlY5tkVLZrSoSU/7VM5XTTt66kF5PY+03XgCaSckT
EdQ4O8Z2npwTbvpg2ohNyNqRFjf+RFrtqNKElzl2RgDqpEmkB7lhVHp+obg1LofW
WkAZ14iraHacCvy5NQMjlgztvzI/Bp6GV6VMhOxC8EgLBwwobBrPviQ36zpX9Fbe
I6kE6N05bSUBgOEZ1iM3zK+cXa4O7UEe7Vv6AUgU4038Oq1FEaO0LUZMc98VaLrA
TBbom6C07Z+1GkJ+2KvgqBrpI4TeJ7ZZa25hV3Xris5YvHfU0t6ilJuYURhsMblI
amirT/B0DlCwInVMEGaKaLuP0aIKq4k53M5CQk5advYxe4pjR6W/yvcjDnCCkzHj
k7V4m7rcTiKc8AqMEWWuUQQETD6sZUJHRsn3G99z65O6xc63w/gg0pu8BvMUxD/Z
dwdAjsQrQzLmof+uD1nwCgldZKuFG+6NPazk+GOyyj4ezy3Susu66XSQgWGKCWQi
HdnhtpJ8XajbKJkIsUPYNe2r2Fj/9OtbeRshhsZ4/xj9/a0Ve2Dk8usGz9Rs0DQM
4sOayaZ/m0tzkAzQRRyi2dbrNcpguyEBMISOIgFWAwLjPkhNkCacUf/nvv25psQj
DZLYhQynDV09aK8LGlS3XzYftLtGVy1BGBC3apd9juPYKcRKu4KXcbNitaDftXWb
5OdB/AUSGDB2YUwGbsZR7YBFsff2qol1BPmKIfcJCgYa9BbUnezjIobkvhrH1Up3
c4/CQjegM2CHrWP4BOqc7UvaOoX/cK9gzko6lqeWcKEJComaOo7EI9zfSnaG/Ocb
cCyUPkQKsWaiEf5wTJ01kRT8ujPbgHb0vNZ29hxSm1d3W2dIehdLfQMydF0hAsz0
N/5dyZVETPOD5E8IJfqKrQuOJ23+uRGtGQoZcq8QOn7RyyOh+CYomk1uUoOc+yDj
AXEjDOhrt0igyKRq1mtV5cV9kPjeg/Qjc1OsEIEqSANu4ppeUL7z7fUgcAxcHbg8
Cpywc4XRv9NDKqJT2fCn31qB3aadXnqIIq2Agw983BWuoAvtZ1mMmvgWRgVi45Z6
W5D5xpKFfQ6gqAYh+bU21n+P01z8I80aNsQ7OO1mRZZkXSqYXSaBQNSs9uyOKk+X
v++s2sspRGRxg0ON34f344Yxanwd0iiZsUbEm7APhl8DTwuPqA/CazO2vqOwMgBl
KF+zmalOpXLi3bg1GZihzQgXapmd38tBahM7VmSDexH5lQRKTYtrfEgBR+wNzKZL
RNOdXVIHeFJUiVCnSK565b2/jaO6z/tbgkZI6VPlVXZHUjwj2NT2nQSlSTb9BPLE
/SLc4/zzA7/UxrgaY9tcuPH/6CjN/Lzoo7vS651mJvF8qD6QF+R6rich5PrrRZpk
2gAaDMSf+4QGQHRSp3AbQU88o9hBRp/t8Acckj9K5235G06HX9igY7GiVEJhVjoH
gVXfORMPBrqA4PiSLqTQOuqxUermT/lm2KTDX62hi0vgYvqFMsrK7FtmELGNAoe6
h31Wxqlr87NIPSeL7rW3PwcvkglfP3v/gBEEiUzGnsr70xN9jj1sS1+48BcwArVD
LJTqW6peiWSTJbdly97O9/dfLunpNERAFOWBnsNEvM77N4Y0eWo8tbtq3G+lgRBD
3qVhHQ0vg+SmfrH9sqx7jPOMfhbN0BrSKGoMFGFXcG/c5nwPHxb5fvnG77QpE/FU
LrnOYCm4HC7p85mV/ZTD0XI/pFcGVCbVyzdntf3fHIt1QXnqBhPg4WTbA0nQoore
VEs2pxZdxvtcEqnSg/vB3bISYsxwz/dJU43v+AU1h36HL3JtrImvymkiyA0BnEKY
BeFv9J8EBKY6uCidRrgORaREzHDkkWXZv/GQlQRcTWTyqOF3LneJEg8cXVXR3z8S
9Quqv+7mDbQCvxfE+TvCIBpBnUqbwKZ8fdF4h7iYTr7emBY4LCiX4hvnglFOMtN9
EreYmd+mYEfV306Ecmhaj6cKFdMQ+d78tIgC/ahRZGdWdG99Mqri+2mVgKjZxQzb
luPhfPpvxD2bguGXIQG377KW/5cPYIY+K2nGZtt1zFMWmfaorAzMVjEH2U0SEcVR
q2RBjZRXa9DalCyHrYkadvhT1EUlRDIWXipHnwQ0bly6AC1THh8sFpycdjWB7x8o
vDBbSlI9ikayG8tLFSRTJF6Z0BMKRYX8Yro+YuYrRmRfGa6atCW1It3FdL2WJmrR
cZSkgF0zfS0uzY0kcSXxr8/GqVNjwocTuiMCUIAlXAok06ss/1iXquHJIe9ckH1N
iGeQIhQl49Slqrf/0t0lYYTssAgQjGHWwTZiTJRzgHGic8c1hLASud6A0ab2LeOV
1HWKQhhLNBLDvsLPf1AeAGN2kO0Hvfjq3FPmWcwkUln72MO2+g4GQg17a/ltI2hv
/nLWJJ5ZaDoqIxS5e5Npy4Td74xHp3uxih5TlYCy6kuduNFYnlILd2cPCAsvLIpD
9dNv/yKL5Mkcjq7FCEy2zI9z6V4BGnYJpBm7/LShQUOVsQkZxuksyBW+5XsR+jXC
4WUFyE0mWrCXyLiZXj1BEsgx0FUFRD4CmTGDSLOCVE0SygU5jjrXetKxIvYuWSGJ
s7m58LJarXcD7zEobXURAaaK38pcmm7IasOKScQwfXPn0yOASTxE83qbGDagojqL
OTcaw0lyqVn2I+ukoS7ZWzzz5LbBs/0yDOvl1jKWSn8Ih/ggezej8sgNDDrFyrlg
oqdz3ug5T3dQoHesy6x//6IpFKUznMt3LKLdzG4vUp+i7lwPOBUBQzea2Erfyhck
UEoHiW3A9uVxwlKkU6osLJwDbWRfHuFW4T9Nkl0VoJYLnT8fImn+wgK8auOPRBta
bKradP72NlFI1UwG58UnqjXR8tO9c/svOSJCkTPbki5mTEzaFFjTrT2vdfu/ieA0
/e4dcMS3qf1/d4+OX8n2u7PEbUkVZUfgu1pHLhdHtY9xuueIbl33gpzwG3DZyoZu
K9+rYJ8DWu2W1TqFBjxjvp2JeRxiqJm6fH+YQugZwsoauKRIHqoY3SnOVd3bjsz8
6RM8izahP7qL0vQPIapIfqaXXxfmc/o6qIo4yGg4fZ8Uk/n75E2SwpVZSYwp21Zx
F7zhYKGd7Y6Fkesp8PdPXpST6U/RSLfh3ZhB5eIv/Y6HNZ2H7s/zHjkwM13c7GII
bs6p+mPZSz2aLqwSeCO0wTgvJ8Wl+fzuzrAV3PWlP2JjTqN7xMrtpXWikBWPoLcA
KkVlVflJPCS5AJoViu/MvQIHv2cmgnz9M+B4nl7iw4IOAhGewYTKqggfeb7SU7AO
bgtP6GPABVQN9Kzk224g+W5fCqgDGZ8q+ItPkGOYNnbk5fQY4zD3m1djOeq0zfAO
sa048d3naqOMuLtqTXk/VjkzDGBJkJJRswB2F42YT0obKiZuZ2FxJdROvjd3V/QG
AN6X1+HVGjyKDk85hPR7T+UibYeLyjKQiTbUGSDxkSlVzJo6Lg++Q7q6EsEGTomV
YRZ/G7T3HFs/TRynPo2VNgViTUzZY39pABqj8KXdU/ZUYAwAZk3iAyGD80DhDxSV
AhySdl1DeDZVzYGHOfvlkucnVOU6cyO1Y1no8bLimElPGrMNUh4N0eEZXjX3YogS
bYPB1mEhf205JuRm82PkA7MndLFAXXT49+/xaFFCGW8cqcwYNuXA4T5hS/FO5VAC
iCF4cuRQqMieD7n55InQ0b7tXWl2PExmi3yGxDaRaD2vrz4jiqb3/CF5x8C9+PqU
1ZyhmKrUD8Mk4VPhIXU3nHjMnKy/P6L0lvYGYnrv/cNL6BswRsuDf5y/Pg4KHR89
3e5AqwFoCGyPFGsWoVQk04HP3n9LlY8VLa74PRnh46XAAbcV77zuM6eoM+3DX5bE
p/ZaNELj4j3ocvHtuA7HzupuxCh5i6j/dB2SR7wR8yYjYxxRJ7Qr/B5N0qqWUBQa
cm+f56K7OD5tYXlXrksQsPJys1B9Xf/pU6IAAN8HVDzH244ZJen2y5Xtbi9tJnBv
vjVV4Cz9icDYVK03EyJMIvosl8lDEuNgoF3EMA5oAYAMpq0X6apf0p8f1AwO2Gf6
E6Ck0d+dg6NY4J+5774AsJWzTldFA+/DkhHXhBDi3N6My+IsBQBw003uzqbG5xWw
eTGcBPl8Ywo9cVbe0l7oAp0tM2kLEJojUs4HTVEyLcc8noptQ8FqQtUglozacXAr
sR3W6S/vDnlq0/ep1Puup8WveRKiUyUHDRPycABpgm4+XVQ5NYFXkPhU9WMoCaZt
SWnfM+6BXTfwce5lh01/6QC5LG8qar5HSbuEzpG3yEWrEhmHLFKvHUk2oUvJDxdV
p4JjBPSdFI7dlLzH0sgqzxfsDvxaSIw09+S/N1IxzXhRbrSXNsmF+x3cNRgo6o1d
075sBmMKkn829IBd+e7G2Ld8H/jVuWRwW6mlfzIJrAUlvRN8XIvLoHOQjEOmLNtS
k2kfnoEBG8UoL54lP3kk12H/LNWfBzUGVeJ6ijvrqV1bvy8w35+q5CXrM1E2QNUC
TPahclpZmACJQKjDhy93qCTuBUYEJgCkE8Jtty/WDcdQ+VLqcUJzpPtnet7g8iZx
mbwEu7211u8ghAVeErpbmmaA65Jn6dlZ+AxEGkAjHkwLU3fxRzBtfFoBjL0K/PcK
QMk2/raCa/Wb/y9WbP3dW9hUcbKuYdHHmYy15bg2vt81trsZoVtDeDpG/xJCOrXc
ZOkPsjHltPL4hDI/VoqNk3X4hZ7YifP3dpyKAU4vr1XL/ROfqWs+r2z0Mw9az1Nh
m0dSpeWB7Igr0/+5OHPq4LaS8k6czNKZayQ/zkyAS3oudyHDPjVQcsZcaDF5H3DE
UaexCBBwWJU/GgKHRiCDaitXpGZgA+aDjmADFBRTUixbZHyir2Y/KTw2W5q2BY0U
F2NRaHZ9simHxZ0DKWUspW2M87PTTBlsRDxiYd3ssN1XVStkGwztQJUfTdvVMxAi
z/bJRSpReiMQJO44A2EFQIbv316LzhSPszWPtOXjlNmuClfB+/L0TmdhxL6FQ4rs
XJ1k47VIdH0/yhaJbYgabhWUmMTkVVb5dgGsk7eOVpkfk1r3RUqE/IrvhpApdUtp
8hGNCzQC8DlZSOF/ulvC7sJayY8D/y2L8hHsrDz7dqAokdCYcEh5CaUDFj7vO7o4
cP/UeXHjb9PsHs/VseRqTz+ncPXhn0Dc1ULBwSyXRwZO8NEY3tczGGZhRAYBHRnS
w2P5x/Ww6nbnG4WC02yL9h3PODjlf6ov8QACj6H82i+AvYMgId2Y6q3kvgns7jS6
2S/a3TrlFvQiLrZIZj/en3ZJ/FScpDHEjk4SiX+Gny1AqL698hPM3YqfSj5GCdFZ
e9p/uyB8TxeFm+VLVSEL5jXzs97Bii2G90HD19IZljD9Vp6KngYyVyUr/a4l/eo3
OwkOQnwUnCrUB3B4OaxyhQ+1RsxadZQfncrogjuZzrqM3DWH9ak1g2mSW9QHjXVy
ey5rbasZnlcfqfO6JwKOzHB3/lzwZSulacoF2ZUdO02mS/6Gv2VxnSENSjF3udtz
a+dD2Gf9oMU5Nr65aexUXFlXD0WUJAkLv2efIEz+oeBJgoKttO1s3NG/Q64MjC00
DG2qlmNuGfvFxSjlzns7MJZtTfi2I7grUgxwdGiT3oujct8l2gw/TsdkJTHqqY8G
uXbfQZBt0EcPa7xMolFocZcGGPnb9S6zKhcrGfLWAoAJbqIJ8xAC2jI1NTUKj9fw
nWpFJaC+L1rs86nWxOd5lDgW/MZnej0lGBEsBEXwW4/NeUXHJ4FvIP/n8koPiAfr
X4p/kwZCDtCJMFs1bHj0kpwvzwINpp5Chtcf8Nz6WP7FE5RrVqmzZCuqgMFeQauq
wRyIr8RlXFCwRh352W/VVga9+V4AO5qfql6Q5iPGgPFRjbX22W7wUNpP2fJUZ4sF
COpJTekTSumSYGuw8PDiurhQqrYocbfDYkoQ0ET0RI20N+udrU9dy1rXK1KQFwg9
Seua1pjzdxkIyMH20NoIJULk1cY8zXzc3YhVsLIUdG97ugX+g1RXPbJ+i67v1LTS
kzKFVkMmnABt9ZUNaJ5rGG/SIsaxyAGI1TEYDtx6tL6MwDcpmKvu8ctSXTuKh+Uk
BwXf5Pp9ibtpsvsxx1o04Wf81xFV8a8KBXbwuJwiE3huHUrrKu4CiILKl37nmTjC
bL4M8bG/kjJhobM4XS+KMcPt3AjPI1yXdD505hRquM00NuyCPVEGchWxuIJ1CbkV
Lefeg8Cg8sPwj4k8nPJrAr2jBKBt+2aQz0Q4x3O+FyZL75CD3wKG0JC7A4AxTwhr
OWm8atiNlZb70HbgOjP7uLjwBQIb1rQgBPM0UC7SM/5m9QKCabhAxBQeXb7iLAAb
wapI9HP5FfAz5fcKsOtyIF4z+30ZObMvkHQRmgYyVHtPAPNWLxyfiQAmaCDMJofs
jGO4S18QGiNgPcFJ/iiacXk6xz+lMGh2ix7MRjF/Cz735IAh1e8K3up171ClwV+J
Woc6H3bXki+KZqai0kt0Cwzy6d2k1C5beIt2cGrM7w4dD7GoS39GSrXYzSneJTTr
i48eRfPgwDTsVj3XkiRlLNbJ6BYSzLWfPn3L5+cGSCa1Gcw9LT2YkDL3N8JFOzjG
/5eo8e5M7+sC6OIllRD8tijl7d/SrFWP5jq1vUvfrJZROdQ+rnw/eHy1clMIXKBf
YQwh+8qdo0hwojDz1kzOP8AhyUmmSyZKFl6WKAKGj0zz/2HV3QkBcuHcyQs4HLt+
Vcz13jxdn/tmRYgqlCIPLjB30OGoY6x5iz99Y9cyxElhlewF2VZCdLc+k2wA+9Kj
y5KTFrB31xAwR6hgAUihJRkMgOY3/Rx3MmyleaqoUp2kW8FV8L4v+3HvvA9i+1Se
DwW0bPsFq7j9Hid8nKQTu3pWoK+qpkNzViPS+7i0MZU3pgU14ZOIzrF4u1vppCbB
dNUu7z6g4Fq6njb/JFES6X3bGbZYtk3H+eSfVqMFDOIkXnXahpJpF134J3afbBW2
8Lt8BrVk7emYmWGoItLJX8VtEGFVmXffrBuVr4xiRO4jEfnm7bxevz3NoIdtf64u
3VeTNPt8drmB2OhNSd3ekpc3jR366cfbzatr4wTTm4cGI/gNZ1LRheq2gDH+dmZE
TiLgeq4VT5GIwliybvjC0DwE7iGNN5oWgw+niF/3kd9WfbMTTQyJYiIyGeTFLNMo
aN6a7cmDDdFxCUoH5Gcq3jPF/YhY2FRK5q4TPOVlDlIIuZd/RLpw6loZ4mVRV9pP
iSU6TND3SLVKcpTNQ+4XDYqdmnDIUwvvCZY4jkBErceMFct3i0wNZWl836vaC45O
r6gF8kZ3cHcFA+iwh06Bf7+6oGLEKnLawfJQqUxjk4Y6lyzsfuqdfiiqU4O4mVIc
4VVXXr7ONwna1Qf3oYSeWC5z1zCxyO0cylO5RlKWuPva7+n2CtdS9suZ2YlPAsn+
IPHKyjA/9I0C1hLD3whBbSTuNWcl7/EZhxdSs8GyNmCWynGC+41vUCinGfqO08Z7
Fv9Gh9wOGW51LVYMo0A9SbTBiBVei+1ze+bjAWeMHqduMh9dklT9ggp/q3hgYtut
45/w9YPmvb70IyyUn+FLQA+CcBLzLI4FMcaHcNheGEJqKOWQR8UpNsLnft+LScX0
NxTpG3wAe0yCGqz7cL9egLPaWGxM9r0px2whn1v9GInAVJvUAdogNmYyEkxaxMXF
sWTAyddRwTqcfX1+VwSPGPtoQiauIBLz39gqepeVJP8rx0gKD/G24lTkviDiLx19
qTXBuvt8AWwvJbtMEoNlHR/TEl+Gj3e98KoGb1JzvygEQcYVGfwzXAlnsdwxaTG2
we8YKpUTigS4NLNwtxtKERWm8g+R1ZBP/ovjBahfsgupqPvXLUprklPRw0OCxCM7
6vM87UZTni37pFjersVksnOum0MEfMLYtJv19mDQc3U+sqHTPq6JKP7ahAYrlALw
KcGsorenZ50MYKRJbr1OogVH/o3PhLA5fEiGSQZlYMLPX4Yr6QxD7OVMwSd4cEZb
GJadv+nK/YAXaWXVD3HTYH4KmHuxptVamh30h3cgrheVuSIU1HUtTMCOk343WAq2
agqv/2/UykQcrwNefCyfhkWuI7jk/MsOn5wLXOIvhwjVj/jO2FCbs1KAFyUkvKJi
Nb+0MBC2PdxG4AuVQuX3evtG6V8duVXiuFUtfYSYAOWZp0EpAftLjnZ5aj7X8jqx
wuokGFnNFm5fFVyh05L3Op7C+W8PmeL9lWMKVGeBYh+USs7kCsGOxJu4IAagkYpP
WDtN8oIekiZF72mg8BYIz+MxCIOLX3HdMF0kHiaU1arpunfTmS7/gGukW3TfBJXX
1OrJrvjDAI0GzQbKeq4yL8KKCB18V351JGVd857DxDJ/BB5w4KRf/3GqnFQovxu9
lxFoYVRDDflifShGz+TI85v36GRpjGqOjQRY+v1JibPEu8s7GPoex/CizN6BBIQP
XpaCtOBu/mHHKxEtWgv+gsfijBYHVEjM6QRvWnPdxXSEehA6ByAMMBwfqlY0mYYy
Z7VTho5sHd57aT1WpDd0IlqDuCoySU8jmlXNRUyp7A8N34f3ylSL81lxsTRyAJWM
rApZ/jtQTNJ2RrXur9OL2I8ijTHSEtsdHsNg/DauyNtN2DJp0dOjWdw6C3YKTu+h
pV6hswJ13pm9bmnw4FDnYb3C5EvzqZ4go15VJI2fWDb1PTQrxhui4MsfwHa2v7af
aaQKYj79bpsQWC+MRTx9sTih4NPgqtzwGsmWNFXBNbcwpkCibxeHdVCZLtCHR3mZ
YBGUdxIho2JkKxEY8w+oy+gUH3mmt4mHPdUd35U6WUzMyqqTUKOLwMD3c5kY/KiV
jklBmnPU0NQW0xomQ5yFH6ES2GA0lX9dsvqukL9nGc/1Tf3lcz8xOh7kymnMAw7Y
vWZpC9tj70jfFIn42jY6OHJrCpeP0GeIYnMhiyH3k6riocCCFWNAkvV9q+uM7JaH
IKKV5W+Bu9qOKan4MUpfq6F8SsYUajURFfLkZjBzbKuiJHoKJr+0HHK67ybQdY+L
hTEcWmvX4Bp23n7oD3XJS5r1p1a+5c4FKIBYbPIZLtipIR+ENY+C3iU5RQneEfba
M9ZMbgnS6KQisREeX6ac5CHPvqR8KHz1HAyJIZb+Uiyb71oLAryCnyYyvHtETf0+
pt7p7ldAvtslGu+o+AuLZvxCa/6XiJh8razoQZxAxBl/uQmtSGjtlVWH1LorxA+p
6LcDgCIGiMNdmA3oqQkITUy8mpfFkhAUpGwtHrhm/mqhHWkOtdMcwur5dhOrW6a/
ejTRCHwQuWRmY3HHLN4w3RvEduICSRc/cZQ4We+i527LlNN7N5N0fgDHmemU1vqT
rRB/iqdgdd2R53IrRIuMT0Jl/0V6Lf8OOcQFenAi89gwOrN57CnBza9w8PLnGnPb
BdpDH2VVrqyYTTtbvp3r6/ocYgLwfaCvHlYXTEO3WyrLO1zkAJdN4uobI+MVVC+x
nvV1KxgAh+hdspO/wluz+tQb2JN74gmEN9jN+zk7qfjce1afKfgqYvHGpDRJ3m0d
o/gaBJfI8jXjmjuEMpwAJ8V7vImzFHaeociQsDXhgQLnHfQkCzF3Y1SXXDf/RWwP
WwE7Du91VwIR16wVJ2V2XUnwkLMqdV7LkkVlLvjHEQPGx/yERjiLW0fbh1bdGWCu
QOlHiVhIkg3vLHV+D8LWgSAGJonzxUUzQM0eqJNTWJml6yyS3w02Ipc1nsx6HOUW
gnq2SsUZKS20pi/RmCEhmxKGROdQGpbe7vT+ORsrWSL5gBU54Ie1XJTtcEI4gjMK
bUeEr3+eLZvlNCsbbrRNmhehnoF0kWspnIwwKaj5rDxPv05cvC8MRKamXv4+zoM7
Hfxz7A114mPVDDryatYp0w4u7NM82D/IAt889dSQzB2m1vLJgwRAMsTQ3N8jyFbQ
/l6H54aerJloYGwC/AjI1uV/ozUwYaPYG1VqSL72c+pQULNMqFAiNux84Bn2Xi20
lFplWiFVhWpwDCvQhcO/G1JpqyjopvqCaSKjiKga95vnRgz18WJ8zR8eIBPXU5jz
TkhwYClBWG9p4FxLgBgb0rtSjL95FhYyJbbQTj5mm3ld/Bi7zIM5fRYRAX5fMLHU
1TamMm+lZyATpfC70/IEwvGHXQt9k+WraUTzt+62c6I7IrdG+27sNdCNdVqHl0MS
FHKKZVDCtpMnk/eKexxw2Q0B3e4HHs7ESAQxJmsvcHuV4Yx0klCmoZm5fF/1ACt6
a1yfPfMcMo9hW/t1wLspIMEYQS+OH/c1ro0PPocTX8SfHrTd0K2HCLK/QbdUgpeO
6uCyT3QEp8hr0w3GCGKqdy1M0htHqVSE5buENi0FKKReIb6aVqYZbp6j5w0mOo0p
akNe4xMjt9gLnI+NAvvcfG75Jj6Nqp67L8ndqVHj/6lA5MHmN/AGieGn7e06KYTX
8ziE8his/8D7kIuNB9MrI8uWcnUG1X43aYkUPtmKt45vOhWInvBwRD+8cYQUi/HI
CzH0SAesIt+5nKwwO9HqQzLDTLGIFaBDUw4pTHB+RT93ju2v7J+2AtsFv89wMOCw
y+cbEvftUichZ8xPVp5NCjLP/Qcp53qmurOEoZKr1RIMahKRjlbEIJuVQCgXkX4Y
1VKOadQli9Z/OYQXKmj1BOHJOzA1NAtOECxrNy7wfpUaF7T1k+u2hw0EQxC1hCSQ
AuX/cgDbYSiFd4qZHf+3NZgjG8HIgh+05ByU1zIZ8gCrbzwJsD5xOT3fFTQ83pDH
LhINgSOMV1vJ7m+pT2LU8Ll2GqupKC+OG0upB5jhOOpEuYLhm7RY9vhH3lvJ4i12
ik+CDcELonhezt80M6BjVBf3PW3DHFeC0T+U5NLgWsJBSqP3C0yUibhr45Lcj7z7
aubWdMMA73nc//EfJ0Tb6gnKOX2VLov4Y5n1XJMtWOyN4vh1sg87mKcc83eetn9k
XNfi82ivQmobnCb8JO1c7UPmmXHWkq+WopdkQ2+mJjCiecK1nwTsEQuPd6VAUAoY
olZDCvvtF36AA5dtxKf/Q+xya4d6cuFoM3XYDVDTBgV3t4D11DL5E2q2MIotP5VV
yke4Gm3843K+9zw5Q2VC6ZOWQxr5hHONFZr9v+lgf7e2roBLVxbJBt+ttJNzn4Ev
7/Z/WPj2qTrMU6WrDYF3WsQwAdqtgEh0mhgxMke0Xtd2wxssQGKPMCvsZImbGV/L
d6Iaxb6YOGAcKtQgTIommPODu4l99BZHzVfNqZ6NMYPC0mTo1RHP54k1l+fAtXeh
u/GtzveYc/pGvhEcUiJQ5JL/o9lKRHHou18SMYHzL9EenUUhFEDefHQEEZALFd9i
2HS3kKE+hbSwH7wkP8POdt8+zYrabYwEvo00BxbIiJmR6mjjTDwUemSpb3ddp9TB
aOpBL36cFiFtqWdVYvaRGbjEzS+Ngeekrj+9AfzXCAAo5bIiOeCIbr2ci1iPlk2L
8Mx8Ej1Y3LJCZLAr88akFj9SFH+p9mX5vHX/SfAqM4b/hyvMNc1Z6LCxwSbEDc/h
6djFY7pBp/EkEoCbxso3TDFTjoHWhh0cNJdx8ayDPsi9SISCTcgDE/FKU5EPszoy
3oi/XR2TfDuW4O+BeOHJsIYSg+jazQYekvom9K+VLAc9ua/unrf4OZLNaCMRWd0b
iT+AovuBnwZlHF9Hu54ctfcsofZU1tYm7+n7z0EpdH3cIG+SnqR83FW0vxAbFYc4
inA/lxkPPFdklpP5RY4uXk/2CPIvDKohfUzTAqfiWBzeGqIFlK0ztiqqyVV7Epns
U4CqGcrSlzTTPAoT04BJ0JPoD1t5lVsw1cyfKuz7OsAOiwAGAoc0BwL1b8OzSUbg
b2L4ejmkJZ8auxln5wImeRotQ0MdpsBXDVHwShmyOa0ckcR+tzIhda+xOZgCTvNh
sD7bzjpExFSBzCA/HBHKIHn/UHwChdOZoNqYIwB0lFuiRlstzBcJUGY9AFOEaV+S
CKkKzI+wSiTG+yYbPCo88Th5K3E6SwCCXc+4SxN3tINAyP0opi23D4q2ph+I2rnF
3CRkUrTcChP0SsAwua/PiAN5WbnuHLvTrYF61Kl9gYf3KmGBYk9LsSs+EGIg11of
Iu/HVPlRpFN9UoI0ytnrmu21eHxz/2ueMgN29NU12QZhE3jgsc9FofrSysB0UqUM
CwqqKI49xca67tMupWVBlGnbq6T3sQLNS+5PEOIgm7fEJw777oRbHNoiGYdadLgO
2WepILvk4UteGpP0AWpJ+cGiYByxUEZ81h3M6g5j55Z0LrZhuFjysZsH5bdxiW+c
XWarJtj1mk4jzuMTmf+S2L4/akZCH2B+D4cfH86QPYk72VqyvNG6XMna10xWOTrJ
WOSAsjgkaiqzE2Qb7ELOLRoQ7AZX138+/fTCElnk6OIqVOs0Ji8/RNtzAtg3nEn3
/wWKmdvw2+JrOT02FIApgy7DxfhS5pT7g9/yZUl9mj232alO7F/nOeg/pWFBrs+J
H2BtAk9Ipte9o6ZXHUUq5VtPEGlg9P0h+bY/PqaM16xeyIrfyE2vTw4BC8+VekUo
Ukv6kKZ9Bye4tYGiRK4krsdmSCT9XF4YYmGbBlEDxY4AlU9i9VUeNF31DwEXm5Sl
rqZfIGTn4S+6kjkqwDSw8ixxnURAsJphSQUwpB5y2ZPpPE2dGRrUZl+DJM6CgIp8
6jYrm03X9nrUknipuE00iIEMCiHy4YrH2l7G346dRYGmfdHwpZ29LHBCrje7IJ/W
j9BA7AOwgbwt+ctJjZbRVFa7aHAJARvMhnDFVNH6P/Y1FKZmJu8GPlMl+KgDgrTL
Qqg6L1jx8+HssH6AEPVIrCRyc5l6foSj2cy+F94rPN9ZS1GK+FvEv49hK08otYMC
CDQOWOBFA+LC5BPYtMlOIcOjxyrjjfBRYPJncw1zC59E5EbrEvh2FEu7wg+vBqS9
/hLps6lQ+1iFZWEPYSp4//Njn+gwE8l9li2/j7IT0AlxskAeFoLpmwTRjIMJkiMT
OHIF92ZdqMuQvNY30HcBR/r2OnBAnMfTQkj+QLRiCgV9h6918KJ5d0LOEOGCrVsZ
dJNlWdkWEY0NGJcfDhaPi0MpK5C0cUC3cPV0K2NbTHUYfQNZaFTBHCcDlm0hA5EO
D8qhrIzUwhlcBCoFs2mR5kxjhNTsyziJLhTxdlfDv82amJEvuKu53TECagne4GND
JhdtD4Nz9Pa+puAMYSAQfCGErYbDagg4Mxcsen116B6t5LbFLmpwGXXb+vShg+p9
s8bsIB9PgyyWOLBWcb+XPPrp0POy9FfY9sM5Hywk84cHOzGkuK8Tr4CsyKRX30xN
lxwpSqS9ieuhDg1fsaXtgHSQ7WnVr+5FJoW+D2ntGBd77ICxjqiiOLAecEOJF02W
YtDAny1ZaeVkvjDA+s8U2vVsAiZb5FuhCKXTerfpxa10ZAYEHkiuToucRU6+YXlZ
GqerFmKB3G74GU1Kxad8KFzfM/nLs/27sFArVLmbnmIEIFOr2nO5TScyxkka/50q
hU9mupp2YTdqr0+XghNoitgJiEnRJXvBaTLhEPMEoYY0yPCGjToklWVt8e2ss7/6
M7D7UzEJSW7QyfDYke6wH15iF2wdQ1EgX8DzXezr0zVvPiXvtUNYrqkWY+nM262p
F7wyGCWut8RLmfy7yIkbEEn3l3TXp/WU4qY6qh3mUKfwScOib4ZWsksH4vAUbn5i
T51FfhSyGlj0SQyYOKDTMqbQKXQ/t/8wyLEL2ylGBDzyonqAwE/i2fLxTMP3R7ca
K3MlpDFSv10KTE2QtykMmTCFQBlmMrs0MAruPqdV32Z+x5acJ4reML528aVPhvkO
g2okBpZpswfTPqJVfe0fl5seT/mNGbdmHKcimWV7LOoj+i1jMLVZfUhEGeKJJUWY
rnlIPPHgzuIqE4PoLSXw3gbIpmhhoqhRDyfadK/Z4to0b7XNdm06Eq0Qs/ea1CwV
Gxb5LGcuziqR/K72TTqSNRWVLsWC+nUD8yF7LLsNB2t3tY0f5ls+KJinErHJ9Bq+
KG1Op7vGOOXxF7DOe4XlO92UnPbR8sQj5fFZar53ZDehjs7FMAe3UIu6+7w4M+JA
Fac++YvAfsOj/RNH6PvOpRBaDBOrKUwtslFcULQykb2ndGiz9DxhLt7wula4TWa+
Fs4YIxWIpyuZ2nzaosHnVFr3Vfv0MO2c4YUc2uduCt1n0Okm37DMEnHHWcaYb8Tf
e5KWSvzQGDQtR2ODb7BpwEh1RjcjRA+Q5oPqhOpKcNTMz0aWKGMY1/5VqjeWyhF5
QkYyYc6hTWTSdZM7GgoaSg/TX5tiuL3iAHZySxZBtcej8UfjBoKCjH8R1OyStujb
ib9JNKRPSJvAh6ZBuXzd35oPanSZMfshF6rT0gYKSaxWw9Y0kAnORAXxbuxISi6F
2GIXFH94UG+jvboBNy0NKvgwKU2t/8E/p+XbOPcTd6yPWnPiaPgEWMwNP5rCDBAO
UzCVrxiU95ZpBtnbP1xSIuvBNMCOujIE078ZUwkW4zr9NMs5skmpfSqfdzoxGTDZ
ISIV+CnNaZtDLFWFqzV79/xCqWagoMka0q+nE7zC4xPYsogLwcXi9gNa5vN2GGEt
vc4jm/RT7HKtb7FpC04BdgKVUf1R2lP/TzcSc2IzYiGdpojX7U1s9Jeya8BOsBw9
LMjJH2Gln/T0F0ujva1pI8vRAgMroPQ9ot43ytlgzqXVxHzJda3KMba4a/kVlQdb
Nx/swlxdOIb21u48fIfGoGhp4QHNowXY+LZEnKu+/5x1+oCZEzmuWho6qJCDQfOF
dtCic6dvsFkHyOpv4W9lXGq0ZxfXPKMRk5iDTWpo7qWeNgoxx8RuwOyvvoysXJ1c
U+KVHCD76ry06pUY+/8zqIlkVC8az2VHNX3ATpnWK6qc8HXuPxFcLKdJ+IHiePBm
uLu/0yTchkNiiPHND1ARcoab2JK5Qhq9kiofPXkdW3NbcfPLtYeWgWmdoMriQ98+
p4VK6p+jvXXMB7FA4rRoja5klWsP/spw6QV3ioyatQEoQqjUhmtlt3wDpAtrhYSQ
Sl8cPrFotTQC5DJ/5BF7aY2ULvvd9VwXwD3CNmqPc+74CuR99UzXbCfqdOy0bXV+
Y22l/Eqx/IVomgWIX03hCF/mmc2VOBHcjyAF5ygoPNIexlrqcUp1oaGzxNVV9L/w
KR3eocA2f/hY5/Fn3QmtQxvOzDi/oWDSFwKblyrSGxCJgIaysEocC6krZ0wTBQdW
X4jyCRgu+qj9aPTlbwWyI0dVNlF+hbSD6LBgJvDI9a3CDgs4g16GjfIo9+1r7gOo
q6Kf1HT0DPAOvw86go79rSOOyXxtK9q95Rq9H9dcbaPcBB++zj6uYWqAoyEnQffc
lhfjmlsekSmXuSlebjFff00K8Mo9RHtVWHpalCzro40RuIjkC+LFWz2LM1okFcr/
TC4dbzU7stMF+xDOABSFrlH5M0lvx41a1fEJKEk/A8ng3c8KKy2XbimscNqsemXz
fRlbUcnMhj+j2JALzf0ohpJZgIru+8mkpDv5cMo7WPMWTHKfmU+oE/yQa8CW7EOq
isHhWmRNYxVEaOSxpUpJiwzYZuO/gRrL9lfRDv+LPlwCTNPHuIcz6lRtqYCds8Sc
FdajlFk8ceLrAbppOwIriaf/5+r721ZWgQ2Z61dPOkwU2PQqUpqijIFoeWTaHKMK
JCM30K/AbnR4zB1SxOSwyQTogYMGvczdZBiKIP4+p+vXiYMCEoZA+2Zk4Dic1d4x
vN/E1yQgf1jx0XSY05o5xTnMBzBkvD9nyB++NtVglZRna26icZ6FrGe71VSg4qej
FHQF3e4MercZantB3pSWVRjvqlKHJ4JhReFt9sh2X7kCcI0TEGEYD2fAFr+zK4Vl
KkJ1TjVCrcNEj/Esie9wEZ3Es2lf2PnJj2dySd168zDC+mvwIbRJVojcVGhz3pD4
TquSP5gl3VoUCV9GabYvEGaSlWcyTMHbbKTwZM75AinFe3h3vDCJZ3YgwK6M+9pF
ZOOQ1ToQm+YISzGAcVxJZUXEnSQ9hyuleUlPohHdC7+AVzZ7eV53U9ZF1ZFng+DX
dWm7Sk0Qu/7XIB5Iw792aQskVkaYd6RSWZKmerlp/dzc6Z4Ykahioxw2t0TovLKT
uATHBf5JjMU4kp1d/j8zLXsm1kwj/3oOkeNIninKRkIrAuc15DV1jH9GCKS731MN
6wie1wvOW8TEFpSHtWasgy6hrtk6xsXPJeU10DFWpwQmItnKpG8cxYfNDJqPuFlr
83OQ4CgtiSmXuDA0b/kpTTE0pIJCDB4p5TCXHRpWh8r1yiM5NdtOvxgmjnjihmZu
bNoA9BkHd+yanusKWxIeH6YBwuYvH+kxiWm94ZWf8qCGb+4pI1sAqvRgcx6hS/tP
iqbIN37Y9ffQwirRR/A59D5eR/MQmAraB05eRunuZMezj/Iy9HnrHUic3GTwroyN
oEBVTTpm8aegunsGUJvOurBwwyJ53GNknMRF8YOuuhxVzN+7Br9GeiDzcD33To2y
r7SoYBls+SVz4AHyxMk32gAr/ohfcKvuzbiuWVM+VkBHiqZ6nP/pKxTbNegnR++5
xOe58RaR/Ce4sztZe+2P7Shic/aHIVf2eyd2vCP9vnfw5/3kxmdvTXFlzFBTey/6
2Pm5qogIF2poq42j+1CZMbiqUjmV8sCunz6nNvcPMvTpwWFboZ05mq9TPAaHkBiB
r6S6vt0x2/nc7TzimJAdjiL39ZbJIUYQMb/Yj+SwnR7x18waPlpnoBdiE7O35a40
tNPpROMKlAyq1J6kvsyMkJJZVg/B9vY0f4jSYA7wNHAshGHaGKjl/IAldI3qmJB5
ioUkrdPPFGQrb/N8KcyiHuprXN204c1/HweOBpfjBqi8alxOAOW+nlMvvip5UbcO
vEXrpDwPqO4NYzkgKMN91ewYYzW9Q3kQRrSgNXPRSTzQ5iwVL6wvrewq9jYqbq3V
B9OIFosJlnlGFVr1mY2d4hsiAVV9Og7cW2zgKV9Fy6BIObaXkd2/mSy4Qqd9OHPR
kRhH5TyIV2gSM9kCFRIKjKdZ4THFunYG70vuMCPX43l5JpNQqMXAhYPhdKP5ZYzo
Lqu8GLRaKUgB4021ZL+P4LNfwftOVVomLalkRncF/px+6HYuZsC6L+cIZxUVjc9R
rLNrwPPJjfZJ7H5bZMC64PWntJDkMuYFWx3uXWPM7IqflOevRRLX8cwaDxe1cD94
WaiMw+nQEvoOBru/IjPHrpLY257CH+OSVPMOcA4d6ETDv/UIq58F8P/h0m5z5W4P
RbEhcKmB+l0ZFfyxJNuii+goxIJFN6a44hA59bEYUPO2pJSsETc1MIe7X+F+Q0OJ
U/zFQGQy40RSN5W4nbUc44NwjcQWBs5Aq9k0QjPZQ1VW0UvoYJxNhNQeAYkAPmPR
rR9E/iyAoWRUiXzitlpnflG0Mu6fJW7tfREAtE7bRpUX5DgteqK9hcUxpPFXqCGF
nkf9XlgLV4Lz3RjtU4wTUFr/RrlveBzB2muuAD6/Ygj500N+HmhJ0gsSw3VihIX4
zbMf2WAC4TnBwEd3C7b0XIeJbd9ApegtrtfAeLxa3T2s+dl3fX9Pn9jrQqdq4kMB
qfRjzfrC9KfHhCZt7lgU8n6DuB31gAYJA5BknS2yEv7fAxybMP9jHvaj0V5GXIkd
M1KAcUWfGX2TYavfeNhPB2JVbv7JWVRCuzZ7dTWMZkLDZZflefxSenGBMnoRgXP6
G/lW4cbh8aH0rNB8gQSr20pLDwpBENoufcc+C8aJ4JE5V0miTFr7PhkCATo/mWZr
kES0xb180tu7SJuYJ5uLM/F9g3jfiizGO8IRy5KEWU7MIyZjcHWK3paijwVgtqHU
25O5NSHHC621bCGEkglr62j/NCoNwJO9xVrDAouLWAP9SEGWbJAR95aTpJUfNw6p
r0jCpd1yWHGWG8eBSzb5hmRJz+bqvo/n/b5ZS6wXVdX6/11cB6Kl9x/neSNnIF4y
XO9hIJROTlsp4vCB7q58meMUvgdHl5tYLSlB4e+EKnZxwn3lJC6WvHvV1FBN9ZLu
gniraUkHjD+IgUQ2jDwGQ07t12qoB3WEeGFDdzmTt1STrCLZ0Xuhox5scViKEABR
cWbXcDR28AUqX0QXcgu6FNFW/iF5bFxELGronCPF9NfiamJdrkmobBib+4mVOzat
LZVvOGXHi25F5d9rpF5cEAj2XGusopQp09/rF/i434j4J8fM3JnmBrAlCO5AnrBd
bkd571YRqZpptU2y+NnojYLZnb+h8LMZ+0qrAi1i2GxUU3EnRp+VxQGKtWKm0bly
I50tE4DjhMyBIDd41revLT6KCXVl0WK+LRw3GK89h0SDOjTwbIz8zV9gGZ2GJYTd
7znOzkIqVzAufUqu09s9jWi+tkLUDawCv0PSOwZe7pTGgSKi8m1RMKRRR+PiLYZc
GOK1QwZHS5WqrpegH5P52udk3SE+RqQMK8dRlju54xf9Qd2GhtgNKbWmQ2a1ONPc
cmergG9nXnMK6wqG3KOMzuvKwW5ReFPTNEkDsV0JC9Kb2Mn8BJRQ438yVGV0lsFO
v8HlXXpMjWe2vkDPdk2HeLpT1nty6kWi4SF5IxktMYTpLqRMgbjyyM7PEf92HoSM
u7F8tEF4gnHaIa7IkwV0oOdaLyOOAm4CCzlhsrhqOHlvtbQ45V40ULpuzpodDQNi
JIUTLwflwIHLyCL0Vd4IKnjrVziUTABx0utt8z8Qb0YR9VBahqoLD8HzzFUIhq8l
Ii9R46DqsFLah6a4kuNcPLhzUorOfVoNk2NgHao2yNNSSUXJmmH3IuXdszcnEF8s
gblhWf+ydHyEbKa3MtRQU2zXZwVHzMe+XijbK76W3r2Pvf/fGtGuuClawhvg4wIy
Fh9QKzAwAhKVVeG48jLq9dye3ZgRnOtxwzoh+9jkzGRW2X7GczBWib9xvpfIpHvq
LDUGOlc9O9mxHF8J/ZiXkK67QzaGr7ZOB4qmRY180vmIY70FDco33R0HN4zHl6nO
72esGGvbXoAqYJa8lgN4XOza5hQ197B6m6fKWzJedmO7EIgyE5+pKlTdrScWoscg
zNPOiFvDawe57iv0AFxJNkMiOvjAxctx+7EFJWPwosZ1Y0770WSLUTYrYEGznLsv
p6sh6U13KKjt9yQmI8qXjFQeuR6asIb10mZAg9KtJOLjhVgEOlVaz5jDKcAYhKC1
WdUfVOexhrUh68xuOxb65Ib4BniSD9rW9pXWQJbo+vFSyw4PqelwFlewRYc2lo8+
uOD3aXRiAc1U5un5n9wZgJRG2BOWAjjIA/IlWEJ7JVmDJHin0f+Tu6eluMRqzRV+
7yAGAc2OGVe2ekOJ8iulgNvjAsVTdNU3CeywcmCcLjjiqc9D392N87Ul55U97lQw
YizdHZBhCM0Pfp6USsJX4jVGLO/07eu9r6iZxW7rK/iEciR4ntGLfD8W5SStnaZR
PwcJUzmS5JvXhMtWVDz0YXkYspRdWfu5Yg2Y82+DMvG5AtRx984mFLb2Y/VQ9oWW
B0kkNaowApr5x3vy1lHjJf3RzQAO/lb+KdVla4vl0eZW1hkczfevRaeJ5vvCSeZI
OhYdxVZspJR+CNdyqgk8r+QgGrv/nQJXj63paasHOxubyWi0Tji8Ade94M4t/78E
GCbabw6RPoLqgUX1cqIkj2pSZwuXBvNH91gPbqCFMsmN4cZie/XozabjbcMpY/Iq
D5uuao2p6izdTmxdOomKFVSC4ateuWpMiQc/1KhH0Ii3bQTnufnTTT93R4WD/ZVo
Oh4PUIrkoC5NQizwkYK+PU1VIR/R7o4sLmJEYlY0iXo/rgCZNj63eyeSSty17/JM
j7jyMv2lBAJhKNVzw4I9yezbjXj7rFBOUkjRioy3Oi/oi1/RxddmbrtbfHEPupDE
mMg6EJId129qDstZu9k9qJfR/i16wcH6LU1CfbjlS6JQM6xLYcQYF+GzC/sAY49s
kHTvZv7SBlsDuffD5tut7ZMYrVLRxhXE4MQ+qSHIRv/vp7+/EUK5lfOTd2go07EY
V5x8A9tIyMeHmYy+S22Rnx2OdeBpCj5fkVEOlhKGBC4wKojPufWdSyWwrFeB+42W
MbpbnjYyGQiDJemevGHUeHB57IFNgjxjcJcpkmOg5WUwLwVbx2J0zqLFSpznSU5z
9eNQwCAQjO5jSGOpRr+oL1gsFzRmHLgiZzZsbpEOt9jXtIc7hASi0EWOAUewunEJ
cxAn3pPYQVJLel/u5Q7rUcdEbN4JSqvmHmqf6bAap9V9uGCBvVuBS5vXB+7HDAav
0FYjGTm9w5G/+CoEeIc9JNHoX5dACRdH+Ah5dSkNvQS1iPZzu5+pxRCTLfRPz7ID
iwDzjq26RPatAfS+sNiTROUu1WNM6Hj/jHoV9h/comlK4T5W0EzhBo9WsaFCjh63
q2xQ0Pjxk8Iu6JIcGiMaFMJseqQA05aTgJ651F6ylSu5gEl3E5VVJh2DvhmrkWVh
1MdLCrgx/UoiPHI1f+ORBAXw/CV4Q9YhchXVO1UWZ6EyH5wNA8H76n1UdW5vu+1i
RMhKtM0X/ZjS+lZqaHQe2i75rmSbSP869td86AyvA96hWTE+VXuJAn6v1lDe8PdE
TQfmYJjRUQaiHyPc8QkK2aPZKyd+VuQHh/xFgJvltGWFU/+/wMIKZYkGbtsb+IiT
Pz9flr7LBGyerNuKBU6EGiJjJ/JO+4umbqzy+g9N51fhV6SbSY1KXF8tYoUefC40
OvBbJYZz5yZzUZ94XP9f8DVhspQf0Wxq3cwLUlrARMQ2KDGmpPMx90B/NbHaU4qY
3Vdm+5dGSffljyAcZFf7M/DvbWqIUzqM2MxZz5AutWLnjvQD4w3+u/sMH7DS/oe6
Lk2pOnmF6Y5oseVSgSxyKP9KWaqvgFYMm8HRxuSVdrZzmN/N9Q4ooA3YqYImvQTc
j0WXJg9NBHItUaDJRRlHBHPqHgGUKoiIWU3EOg4zroW5dao92Wql1jbjiqsR3frc
nmkVZj6jQH8KQKX8BM6D/mCa9PR5iQ6t4oEdgOo4V7jhSOHez2rRKFPnoj66qpmn
5v9Iq70R5VbP3D4SFjao3NLda2uevdHTMFfCYEmObBBjObwKsZhM69RyUCDb8ZG0
wZI/+KSUqAmmCw2dg+7cg8xb2eyv7F4rr4Jgh0HYc3YLFv8YenSfUmNZfK0GrNQk
24pum4R2GEdsSFsDlTIY21M/lq8r7jE0QB3pWAlC0h2JNOrn02cgKyG2TqkXmzhp
CzpCjtFrtk0Kpj9iW1uilH/hBrMBE0syR/QDHGO813+32TxwftqfS9a+HsjvY3Kd
GW3f4e6KRMuaaHc44dGJGMbImAcS/l0jNZAlWVdBxXq3tqsapfbNtbhR6AyCYUEB
X1dy3sjrGD3WBhGnR0Nl/ZZHIVTBDNsY1feDvODzXdsD+EHhCyP1+kGi3kRoJLS4
uDJGcJkU/YyseyaSAdQQlNUkXflgFGo/Lqxj9Zuo3yjHtkfsoHjq/VAsLRYMznlc
Y4aqpiZQnw1Vxvm8AG5/zqcuWfSe2fYQi5bDzgDPEY1iKC5yEvBDKJ+qfzfC7G5C
uTRjvXltJ4oZQeof5nldm948iIoVuhSV2046MalNDMqa0OOeMANnLGfYgyUa+c4p
t1OCdfRQtsB3gTth9H37EeqUAVR7JvZIe6vGn3ODufIKRrL42l8uVIuZEaanz/AN
ne39mIPreYFgaGzSzWN5ks4pfYlOdcbvgGt83Sj7qlM7nMoFWHlPVI1eSbFnmKMV
Vr3FJQx5xP+m2DnKxQuWT+YCJgjG7bNRunQ9pqVZWox6zZhXkT0wNbaWeXeQF626
XWgPdws/yuey2yQxuSnLpJ7sy3DjAZCjKgEo9gRG3/moX6b/OKCUQrXXCWsULAyL
aQzELqe8WMil7n150fH+bQOdLfecRQxhRJBKr77FNpv918/p5mgFPqLEUeMA7nqN
3U3k1SbuW5RhgCZU5EBkQUnUhbddHzQufcG41LWNQrvktnDS/GYFeKNq+mqJDbGF
mVst56PQtekguy3JptxLWhtfeStN7cGVKBNlC1lRC0rAN7FI2Brdwl7hDHxC9WWV
/WFQpt7YhxFwQJDPeTWRs7+rUwHBjLTYgkzSBNg7fnQ9WH2VPcn5CzBDbVIglA8r
0kukZ3xIoEaIZ+KMve3Ykv52jxMLsyAzn/aHBT6CCfoTixeU1wEWSu0AO3oCo7IW
pCPErhcMjrQ78zvA1LRR9bjGtotIFg7i/qeD+h5mUsxjzDfPE08sUj75H1JMs4bf
UO85RWmxN3ML6U587VMuYA67ThUmT8QR9j8iSOV/o/96XLdIMCyKeqm5lqOhgR50
cp0Cof0d+5AbImMtcuYKXCfqIdokOmPUzVPqxBrZh7dwhZq5AnG0N2fKrjIfkxXP
XWhVbIip/ErBffNqsITwDSDBrDzx0wZgUhpUWL12E3Nz7fux68IY/+/DfACoix+u
u4UoTpHMKiHS5wvzuCMrMqlf5u2nENRLBApiFcNYyqMt7+VAgGjVUMYNZsKEgm+P
MNenN2dEDXdYxF54GZV7haRC/UhsTrQIGbMe4JZt5YD2L47hhnQA9iZUAz4VwpmV
L+O63S4o8ueOv6yb6XGI7xX1+bJ9PhQ8UHnwTZxFNr7kOJLCWCxLRr5OTqa1W5d3
ESo162QiA1uOLuoqyZfurSvjeBUPRh66WlSPiLh3E1sAdHoU63MAP85xwiyblIiI
d7uRotjrCKsr+BoCnxK9JmH0AoB0Z7ao77pEpcUZexYs4DpZnpF3w9mn7kZuXMro
d2h7akitrimYcb3gWjo6c1CisvpCR9Z8WFaB0K4h+imMr8ErjNmYw39RGcQ8uMPa
tiuun/Hsb0IoVge6VcD8MMiquiPxrAK1xxIVGmwtAx+cOV62r3AyraYbdEApY8yl
iobTVSzrO+Jz+UJf3iSTAPMEA1WINkTeGnVbra9VIPfUaHZTFzIBG8p9uJkGNJQ3
kBCy9xVnlkymoHnYnnSv6LB9QGW4GeCBC/UTD6JuxaWUTPHedVeYQkrrxK10raQt
76ZBLZGTQW02eqcs3NzpURRIBBfKkAjIjmhdemQs3StwGQAEmGxg0aQYwiEOh6BC
b22JoWF3KwuT8IEkuQElAx3ZRVYiWHBkmrppjDbOSx8zZrvMI6wQSjCsvF+vleWM
2SQLYM9P2vxUsqFwp77NFmXZkgX5P2W8vPvLXSa48zLKh8H5m1j+i22eUqTYnIgU
D30mBn+CDyl7cGgaGasYH5Ad+qKaT0ahR07Q/w+w0ujY2U6tAJW21l4iiefA8njF
U/An/ZCVeV10vij7hjJ5uzNjzp2fiHNnvmOX8prjJEdtfDm4BajmuLaFOjoFZFGM
5ZdwBLBs+ZDEalvYVGqqZ8TpcuJTz9khihYn7x7oERk+iOtOHr68/Pal3g4gvyYg
fYOwzLGOqrfONUfLpvCdFRcg6i+GqE/Pxo2vOiVTKKPAicAfqIsgArWkzrjqZQd/
dXlsefq4serfpy3NWitDDr94bzu7Wf054ibQJSZMgYFZrIGtTcMR23d9hMQJRWcK
jQEo/X5Ixouj59EcxpOE6EKrWh4QMTJoystyv1/NsWBdcSq1JziwGZfYYsh69xPq
TAfNsVpGU0kWD2vydwW0htEoZJF6YvMelgdw5OSnX5NyKZEtQ/CBA3kTy9q7WU/Y
oygVtuJUbPBGnnD8VuLZST5lPJBkBky63oeJVGny0dKazbWO/PX4DJ0mFFBjO2U5
1EVL3gAkIm16WeOOzwiEC5QVRlx3nkO41BFYEAUT8NrcUrV1IfDA+neL/jQaiJPy
X78rPjoOBsCy4MASFB7J1mvdIYsnbvItOU24nEpJktSryfF9Gp4pHzfaZjlb/tIl
MnMDoEeFe4wgvK+ww2g0AUvt1ohhgMxeoJEqNVOyFBzDf/ev6txTjJC7QG/CPuri
RR4BFUHkFT/pN3gaC5xH0U4B3SGMvCw96suxuBhCoQnboAqqrbPuVr6k+5LeY9+w
zPdCLtFcS2dAKo+gKwXpN6nLOj1Pb9xpWmfNAPabcOVwY8W0vZ43gv2TMkp7FHnW
tArohTxyRgtjj82bqtIFJPKLQrWEo6a1qJE8+NVjxy4MNdHIw+Y087bJ5uJbHqqO
8DdLtZLAGsSqa91VejhbmOhSGu6J/AMCLnHgkQF/cZTxxpDuQgNg8FAvputMAADM
GRgC5SeoKBpoyu7AKZ0GsArqUwZAXdlELsLhNwA0qDa0VcS2GC6zcy/bL/3Cz2m/
9wiO8HPhCNqvQPNd8fqOvsGlkbyqpW02dHrhYVLxCc1rQ7th7TkzGokcR/Gui2g7
xivGmIDxMRoX424IJC0Zfpqd7JeFVjaXvHZVH9IC1ymOiLef6mGfu8QW4ocVfaHv
ZHVBEJZ1QP4IO8+Ll6VLSt3gvl55aBecrYKVc1wAoV2xmkLtVLptOsQLjgLc4MHl
L8vgJqzpg56nkeORtskEtZg+EmbmJ9vMOBbwIiN/JGFQMbwMW4ghEQ4I8YBy0wie
80IiGPY6MQQxWvf7PTVIbbbfTREzn9MyvlvKbSaWthY3OCKluqJ5dJBuK2/Z8hfc
PXbG3wYEuaavfND1sW/2Ah9Odol05Ri/xbxa+VV7qO6TmhiIpS6DDVLxamNjhfsc
p/Q5y/Rm5t7xLc5eGF+oRX82SXG8FPdphXQNLvL2B7v5FZdWjrssv7i1ioCwqkug
98S4fhIsOjQ+GRf2iCVnSCF136D7PscUbkp8qpb/NVrSp5Oyq6BkYtWRlxFjCTVc
tYDVZqnV+eovIg4E/FtKEND4kg7lwi37pAj8JZYhMXDw3tRal1pBxnWhQRNre46n
zy8Pihurtm92YhxQbNagVY/6m9QeTbDZ7igHnVouAS/fCIcN/EOw+zEQ66FyFRUE
qkLHafEfiw+NRqLm/GU611/TleehWeQ/35KHCl/rjGDFlJrACAS3VT47mlUUB5ZY
2eASZ7+XPi2ZnSzNuJ07hm9xMb/1Waft5BC+tGKBrrQqBanrPAamAJOqcKZaKcGu
jAs+vVjgcfOWFM330FO3/OBU0eGFBkHBNCCpN1zzi1G1Ejd949a7ERDTnKRgZ4XJ
MtNdsZoynOOJy/eosGgqSYtkmaRFr/NHnAiLnIxJoJHzaFIR6w3RqnpTpfu2wEuI
pWI8cOTrRzYU/1HQDzd3G3Xn6L4+p/YmaKkXmi0JIzu9nEiRCehfzU56NIq3eZAP
UxcvNapAuO6qpXCdN2cd86h6mpcgqjv1XHAriVwguxvMk/EvmU9jNg3g7TQXpLws
1PqD+L1i1AmZRbimC3hhifj46iPyUIW5VPLb7BtvpGFAWephDMNDriMROGN/Fzt1
ySNWSW2w6umGL740lc8Ol/u8FaOgv9M18SbUtzZzW4KD6xtbuz9mRZVj6WV2zx24
LlgVX5AsNUiYzGYj109a6V+JETdtkSuq7T6Fl+6cho44CksMvnajXzs3ECxsOIJn
1LVs/30VcL1xpOR1EYkl9jcc9V4sk52pTfwWQK37ZGj8kh1nY8V96DC+A1E09XX9
ZfiPB/6zMVTI961O0hOmSvMSwN6m16o/SfRCRSjBjJWh1GxWHRMDGq8D7EUNztgo
8Wi3gbQ3V6mFW5APONEcHjJ+h3bsPOdB34PqpLIVNQo1FGuM9l8qw7L3PSZMkGeN
yYdO1PTo4GjyzBtHdnpe4TyasZYg70yxjI6cCSwXuEeU3sUORYvMWcXh+UmNgl6C
UOLU8fMnEQMq0ZDXFj6h1xfC3iHPkJmwnIXbnrqX/Bg/nrk2uBEbPH7iO8YhsdB1
J/JOVEBVfUjtU3AscZXY4c2rD26XQ/4zmdJG8ORUeZXrFd8+PbGMPpIZpVqgCSMJ
byq/aMjMKWC107o6hI6sz6+wvQamUNe9OMc4CH8UFMy2/CnbRRr2wuNIIUiwWyIA
3ZzCFY9HcrGveGBXtrTJJUWvm0w19BzJZ1JyxIcobNmhgYUzd+KWk273AlA7OESm
rIT8c7mVrrR9Pch1chm+6iJzB9oIj9yuYz0StFcEawBn5bDN906qM0v75X1rrVVL
bu6nIiHK6Iju39IKjHMJ/LyHIOuAv9OMbNVbNCH/R1fWsT7Gzq8y+2gpl20PKggJ
4pRewS9QaxpGn+CAwGVCNgUTIs9jmNByfPHU+Jmi165aSvuve//46N+FRBOde5vb
zDx3B8Mg1s79c7yJPPl7qhY+WYt+YXJzeRltbT1PXR/nQgMw0zPexVOmsdlkeKQG
YKpXtUfaPjXR2HKIrsw1fXSDHufR1rOwCmlzKrmiWnGEM8R/V/fI/MbQAShsl10j
PBn5ZXwi46GY97qBt8VjR/+slUjq8hY/KLyMMQB8z06XNX5yoUliR3+NlXQbLjP6
1zU0+wUnBIvzloDfSVU+cMA0FzCtK/mSHvfCEz4Ufxm6y/IPNg+1lqfZw3kfBa7u
5JXVGyUeZ7lLUYmYUmjs288KQYnRRhCXy5kTtvkhWj4hPdVxqPQSWxjlSeNr1nPj
DlC2PN8MHBL/YJDshCt/jbWvWiP85iEMUFJg9Iu8Se8WcIVWTltfG/rsFMfTOvdN
6F1OMYHJya8ZDDx510fbWdrfym6xJcpSLJR3+Z9XWLFKr1DJ/BdEAIKIxHbR7M9b
4ZTOqhFwKQ30soi/qGh4ZspdeiPW/cAPlJq56YseqwLrCl4/nd/AWgrIb71EmOMW
dUqlJNBD6eJyQY6MO9F+MXrs6mN+SQcqr3xgR062fVdqwOws2k0QIqc10yLDrTYY
VHmsc5UM9Rttv14RI4OXVDw6YvJgFMIkyqPTlCUX9bvhS7ebEvzhqfs7h5/tU5Uw
Kba/yr4xJOa4onkih+6UAKhszeTtB5p6j13jffWgBg0YZlYWp2xm332kV+Z+/9AC
fTFyfDz9Olo0qjyrCCqNNFNvq66SP5JKtINH6OILQKFTXLzW1GpX8IE4ukjHes3o
93Is758eL0fAHEQFMGFU9FlK/WHDvBJzO0MIExaz/iDz5+4vZZYntROPivEtLqhQ
mR6QzBgFJyVSOf64zNsLI7k4MXu3kKaFsYICLuYHNf0Pkei9x5vYNDt6HVRZ8rF9
93Ap/QopeSglRRDsgY6/DRJP2zwRzqm63ofDQ5+7G6btlnhdCzUSKcleUcXGlYxK
byNs+deWCIroCn4mfmf2TOo5h8lXSJT769XpH0yiY3wukD/3whFd+06TwPwH5uyt
POg4bRaVF9uDULAxufQ4QAA44U+OeP4zrVMLwd8qiNzcrUEYG/iwWanpIpd8iDcW
hoifvYeqzKqTQCV2OZnJLVupWv7SA0+bo+0Or8pLobgefjiJZgwotRZmWnydrAP4
ePWMdHhX/rVLHDHzslE+zVDiHtrMKp0JRi+UvpEF8jX3D1Xwg5jYlPH2SI22ofT/
8XnsGMWcue5HJ6VHWSMBwpNaqrf8CaMbWIRZRij0InJ/FCphiZaoaoCEvZqO4s87
A8Pkra06wyBCtouRJXTU61coJuMGjio6Z61FIcXgiCfgfsTBBpUAzENMUDCF0QJy
VGv/7GUaiJZAEPvAqzWy9sAdyYdhos3p3IcsVwOM3cZ7WPxYEXqdkb+gA1Hsh/gS
nHbU7CXHyK6YyNVwi2WdENeJpHFg+4B5IHACuEDSwMP/forYTkdswwb02TWLKVK/
XRxbiiKq8rQOe96PNkFLfTSoPB/7vQuUXt1oVYcqoG4Z0rsK4hgAWA5JjZaHoX+s
PQvGMh/PwWBzz/k+pxOZrlxUL4ZscD50V1SZnF0o/IqUafpQCO1/wiA/VPFHkjz8
CUaCUgqheT1mDbYU6VenZhS5NX/rh60RqdHaR7mAF6OuBZ0PsN/EC1Q0U8S4ySMI
ieGeFlDP/k4nQjvGKu4n+mU65jaJuF7/zOnZfIdYpY36UyLHWwisCrS0cQRci6eY
1NYa0PyPNBJ1kWSl7LbH0MnYJ2fiBnE4i/hwlbqPBIyjWP4oPvL9CfwfHTIfm215
qBoU2FxEQ3YBh61JuKiqAVa7VFq5BpNz8oSp2Meyn94ZKNkJUMc+kAy+dkjZ4hn5
KJyaIcpCN8NcJKOzwio4iWyNKfQQj7ScwRX00e0AczbhMZmOr6x2LNXEvVfHUIHB
AHMcuJohrM9atXEM4ouuO4l4Mx4qkjcC5UBdGtZsGRTkEIj70Llr/QBPn2jQM1we
2ow+wouBKLoIvVQulwjeQYhZRMI3X0L7K5fDw9DRndAHkVYQFDw/dpc5MyuLQzBc
qE2SyWqAqJkodGg/8U7H9quLJZS0zqYeB230NeiQaeOPypFEs91Y2RUmSY9bZiUK
KnlBbfFWuSVdNcekODdcx2scIvRZDYxnn5mIfbgDcbeXDMTy+x5GpVdB40jw/In6
F59eGYmxSaLNqnJfn1+DKJnNLgSrNLjy+8E2ztv4M28YH0O6Or9jqk3TRg7ZjXtK
rUrLnCxW428Qlm+9s/IjlUlbxqwVYXOdhyAR5Tc8aP9KzlDopQI1N7z6EdQecvqs
L6jIROTzc/HcFjXY5mUDR09DYd9C3IFpiKaVEhiJn7HsP1NDQ79lrl++lPlAa2D3
w+c4AcNd+LvK6LrUPi1yNI28XLjUZxtPLo+HPBrWVSfYug80YsEcWBfHC+1nVvKr
uVO7UxHBn5HcR/aaPALnvoYBasziImX/OdOszyDfIkamHzLi1uJrS5Qt6PREX7MO
9UoBZp2n4z86yQBiAQPyIQsGyV6nAQo+fCbqMPqfAP9GfFPQaw/UllpAzqrhEUnK
kqGqXeFoIeQRWA9wnYIDHVxhCBvtVY3f8G5yYr3YDope6bPdQxYLqTtDQOqqKHuD
NbrL22kX13RvfbSjttWRFgxfXP/T6Aj+HwjudasCmx949T/9sQykp3lWNwzrdJQV
oPIG9xMm53qgHCoc5hWLlVI3qzb7kKirz+N+C/4v3xfbLYGxnJ5B3QsfTT3LWOTO
ZU98n/JeEPROEAWr32+VJMMRTVterLtxHg0L8uvh1cELzs9adTbXuCd2goWptL6+
aH/Nhsdqn303IGeXAieNHTVoenL2LMGL8kLpvRMnrd7jnLU+tFGC9c+KF4+90Vgz
Ux+ub7iAmlB4RJ3+REttDHtFxtZ6RIO8V+R1cjF9JuGjIVhbLCFVPA6WyXDDrGiB
23W7syCIDDbDFFYo/8keScS0KcoQusbD1327pTZXM8i/VvOvtwu0ftNHLsgFBUjk
AWD7Yhxsgn89b3QML1IwpK6AhNvXOgte0QDy9HmZj8o9u6awO4b6UcPQu24Oymog
ZGflCXjdSxrEzQwLjemY3/44tVso872d1FG60FP0Ihu/MhT8Dhre6yqdeXOCbDvS
nUws5W6dHD5N1voTYWCAJDErDszpiDVuUAeb8s3RCGNb0en0cMdI8R6xjLzl/a8n
oVt2UjmzT4XFZEsobTWCxVgUDwptil1pIRjLrgRX4ZSSV41XcIdDD4+lywPtmQXN
w67MyLTsTAm0BACOn/fT/ILw3Nifcg2/UKOctDoHHv+kTFunZG87aP+rzoj291J6
abMb0di3RwXufQIvVIPbCiX9EwhsGjz3KGPZ4u6BMLDjClL4LSDBa9o4e3tzsYIR
tgXxi94sE4/aE0nrpDsGBj4Nq2nHBbJOswZUkRlbu0PosuKS/NbOjD6/ae2RlwlM
xBbnkwIY9li1h8iqXFRMplpUjG7AhEntZDKxqqgT5AurZytWkWgLb4Gkp1sdS7j/
6hUqIJ8mUS3Ch7k62mAiKoqI+/XX00TtLXkrXBw098HZYd4VyxGq6J9dNLZlpSDh
EaNlBSvfkGUUwnslHGockHkK6W0pYLv9MAzm+52hsIhylv7OZkZx1HRc/vBhMlma
T5KtGsBVShDtISH7My2fzcsUjGgAlcGUdBahkVaVvQ/8rc7NImD3JXttEYgcFGP+
KKbvDJaedec4EaB4p3rIoKiKwnJwWWmNEva5AbL2wRaJar51/cd2D3d5YYKXBN0d
v2OauvC2dceZQkLAk69esBSieNU9fq1ZyhepaMCxRwYJmIvewCbtkDcv+UATLWWd
IW4w6q8eSpOXB/WIdvNQQWBgxSiCwap10aDPOloKBSILCVR4At5owpXgE/CLn8tQ
wyh+WDMKei2nEMCINUWBo6yW55um9AYmv+LaS5s1YMobfOKUvCwJsGePFN4uoWT5
SmepDphm1kORrj9kVqsLD0SI0dKqFEz31QWMsP1mIlWeE0ssJabWbiYZv0ZbU/FQ
fMves+7nJY/lX2MZAuCZVjSe7g28PXLyD6caqBtN0M5eKxX7dIs0IWvdao5389G8
Ngdoh7q3nC2LdXOYyRs0Y4mF/DcvtIK1Rp4IsxZfSdk6czjEq2fEmlyrPOIuV981
+0dm2bvRHEk8CkAZYsXw9K7KdK48WFL5XIMDJp0AJjaY/vULhIcoelbNuvAKG4Cx
IgZyx2ZicN3RwSqY5NsWZoH/CYzRCXpoGZedZ0P/vDGC4o+L+v6jd0KjvX1J5P29
R7gOqf7a1QtTdNH+C88AIYDssTwSMMgrZwHSPtcVX789mFzHXS6b7k+gBPie9+O1
EH2o8zYxs94s4gfaOgEqUsc93QGiDaNKgrSov0qtHaAgLKbrxXSNPNj1aT1dbnM4
MgjMjFSjBcX3e6PeU2S+nfZHH5ayiURb5X4Rl0m0HZWzCZw/Hjg6k1wk6iB3FhK2
SbKhDrxQ1NWUzAMa1uhbLCsnIw4xDbnjGO0YzZCYyOlMu+6APsJnd6EchYXFYhHf
2INgj0Fxd2QCw2khq9Jv+nxreKYFw4yG50dQeWFV3EsbEOl9XXUUFg4N3IdUvcrI
QRJ0MXIiE/HPVh7+gKLgi04Zg3u26jo5bROtFQ5m3o3lxQ2A3WtrooTm8H2HhQUB
F/+536uKe6wfL5nxuUn1kCUC10ByYzAfdcPmtSSIMmNdtyo/h71v9Uyeo4gf72TJ
0en0Ofbsgo3AqujQQQTk6e+dgdRuP4IuXHjEDui6sZQ5VJ+PoDLrO0YZfEUEabcg
Fyutk8TBnxKS/GzWWhNZ4+41xXCX0L8TUrsYr50V4FIFPdoUnLmRsqIuuWrxepDQ
gveTBxt1C9lEzaHj2LrWwoO3BMiRVZymH5PjY2wsv1mx9iZ7DFb+Dk4+fQCnIEWD
rziAyfQ7rlAJ4fdCY2ckTR6AhcybSjQD5k3fiE8/IstVrw+mU3kGhSUHxxl7VyFP
PFWoqA5QpeCP18zj8SUPPxtbWhNIYP/VVcaajCNvQMnZ50PWOn1FWGsIa+qmouGV
BfTEF3u71Ns/8Jfe0urqCuoZ+aGknckieEv6Y4P1b67aidJPXlrXXRFwHb9u8HFN
I4tru1a3asZgOOJReC/VLuOpIjLZSSJvFCdZ4GHAim6Y4s9wLUcp3KnXKaCZwAU5
rC6iqpVm3rDJwtlDLEful1yuhfMoVhpHeN9jwsrqiXlOqMkxSTBNIsY87Ev0Z/Zp
3gygkkkuXAd9+cbdtLgTYjElXXCo4OG6q102BXUVYI0vxIzZegjwLcPEQdgLqlGx
aTLpLiL2updWUxjfy2av1tWE4T+sERBLRpy8kTn1G3PrpNP9xDZncuvjvpQkjZsR
0EVr3hN02iV9Lz0LsHcKlnDwn1HMBIxfM/sJXOxkZMFNwFkQxcvl5f39ddypAnxs
d0Y23jiN4/i9TebgOyjmx7QU+fvXMMwgytvIi/fTPfi5AfItRc6PRdQ8KcojJzBX
fg6g4XTTNpqygnwhBFkWbgXqdE0ACI/kCTqcXrOY/oif/LoBUlV0OOXTuXgJ9NA7
Tu9VWS/4dzs8ws+MBoW0Si9UhYvp1uLkWkagw0XFfztTuiBqUYh8wDa7xWqMNuvs
mxkQP1pWV4+fP4cgzSdIzOciEIpka6ewIYf+JSVhYCBERUEcAG9I1RMGiunkwb8P
aDKEUIZN+ALLFhgInqTDVh6TwFjAqoSIuE4KYA+Tz+7o6vYpTuOBw9ZYBQHPJqSl
2ojEZrhX0unFPhwQr8HPufDPqHvNudHPoVjNMB3K/lent66txfH/Yof5oGybjCYT
VW4hBWYyk3inGozKL2iewa+KZw16aZ9eQqbAEJT1vZvRozYs4EGHtOZdfOpwpv5Q
QdJtJhURhrDAhLpTUBGYgcB+jfr9dqTKIVdt2+knsI2/xTt8cVsCTD4Dj6iAqSjF
dGCYnBKF10V6hznNQZSjv7B9M/GMKxd5hjrCVstflBjpaGDP3a7Vd7U5Zer4TOH3
I9srnTY84yGg6DOXkfsTvcIhLVFUZQRNZ/jez+wmC6LKGqdHPDLJVE6yi9XR+ZTc
chfglMXcVrr1+ZADbBmdwBECHC1wLvfDuDfnF+Z7+fmsoDVRyS+m0WYE85c4bmis
RmZXqo7R6XEEFEJnVQHh7Hl0hNgU5hAdqr8Dj/YMU0OX0ZV0N7f51gyjW9v42z1+
DDoCT4f230iyLuQsBU50e9wdBa8IypYF+wc89doNOIhF6YJwOYxqG3K6zaEcCybI
akMQbNXB85JQja4r4bJxw2Gj2wrLkVkBdj3sODcsbVXdX4zeSMDRIrYE/2wPx+pJ
4euu2RiULmJpMx8D3Fw5Cio85bR23lgSjMSf8aOa4a46LQPRBlGXt2eS1sd7wnPV
++p83owDUHfijwEJ/Nf5IL3RaLoz7ldz7AOsbgvLDLDL8AvtGhZYHviV+Vg91foc
mLjvYdQCIYzZ1PQ5pZXdMwV9uUatYCr1IFIV1U2lqLzOPJYP6Zzw0MwfPMlfKSZU
Dfkj/YMfvw4YYHTcbccULntrmU+3R0xQ6jRDpR5Xi7HicwuyqXs5PAN0blwXKbtO
UoH0ha/0o5SsK8JA1JW2nOxX3r2Eq1e3YQbVHlNeu9gnsrNgjYpUaGEIn8BC735/
K2k4zGFB2Smqg6OhKH1W+pZmcODKrJg00y/IgaR2fJ5zbhv2C257bgBGib9ezV/L
qB1arh11/SfqpsKzjr/w+APb5NFCE4hHiMM7QyV1qWMEC0LRLoQ2COdpW7KaS4qO
zkPfpwakwa0SvXYXv9EgU+eR3cfpvhmZVaprg260Jul0XarHRlOrH9WCJdi2GbqE
E2+q7D3AmPOSaEI6BMC8tL+Ydmgwpwy+k577oS82p6iaMIngMSpv7At4OKtFXd24
+qPihnYBVKyo1uWdxCubYwfc7mcq9QZg3imD8L89Ggys90RHWcLfntaQQ1i/Zmpy
kbza4mxaOsWDEa64sYcZN1EKvp/2Zbk+EXEhq6+CA2609gdUYjtmx2yud2G88fBf
S0ODWrcBsw4k2Oy47sEnvtrfmCZLETHSKulcMab1s7jrTaJpZSfocyE2WlFsTpWf
l3k2/OhUsp9fFPQuRG3HOjAR4PDUbNWURjoRniLkgOuLs/mz/Yym1O/8o+LlKRBi
9sQzWL0ZFcGOA+gkhVbvak5SKX1zAnsBAUzlIVo13BHKnBST7TQippdS/xoAYNjB
Vc1bZvAYNzMSy7zdFaghcQYMsdhnySTq5pW5Y7koMhiipff0WWFTeRVltPk/w75p
5Shdb290LlS7VULiIEFRRjZ/2ilmQfAjjq6H5bIwarEbrOo1raTlGIg3n2YTxNVj
Dmbout0g3PlPog3QWGckGa21EuEJcba63rJRS3NRuicyqa8JWrMCTQvyGNQ4XPb7
/MDNRtkH09Kb1hZ1D2KTK1SWUs9YD7QdYw3p6lmJDf0fhX6ZnJv01u0M+q2HrXH/
nELEMAkDRVVpPD+G6M8l6t0vojU23OZ9mmx9JaiA/8Vt1J4Wc/HDMrgDA3M2XDvE
tsx+P8WCh6DxjQbW2wTyGuzlYPvAXvOB2Gywudmm+mBWWMUjL2EgxHlgBn30jA5n
GvLws/InFSC0opwXUxl7mw/klh6JP5vjkVsf57x66MaE4zdRa127gAEUMsts5ENj
JTFgiYWJja+Y7oT6hFu59MKwVxQeYPN7L3qJFVZ2fHQ1Gc7ug5XvSvXy47Y9Nc3F
E1lj0ZEo6FNfc8yrvQewW+mY2CCeTAsuX0Pfr/3ac1Sdku7tCRhzsMPxBk7p114J
tHeSLeKu7wl4zhLwFyReJi2NqrKw+lmEV5ZeeWWZ4aqHv02lkJuIYLedwCkBOuFU
9O2pTBFBycNAC+8W6ytmSLslbrQTEkluGrO5QEAwBdAHy8JAv+gR0/+j0TrKNBQ2
/HBpBoxlgxn2eU0rgk7F3XgbDf0lN1Izotmm7AOLUr0ztv+MltQ0LKzlYxj8gBvG
6T8dCYCo0fiJjvrkTa1xKZU7VzvR6Mw8Amtrk9tO1Jfu3vHYeYUBnhGH8YiYsb6f
xIn/rrv9401fohgtoWZ5voXZk1pMsE/po91/HVVJJe2G9IqjR4a0NvfyV2yBqhkH
cuhj2N/U4Tl1XEUbCQXwNWqGOgL4kL1L9IGau8ubhk0IoMH0XrGBbmQ4/9VTBLmA
9G7WUJJoGI8w3mBlu5KzDqKkzxS+OnEWeSNkHcYOk/hLugIXnXDuLWgwmqK7WsRh
s1BFFT4jWvfV2y0kQ7Mb5p/DxdxNMNTsnVzrra3B0CnVjgWoIBgg6eKJMBA6zSAv
Y++ORqlgn9yKQTRX8u5dx2d4NA1kjZdxcT2kE/C1EC8/MypzxlCsmbv4FpyIUkwF
FYuZfX2BNsE1wdPraVNU/EKCgKL+uURtZBwUZKn7P5xAeRAQqi1KCBEY79sNLr4+
tHFQvmMA3u77kiNPdzZxzHtu7WlDi2rBeb7j7NJmDNNmslcxZiov1LaEDJiI2wv6
4fOIcRXFCa8waWdGgHUpRAD3f9a7yN9FmFBKSnWxw4FbTdQJOoPPbo+OWXObYHhk
AEJzeue5+BMEmut6JvKXXlqpWirE6TwjIqnf5tCp6J2UjREyxk/4s1t31wWcq1m4
0GEtGgvh5Wa/l+SUs3VFo2eAnXj9UKUtOZ2U0v1rJjzNvPuKJtPil9YF9BaB9tdH
qjQNiwdgwosZSFl7pylBK+LrM9dum8N1ywcqnCUZkyEm1IAK6LoRDkTy+l9C+CR2
iWCxtgvoQAJcN5jc/6Uw1TRPkindek/krNwRlzIN+LjsQOYK2nyU/WIQD7LfQyhv
E5jzFKjUN5eR7QjtVV46ulRLLC0VBETYOLaZAtlISWuBoVpTiOy6HTzlyKm9wbvv
Q27ot8IcXokhzlgyrPqvnUF1UiRK9PBuzcxqtKyijUiwrB9uPU89TIM/xtLONrc+
2q6vyb89veCCIFqQisJ/WyDc6FpXWwPpx5VYV3NuuKj21cIgepeAGPqvRP1yEgF4
83r7Vw/5ZKngPSPDQOg3V7UfwMdyc2bhneWrlgAFNZmNqnsu5u2Rm59AQzX0fgyD
+Kkiiz4FFthtpg89zJ5VNeeIMSFlR69kn4c4/ya3ik4mhnpiFe/IbbPD/Vy+OmLx
8r74lfrViVePT3fZl2nHd2Z+y4hPnZJfCq4Kld7Ahr2nkmfKMgNCaHETm8dji2Hi
qvq1DDH/KhV+SxW6GWFcyxeQ7CWQF2vpAaZskMpHQnar6HvNQiB9dS+AdNnkc5IW
P7HPU+hc7fX6SH9iwS5MA935BfVniWLMnlRKBcEeJymCaygcmKXVXm4Prx3KvlBu
hFAuVOcTTQTKzHVvIY92aAp9ub2Q4YZv4FBxYa23hLT+c7gYeu98th+9inlsDiPx
kMQjoyLBXwpgXZESQG5ShSie6KAVtZpOkdDMmPRbA4oUwbLVT2syn7/oVN5+6bP9
niaAFbMC49ihu+M3vX6Edo6cnv17XyfDMmPYkGT/COT8HUXGTzn8EJWHd7HjSeg4
B4wMKIAYhkw79XDYs5pWLJS1irI/Gpy4nQ0FZKcU0R9TBtyHTJ5ClWpnhMeWpBO5
8FOp3lkYbwuTBjwAx9NYdkbEl9LosOehlJFaAOMZIFUQCL3SV61qC2dsN9M11jdq
FP3w74dwgWL4RXwdF9+/vnd4ckn9vxZQcczy+RcUrx/WYqiP7Vj6/ah9y5jUCaJV
sjVQx8DzejeL84B0XnLNnfUSerEm1TvP2mBjQ1I8YGkb6ll1DIl5ryT8ZrGqv833
1UEw2tmTc4A6tXUBf7QFwUscpOYwm9PHHOyMCUHapYcdIEWM21wE3XFLGwktcXO5
XrtejfyU8DV5PBXL2NkYSC0zZEVl+fA02QOlfpyVX+FhEV3PJvamVpB7BTmiOsih
FIWTTM0Wbv35Q+xRW6xT6FaX1G+Bs4t3Asr84aAEo8YONLljKZMjV4iMrrCELIBm
v7/V1LOmbfK7zr1azRGb0LTld9Vn0WZflJ4+MFNRo0JcM3FFW/ymuV8aTVJT8bLd
fEdUqggUcZlnSZbyUSmbJ3d4AyA57FEzzTHB7aUfbWpXjsjQoiE5XFg/j71enGLv
7o8p7wnUq2MD3rd3DsOYRfE1wQSs+fFBmXb05gSaJaZtRIZINP4ko9h+u7TXXn+a
6Bg/FKeZaz3TqSvlqAIvs8haJSjikPsHCKGEuDzqg3JnvkEtI8V+Zejxh/qQFFcZ
z+qh1kpu8yYmDuFFBOyZBhHK2XnYF2Sh/Xp1fk4iWobrepfiNJ248lT0inSODnYa
M4mVTTo0f0xrGcBZX6cWRgHkP40nQqz9sZkF9dfVWiVtoO7kzWptZdQoXs2t/ilN
u7St1qqRJty67qqfAxiQIWWMN04KwavrwTnPKkkyyechxCW1ZqiyEwSxEi6Ly9UC
N6FnjkokUwtyb7yPXScuBHcOvsn9LB0weCSaDZZOC9zfxafZfzfQVD1KRIr/9+pa
2CrZh83NBXg9n4Q3cD/5wbbabQVetCenhlJbtd1VtJyHl81yVDW/6SqU79LrSO2L
ceAEz2Y9pYe/7n9ywhB5LhsmQ5rJ9vKGssQ8e/vs68hq7NwBuOFhe4kbIUxROk/F
a+6SFuY9sLc8hT+KqjIBHSKA/UMeAS9zzUdQD06hhn9MMo9XGbtMr4EFDDNtzYR5
WtXM9GE3253Thsh90Bc/I//ruGiFVbtV9dD00TDSFDILb9+eJEJ/dlMgp9/ZEjD4
MoyY7DZRzwRm/E5MXFouCRri1UQ0AM+bCf5CW81qYZm5LcMKXazKF3Gx6Gj4J+J+
/IM6Lt8nUN+1UE+lxIi7P6c3WoLVRQTP3npUiPImfVrySreAzlTTRNHZPYMQvTEe
YHvTZ7E7BLD6O4Sq792aZURm7qBKZLcBJMUcVChHYn1XzA2Zj4CpiLVPEevPeoBc
wVJYSdj0XGhhXhc2isuxIsn1hZ+s2Ohd9WQI/XyoEe5xXVsWsZtx1GnFgWoFFQl2
/IoJ47C4ufOh/UmWJLaZLrR7n0Jz68NkGjsXnu7f5pEBFLNOgIBWZry1+F0ByAUM
Q9Gc4FehsOUxw/cQAILw5n2uOJhZ8lio6ceh678S2gBG7HwJc6Y8q7oSlWi/yjj/
iyX/BL0b2x2I8TE+PMWjWiNps2YKLZ8eU0RQY8Q+W7B2JySb4QGuAhdWsIsgf+sz
znDip9bbTX92bINZFIFwAGw1TEdC7S49GkVB77pMUZE+wKFP8q8uzmKLLSW8HWZU
iHszlzEp5GfoVwdQnsIW8s1YEwnTy51M4vQoRvvU5MgRCAOrnWUOmP6a/+gHxacc
T/OoUzCGAZx/gC6lcwFwtjhedmKhcJb7IGg6wJ5PoMb4jPk0tQOVmy5VfHXidnNC
doD6RB1X5Tw7esIMY+9pYJURgOcYKqjymKSYV2r40gD8F1l7shHIrk3s12GAi843
BehCAld8ylzlCu1VSx3qFLrzdXKFqU6i6P5CxQBb5JYSI0XumesjOm8Jufczl/dP
Bwo4CD5cjBSzppzV9T550VMSGZ7qM4A3DnDTww8pk1O4TnCSAuCoKVXrRFbq42WT
MFeMy7fYMBaph4eNT9f7SVTFiEmSP62eaoCXf2JeWwFNXHbJFxukoN/Sm3ZHcVO8
ckcBW6c2EgyOiTERWZPUNq9kKJV38v752We8dndH9z3H9ozzbVQlZ0hpRKaWi/Fq
WO4cTAdMDBBZoOhDXB2J/HGDv/HMWH+NobhDnxNrbTi7yajKw4uVJO2kSYx2EsT1
/iea7/5bO6oJSH+DMeAyy8gc+uqvdNV7167fSMjK/b5dR9Dbig37StThkGRnr8Ga
YgJnCmDl2tppiqRDX9o9uPLs3qUk2LPE5RC72hBOZsze6BhZ9QRPIQkVQ42E5otv
v6jzbGhQRix6YJafS/iZbel0sdzhZgaGJQBEabXO2TI2jkPqlTRCYDE9ry0mmH45
DFXvXix9IKSV0O4kyN7JOtbaIJxzIQ0IAMjQzat2TIpnosBYLm56n7Gtw3IYacF2
NIPIoHTwaf2G9dJ26iigQ5jWVpxxtW4lsEXosVg0hcW7y6Fup97D+iIH+JWrynWE
M0VR1ogtVpFKyCxsdqW6TooBsfjb9KQMv5drdFOeG4NXXC38uoGothaN3z6chnhj
yTUd0lCax8h2FysHIhtxmfp9/UEbN+by2sB8BVll70mgIPEGmgNt1joLXl18HqsO
X0D4YL6NsoCGeJZJL/7T8fYRB3O4wCJ2FfbAy3W950Y72lpQUuHOo4pBDll9Qkvc
pPgvu77SEBjriOofl9ImCHr5MUnborbwxhp6nex0DsaoJuvQ4Lt8BScVqgT3RCWU
0/J461vTk3ztUS+lmufuaqhuOWdlQWlt1BaghlGKo94XlQptc/F8Kd4/s0gcOdK7
MsF8Ak1HKY+4/xPmopzCaNa/sqpSVmIsZBZV2OdcbRFjFqxizgJQgU6M2bQE0eoz
pGXhCrUxZzZze1sgGwLKaiaZSZZVLetY+4bqjY/lWyij02JcRidrp8n51nb/LG+h
2f3Ek60EkciipF/1PNXPbHX4dMbKoARWWI9E9oqiXPcR12l/y4RmXTkhH93m4r9P
Z3ix3+4yy1QEnoODgGhWvwBWVd+PociiKR9ZsCK6iog7p8Akz1XENZnOQTRy0rZT
6c4PmBCDGbEmjmgd5oY/0/l5yIOcPXRqWpxpJBDwHNW2F3ni5dWTDAWYxEWtq7XM
wBul48sNACjdg5pSx/fvjqSCIcI1oMBBDvqZ3jjSdLzXwC+4pgGmcYPFl3vHhaUB
e2zTkusNiPxNfGgLfPBi6e1OtNe7pSOcRFpZz+v6SmdcqzQep8Glh3DQex20KeFW
h2yDrpij4RflAtqs2Fk44smev79vvUpnGaaxKDh6BjmYOYPlp50XaBPgMBlXX6jV
QVgTzZ1hpIwMtXavJ9VEP95WrmdYbLOgl767UHVN6QI5SEw4kWzo1LuTCC95k28i
KDI+9gTrQU1Q2XRytVoagQPWDewjZB3tThJCbF+pvGH5YCGHAWtlL+jdXhLwsY8B
GytCLq4u/hvOXuoh53ia/BETXs7TB/qdFeyhACc2PNDt3ym3oqspUh2Odpc0Orxj
7g/jCO1RRXZ5Rf9psUhGVBRD8gSWjvmiCzfK0gzcxHOfe0zgPmI9Be0SpAguL0gg
1i/6ZSckddKwOk6Kmc5FE3N0le9evNF8v3zlw4V92oKgGaL+z3oYrd0YzMvZf2jp
+kY5NopAofKVfjYWgbpvYnQH+xhH4V+EHi7IFJfBrcAUqUVgswJJpjd6sW1VHb72
uAZCKu4QSg2st2w6b/1GDGcft+8o4/psgdqvGrfrFs+UbmLxKFTXUICyHcsLKSLe
nhp/8YHBl9EloAQwnOtsguVHLgD3QMxKHKZsKagRdVot2t0QsCyxvfZRirUijnjI
tCN6MTHaf8hyerDwN2S+1kEFuyYCY9MoPKQGSO3GyzSdE2uKHiSMUYIynKeC5hB3
Oyh8JVfuWZBeQJbjqa9g2PeFly+nmYLOkkj6BeRyOeejavwTk0wJMW61xzFIFzzK
s9xPImfKVv7/8dHWRM2OycffBwGdWl6JYsuZPuzV4aSN5ExCa3V9vGnoZzTGPdk3
sx/5lEm+LCHV+sdivZmryHI4TVS5K4zl6MaYpNH6fAVXRhLLQkxfjqPzUi/Q9wv0
W9ywjZOpCCyt5+Q+cTZ+0bFuWbd6mt4CYPUSZuNfiiyMwRLlB+eTQWfFuDMNuuct
DGCHBAjWay7BR6aCr/Q1ema3n06m9FBw6FrSL/P10wg1XBGTmDqAYIjG6zVoqKtD
wpQYfjxSlKzSqEDGYSSZK7ChcBpX+cD1gjN5aC2h/fw9oirZHyVSUn8lA9kpXWC8
g3oyD9prh7i/xAPhG8zfe5TFlrRfvKomAVt83sdlzlD/33eeK/YSsbEeevYmBOsj
KvLQueq8XCLnv+E4CXQBoEChzxkLoKmbhQnlUaHLV9Bmh6pQScln8qROGYK1phj4
PzQv4spzA3/7TeJtyKg2rBCPOzobISKPZPcTY7aPbATFFnq14T0hvnpwfv7HJdl8
i5BlRbk2258zod8HM3IXxdoOzgsml1GD0OST94ga2e/vu0ulQKJSnnfojEPizdo1
CoiszZhQHqkC8lXMhYMZEZBq6a6zy5LzuQYQlx4RMHWlCKa5+cHFaincLYIeonlE
CkVbi1uecYP2IKK8xOmpNHk2VWxgulDy44FFMsas9x2gi0xyTszyYM55Ct2ygXzR
VnaaHiDTEH05E4SxcK3Znbw3L3mshr1vxBO1Lz5MILBqqL2RFzV8vam7B1vSETzD
kF7Zb+kk//Ji9a17GTW4zMaxzYIZUHlSyE2C7mujBwHF+atxgHl7T/Q7OjrFu65C
cvKtmClMKbUtYLeIzE8hVrsY18rEsZH0cfaLj9e80C7rYY1j0JFej9+SvABcEptp
y+2qb7Q0uopEdcfPvvFNezvtPp0V4sdTIdnbtNMn1FCdZD2VBKEwUH4bg3zVGf2/
R2RAQonsYsqlIJHLTnUcvDpGS1Vq3bkrFqKIAcvEWczpbklVrGFx6pXqVq9DXIhN
MmxJ8vsnQl0TpUyw3LFQJMEDOrd3YxF8igZIXS58pNNihVXVuJWMeGMuK4J3sz9E
0nNcuJ9ros3f9opQ2rb2buFM4IN/Z+5jZXH76sea560w0opjNkU3HlV0CuRWr11z
HFxu7SpxGQJ86AXqtbL31Yv8fSXpdGgO+l/XCqKPpfsL7hGtlDnfuYtgu8Ek+QG1
0I/l/Mgk64tUSHCacR6iIIEDFlwTwo4b8zbdxG9YN74fhTfOYh0O1USCKdVcXktf
/0qUCRFQF6TrP9vJS2Elnh+ltzkNFjmLTKO1eg1b/qsphrcY8H/eTB84ZryGPeZh
dtloSzXDy7kFdVb0lORPHoOQuXgjtiB1rxQoJdrXaGlmHQfPtny5UOr9xmKMKQab
wWPk2V7O4tF6VMlKstoT5qOSox/XyHbUxjRdJW2LpuZ1coTAQsAChetBdMYkMyKi
Db4xu+Nblzr7g58mffwDPv7hblx2/CFEcf52rh13u1i02BHhppFPqJ+hif8uBgUq
w0wXDUTR6r6DwAAI2YyVlTqms/HN2lOrAfT/2SdYm/BfbOmYby0pVLHy1qXcowzZ
bxMDiOxrAi25YoPQItq+OHCojA6S/MlZIQUqmxCIs3o1DPidpTmGE5kLgqiDgsAj
i0wIns1qo6odNgFGXhqvdmcEuxsO2SjklOYsgCpKcE8XXMLyRI+/mj9v2So0lpqL
XA78uqKJm7rzK43SkCE9BPxieMSyp61xc1x2bJZX4jm8eOHwn1KSzwN+IkWbdlW+
S0bX91Zx3tBVs7oXmuOhgedIxiexPSgGoRvNKFckJFX9Pw8ZWvwXmEisV4NVcRXL
cB8Nk0UPerO0s++ugsLu4gfY6TYzSCDWU6/SQQUImgeOcRbu4YEKR8VigYP8D0oN
W0HLyGdGxdHpeO91ZnW1ZUpbY9XA/o1lk+FaMHcLEP9SEpuqWcxpkeJHpApl4J5s
XTFefTFjsRJaFKR1g1y28Xz+Gp5Bo8xwEnZ4iRL6ilRmuK7MOUEpVcDJ/q5dd+gF
WGd0VJ9nNCMfMP1+FrUgdLEUo42/C1y2ueIrBqz+JnKaAGGjBusV8ai2ckayRQka
x0cTzqesovrX4zaqwsKcxJm2/7UumeJavNh/9OpEWZHMj83zsxfYW5YbaQWGaYJ5
1DEU7cJyfywFxUswIs1vJmSm+zb2RprJnDGUObxU5IrBec6fERqKuk8AYN12CfDy
EEFeMVpdoxpUWM19NBYgWtBaK6uCgr5hclHj1bB8amJc/LY+uJyrnAvvAIB/gYkx
0hxlylVrm1XcIw9AMI6tGJZky5eAdI/HYRF9c4VzV4olXnOlhJfmvMKVdwWtwUa0
gPzaOZwKzEaI166LOgwyC+aeoUUts0poxTJSdkNv3Ax0fHk6oFhsdVRxcIVsSxUr
nFcdBB3TPjE4OjHqJcgfOnU+BD5MkYqvTYxj/8HrBfQMf1/S3QL6/eZfqKSfSEy+
gEH+c/Ip+B/LZNhZofKIQmdxZR8MIu916i0Ewbf5GCVgzbGqbOfAv8ImTs6WDWAl
cmnPvWJeaqGZSt6Kqrzu1jbssK77sQh6HLjo2TXPtWF6hkUPd7NmKpEv1JzJcQYT
7Lb5rV2R5TDl4I6PWlzA0FNA38noM6JdILbtkt9c0YJ+gTlTQ5sanEBV5+rRSLaW
Vkw6FFntvQ/vTwY/DYDrcKnD5VSwZqo70sctWrfnIpt613+73GMvmje7aYUXi/l6
HE0Ccnib4ld50rZ6Qf4DaTrVCCvhsSovcp6332B3JW8lRCazN8uad+i8IfbgvBJA
ytTq4qdvxJgeewVZIBMfZAr0F31VOrGYvsNaNzm+ymeSEtvsCttrjYwoBByheHmG
deSoTsbXPBdiLaUeyF7AMeMfDx4mAfpTvIDPXOGd8VMwgTk+oaKnL2lJmBOxO7RW
qE3Yv/s1snestJjsUe4IawsVvHbpWHcVj3iX6KxoWAt0ubIGFpvJVzxPyIVaxcNF
Wstc5p5amo4g8p8FhZ5W0uy9iVOTBrQug0mGn1meI++9LwygVNGs1ftHvkqJSq9e
RJiyvL6ol5FUg4ycCEI3lKR+nAjsBJxJdwYa+DFZb41r1nFrMFB98eoTwdECSYAV
jhkPVCOopo/43pQ+IzqOnJIrTTl6yog77prrQZ4G/nM1T4TbPbm9axWBMxeqprN0
3sC1KikYB/tqZFWHHKTUk7cYoBEheCL+/xkvOhWFag9RURRLoEEJ97P17nDi9jkB
9TOAVykotPq3eiw30bCDB1y8X8qwaEEHQ0V6VEcSrZy6b/ik3aQtZqtcPb/MA1Tk
KXuTPQydv5+DPyc4e32urqvMowImEtLaoIqLRKpY+zIsRa43GfY/k5jkCS9M6LPv
XJGhiN61Vn4j4Qcd/xwlkRlLl7w1Q6WksUf9ue75WSCTH9OMThmhVXw3mWhecHeN
HRBjwacA/B1DHT52Bi9nI2D11gVKd+0g3/wknsIu4EYT0lpJ/A/dxopMczWsR/TR
cDarkAKK1m7acvvji0qdU5WIqGcI1axU1oFhaNhuujlvbEbnRyCFHiMrDy6qDT5b
xlfuGWDX7MxCkBQjd/gRJIpsX0cb3xRv93HU4h8KLwJ1fy69sXvz+0emcu/+OHiO
rUew4Cs5EldF/GMLoOPvx++HieowtFtPcX0ux6zlznyhXVHNAJtsn1KNPr40MFl3
3MPhl7S4ijt323nppYaqhnI0axN6hH92L/n8EPdApqBYnHy9qIm/U9w1B9liaj/W
42fuU7/U4HCPvIV1qcyOI9aSdxMcff7XAu+ZW5tMAkbC9dcsGJGkgJAC4LcCUB0v
OmvQgpGlZb4Uhj6e2LTzyGn7P3TVUZ2Nd3yusr9nRjHZ3Ug5m97nYB+Y3Fs/gaJ7
c60d5L02yNLrfgHOwAUUMpHeRbmB2cjKEE2MYqsWnE//EQI5i+7h6auqvCJNrCE2
mzNDpB8LU1uhHE/X8OIS30+Lct0fyQVqiJ6LjodFgPSzL6nd3RhOKTQw+YgEkiO/
khK4j9y0tZ6zHWyr23EwNW20zN2WNWST4/KAu9EogVyOuO4pwdIodb5dIx3sPnWo
wOhVGZslvKE5fGntqElHvSelyh+JntW2Pm2qI1rPF0xBtZMU/u3AmL1MvE9K/3y8
AeHKgzLRHyfIzvx7gIOoik7PR5mltUQLprLqqdHiXYpahOoYsCIwQuQw+qbm2IOT
GIDv/IZ1J6fvhA6eJpsV6mODld7+VRvEdriExtu6s9DPsjsaOEs8S8cPOlShln01
WRFBQpZHZwoH4/0WBJDIQQSXh0TZBq+Y612op+NGA3Qztq33wGvwMigr5V+WMeQn
prgWZqfchox5pkMOyXJW5lMANMFZQyVB4izvz+Kc/AnWsOKskKR8/nELM+28eyub
5/o3tg5CWydMjJb6MgBdXyLJTpyCGaPYoVCwTMJY3x3guBc6G+o1Ihz2Y4z1xgYA
OcXwJaWvaB0BANqSPKohn4h9BpXKrPfu1pvp6cQlGHQD7/QeSxgdu+/y5OsLoKp9
b0/V5rLhCwSFF1ACZx61H/GuwceFZOjtpSXU2uQOPC4PczWYBzXHl2c5228hv6vj
a/RfJtbjBj729RtEltVXCWcKMcWlAGf7zNoloGKa34CHzdNuk1eu/YBcAP2vo2Ke
pFUKnmJLZZzrsCLh5k+tAFycTTRBMozTFj9ZYrKb7o4kmMiYxPrAMCwyT2C5p3h+
jOB5luA+960qjfH75a6i4La+8Yzb4DJZ2g9VznxS1tguFdUhQjHQxVF2VgfmM40c
+9oSmwDTJc0z502luFcJOLxVhq4mQ2dAV0l01coNFeHkGnoR7qiBEdL5Dk8PINdv
+KTg56O1JwXTPbqK0+QhKMJ7BgIxLqUOTdu1rtcyH/YN6mXsTmqYAEhsXzp530ix
5r1o4CaDciDs+LtPw4IzK5NFh2Kc5UJ3BqCnIliyrrPPuWMeoPLIdVlts7g/hAyv
`protect END_PROTECTED
