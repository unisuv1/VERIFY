`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tL96RoGgG2t3mYIGgGbQ8pQlrKrU1Ys1fa7LkgD+wTcwRCG1aXyARFLAVA7Ct8kJ
p3IEPaW9FFjJ1C48cxGT8usLhwbWWzMrw3+waRcH08izb54gSrx3Tk5cD/H1Yib3
cL1dDt2D21XtxWHE/4h6BymQPqR4S+N9DD3AFJqX1ScR2XHnQkYCfhPivXG4Dt3C
v5e0VoBjJYSMPnsLfTRru2q9XK+x/gq7sodB8iajsuDRDjFhc+OOeDAIYvqY/qyO
qMV4fIqCG9z1OZi+sqzS/WJFZisZZau2sSyiKG5KbRUHP7h5a72lmAG3M1P4Sdwh
U+s2ca7AnslY8RpKJ18EOHKCZkmCYmJ/7xLSf8OonVX+VdBMnEGNPkVs4fZJnsmQ
U2xkkLFIFLEjH3nZUUglRBE8Yek8FxMR0Bu+stRtMWAQM8ZxOecEoU0BPYftqdxK
99ix+d6k/cPUFdhSMYNdDg==
`protect END_PROTECTED
