`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
A6YH2/4UaiTbEVrdqey0s+PY+MXnN8oQp4vre/ZslUs090ovx9mrDvRuOf33w103
aeVOrOn2wKviLjidZHEPwFKDuDyLkDTcaKtvh3aNIJek4f8f0chN4KzkFZ95PHNw
a866DS6Rs7pRTf2/A0c6ESsOcUXc7Ar0FGOSjsgluwpToB7g4appJWi1a3STtDAj
pOVRFHmQgSxQ2keXxiNKCkqcg0MK+b03z41qNIlV55veBhKNVszY6zckJ01beNjv
xRkF49lqy/NUOdzf6mgKEFyURlZ0JTIA/M+NAENgQzJTxLQxUIX6SczPLtQBrw8Q
OZGMyTArR3vEXJGHw7UgFN87ry9XHbgO4xasVRFkS+JT4gaaIdpdYAt/5h/txJlO
YpMn1MDMq7RpYmCEugXyLUy4Gt1/+vTtDLjgva5SHeA462lf59m9jIOR3h1bFCzH
ubG0F9vsk0D73cvp5wnFZl+2kWvM+PIXD4iuXf0ccZ7xk6Iegp/ysGTIGLl9Q8hL
GxEYxyhzIoyRlSqebiYtBd/7ML5Xble/B599dbsJ2To2OjDuMFAcMvgbDm3f6t1T
9O+k3eqwDfWZ1zHdNoc2kxsVnYGrcFMhtsCTHid0oi0QeG2L/R8fdhZLdSY/WZCW
6OV92WH1MmccFqBrxcRpjIEIxY5rSizN4CbltSC7GE90vZ0pelhVOya5PGDMGzN5
MEx0jsvsRa240jZsuehyY97E6bEOy7/z2I7vXByfGwJCSIg8xPo4oVHY6KtwsV9y
Vtt8CxPdlTGYj10yTooV3MPQnu0lTKGDbiYJtighVMzrgNsIB6Rfozgb50Y/SZNU
kw9SYu1KuvKHW+285QFc2ld9n5zvHf+OOgvn4z/W2omJG9+wmZFr7mZcTUe/dWwi
3UXVl7peeKQ+jfhbSm7XBf2fUuDYmRL4WgluVclVEs0RDYY/hc5wolKPniDvxSzK
wX1xIT8Sy4U0yxHxmcoXXRBO+3Jx4IWVGJEK0miXUXxondDuAmG+Ebo75npSzqXE
F7gYlFsEel+NXyqYLyrIXBWRx+ziMr38fZGmGdIEXXZrVXFrfiCsXXORuGpK5+i7
sVu8aDr6tgX6aj+WD2Kr1LnbwLQw74J4XAhVBLIjJqbbQKvIdTKlg/J5zF071vlj
9hAb5QF2BBt/AOsvURVBJadA2fCDE3YMEgvqblHlC6Za0dxN7lk4UytaFZpLVMFL
/K6/XtqRD95Sy4YIRemcNfTqsDF0GEoSL5a3Z/ecYylXdhlNuP58pRlOEPAUS3Dg
U5B13awzfpRiAaj/Auh7vTVATs38Uv3njYzBl4uaq+AhROHTEJtrq8L+45SYQu42
S/NX4A234eDjU2JMpVIS9JplTHrfqCVdwMzJNgGDVKRtPOfPRmzXG+rnm/5Y9XsL
RnGCtFNevOMbcNFj0gJSWSbRQ2A8VHGPsgJln64Qar/aGrRg36STQPCdQHn8KJNO
lfGiQPmj5xqA6BF5hWOVECCBXz0kUuqsQiSOI/Vo4MYh5sx5mxmbQpXcmyCdLvQE
FVCYVFlwaodeKuKB1XVihVPaViv/Vflxr25e8NmXK2o10k+NhD251RdUs5V8Ul8A
wrCHVt4z+ROQMKi1fmPTGF55rbZPbaDzc67q1rxXQ/W6VDZ1WlmcPdIvxtsXnlnz
uUvVO5W+EnHy57W2NDFXpjgGFBsVlWq+HWIKae3k5Juo+cFl2w4/zS99TOyZSm3P
fRiDXBOcgPSJ81tBJm1rsDdKiWXkd8qA64KdKskXkah8fp2f/wxWMeHbhSosfvk1
nKsY1eHi5i28Q4h6Effgq9VuqgoQwvfPlllIzKxyzmTcTM3BwgyCs6TN3g5Jf7Mw
UiLnwFlDGkpsb3vCPkepgPu9RWWDZIGEpI0dl7ITZSGb9T+19lfw9IYLDILMvduZ
qUm71Iu5Z9okCWyF1zpYTHHgy3fu0VO32C0V49L/DU8lVhhSNhVXJaAzNejBtepF
lMddcschOOzR0IIcAG6NVV1W2RD4PRrndZ9Jh9XxC7ffk2uzJm4VgvCmWCUG0Oga
TDXjTy48EpQLrcUL8wKhoVmt0jVAn72zYnDOIl/JpQIMMn4VaqJh8t7giNY7xLQk
XeDBFcbeE9FZi1rzXJpk2P86q4vRd3l8R9b/t1tnym42QCfAXtmL3laxmpSArQdl
bSg5trJd+kDgTUkQhc+AefuC9OgLjWJ9eSRCG9N+vUAcHTE9uSKrJReLj/PJJQx7
j0afxgsxk7Tay4YJhDvrS/y5/+1wpgBMiv5CWMgLKWsxI5Zv13q9kl47+0FFYDVq
Q+DKoZwL5iLDXrPf0wZy2OD9WVxjNFHZ3DgGJcb56OfKuK0Y/OUP1VNkxEdNtN/h
9Vs/0LdWRWTo4YlbnaMwua275CBFmCzdtXTOBXieqFGGHQ4ttdDIFH47XoH4TM4M
Xaf5XssyjoKH6ZlRvzpAjsjZiP4ivzyHQ6C0N1/cVCkrGjgW9xgwf9d5Dep9UW7N
fx9CcXJu4qJbsc3jyswZ1zziWpxH93ALAjFZgb0CtsRfu5Lt0C30ABYeKkh3GTmB
VDtxacwKPY1D6osh03QNW8nzFI764rvVThaK9ts3iEL3rg9veaMN1yHk67AH4Kqi
jx5+DFA9TBg8PfkQ8HqXu+m4NxIYWQ1AOFZE53xGDMHIm6A8MTLtiwrLig8aTJBZ
di26d5qDvvqan/ME3lQQTRnTrToXRHJfHhBLx2Vx/lvM+BUXnFtOIOPB3nmuwLlN
uAHCaRm6O5g6jEUqdcqbsOl/HmAKWjeeFQXok5CQAe+/VbSeQ79a7YSPn8tpGRbq
kj7OZiuXzzmKvVlWCrIbjdJtIvVrQ5MrD/6ROD0zgG0cZQIi5jp3zNdN7KXk6jd+
pMC+h4l6srAxVo+uxTHcGIepLFKx9tvY8DFHaZxPl858ItAkPiaBRifHvoYUnsQ8
sQPySzo5680LqZXdQq8o2Q4A/e27rVUr9iBKevgyK2EMSfPnuicZ2/iXzGzZK4jg
7KrMBhAefuH2wLw9iHKTtf6ESgRCI3p/PgFMiUyrYlTNHY2i7PsT2Jo8SMzHl/gO
KrQ5s2KhG5OmYg+wIZvcTiCVzUOC1dvs8OteguJlzUZVsBTE9xEBrdkRmMqq7+ZG
cOchENY4WzyDrLAjTslNzbcVS7OD/fswfARU4a0L0nirR2/vF9qccoSHYjxOkNLO
l9uIAkxGMfgNwMJ0QzEG+HxPHmVx0Hc5jgxaPis+LF9PYmH3fy76A1wxPUJywmMl
rBQ/peVXxz06hpE24R58OzCGz6tL61AoxMml1YqLNSRMaj9OYw+BjhIn2Y5me1RG
y5OxeZWUu5bk7yK8jlBmV5lLVLTWh9uEG8ZcVX2rpdbvvtCfHiC8FtRdUs9tTe7n
dBKYMojRMezZLwftyHOdTWKGFOTlChqyP0dvxj5mQl5ZWAbLo2U34qjXnAJrXLKI
rDgjxiaZSf96a4Pwr4R7rxxoLJZ51R6X7l/PDbyD5e//eh73HwGkmMovii36GBck
IiFt3wDvrL+OQrNrm9Vwu3hJSsczFvxi0weNZAeoJIIc0ohI2nPU4uspaMVcg1j/
giDR+Xjhym0P3ubc79RuPU7S2LqEJMclTXLTZ29paoAJFudSMkVQ2FxXdKuM3khY
FAs7NyU2iaXw8YZp+eA0wRdzpyfPLhoBTPSE+ge/XRrPXJUaE3Tk0apRaLKQbgxL
7OWOSktV9DyhrSm/JfOS9EzvKg6mONUlZj6jZehgI0DCyJlMKj9A6v5OwI7XUcZ1
xcE4AsXGqDoMJ1HhP4/Ljlg+g6UhsBWhVonHURGOuIGJfDU1IF5ekT3sgxe21/Z6
4YFlYRgTWtgjtqnRs5XTmqzup917RHXKzNIKJ7VpJ+MT0JZCzMKvpDtpRQ21evle
6WvVjMCtWZ2UZIG1Szg9QUjxju22fZlNineYe7cta61DkVrcGoVjRs8vOVja9WNN
xas/zuorwB6SDUEoMGqQNadaBM+5wY3Nfqs3tNWIZI+SDi/7aFCRwjkRVsvjjFSh
nu2/VsMVfRfF+3Drq+kTV6OC7WUjY1s4dgYXM9RInL0dZDAtuSpC+gBwq6sXFsgX
ohgYLQoOHL3jfewRSBh1a+ew/3cXsnGReNldiOmwT5NjacO1Q21AfIXJtGKDut8z
mXhmggi5oOxEU5iFm3StZcR457FSVWXK7mtRwkt7fdE4g9otw4nL4+J4cSfLSBC0
QICpdorwC7IB6M/YgcKVkW0QjAGASLy3OQhpQXh9gGz399VEMBMYTYLC0l73Ad3o
JOzb9AcTUOr4tfCo28jtjjoIK4TqfEgEBGFeCj8w3yPNp/gN71NefrkiCsLFy2jF
QFXLCljW+OZqW7q9qXwGRtbASjyMQm8vv5Eb0xCvut/FiqAbLJn1mo/QnTyn17za
Cu0SJMYQ7Tgxv4hCnsfmZ4jqgJluYn0s5xDU+s7nQqhxIC2YsSt/11k2MT+Cqqai
9/6AjSCHo7KLiNlPxBWh5GLrzku1l2aNqprg7KYKUVkq+eeDojNgj8Rj0lB2v3n+
5R8w+MceG7vHDLhIfOG4z3XBW2tbQzfUDb3etF3WtyGTnlLXGl54cIxXrhIX039A
LBkcZRqPwAGRWcJIaaDI9CNVMmRk6XvHwNbXIn5K8kFQFRZ1JywHbuhkNto0OK1y
d/6wB7UrIgGoQ5XuY5dE40bUUXIS9f1b4e8U7/2OMdiWF7wPcbuF+S/Ei7yqaPAm
GgwumpnE1uX+hxGkb1UbeTotRiNecg8af2J/2bfP9Z5qUniSif0rNd0xyKKCdrts
KYOhxcLuHo/wrwtMHNmP97uaoDNoDnBu96Ntl3GjjjR6rSZujmDKvuYvWrX0gPJS
5EQrVkqyt/pMVD1mKmIfKOQ59njTjTZH3BuvADX2H7BruTyp11Hp5DOoXbV859gT
9PCyi+LqIVzsVazj/sPOLQYb0qoGSIAZve0Htmlal4goHtmhIAoqOMnWLTw2fERo
/Sco8YwXhcPqdBUR68lslNpNBQObYex4uWnTBMaSAuQM3prKaI2rb4km2lFn6QkL
ZO2PBqztm2FzFc7e74gSFa67Y34+3U73PAQ2sR1jQzRyG0cjXHOX8CaYMRubEvrK
4vOOND0+rgDUGeUPvxE9nmZ0m6q/cnnDDvmuYattLiYIr5+V10i8ExeROTaDUrMz
tkHzNcQaYlfBkKxWsfNLcMD3G5yXCFG6ctElAncbpxiktAZzDrXi2lp9aTI3KUzc
X3og1hBntr3w+3K+k8VNmomdszQfguQkYBRVKnxXGl5foEmmEp/JPTs5/eAit9qC
LFjrMyRahc6jM1vxme/t06tMS8ETgXBtFPu7cWzRacqaoKw7p0gukxqKvIFoTQAt
bqOSNZf+JLieRSVh8/a4HuZvrnOwHQHEFV9IgyQMzSmvJo6EtOlAcYTH9QkDV9Dj
aVNmqlZ3t6uv2H7pMEOQSNnHwZCZPxN7oCbtrJZBF8wt6onrYfZ4GMGaYRutZjcA
ty40jIHr0wiL1seRNsP9/1p8UrpuK3IoOs5lcM6mo/s0Sz+dUtpu+q598+DJFl2L
uifEdi7QIxPYJazTEdgUrat/RLd1h6FNLZIuErZCnCju5t0jo3y1SYXXfNcwpjgy
Pop1OLVxTOKZPzG8gnHVxFGBxJCudyIoMXp3FYnxTurQbupaSNq1bS5WR5UJlEsk
2jFrgBrfl61FJ8sBsgwOc5fFGkh2V40viH94+OK7FCYFAVG9Psehr+Lnpek3esMq
r/NXRU2pqutyFiJNNhmg4Z5xkpIVE9GvEanUV2L/d67RrFhFEZVpSN2GR9b3jNQ6
XahFwR+6qfcJP3Y906HEVWn3hsVHYmyS6V+YwTu8YxVBxNQcKKddDAzNKsu4TqmC
G5aVRUbbXeT+wR8IonYhqLP72GnydkEZMrZL9vgejLumFHtJbEFjFetmj6Ul2p2n
mlz5vmrx3Rde3CwrA89c44n+v3XLY6QtbSHL7XhZ/2Sj+R/bBYXJizRP1zGNp27B
+8YpSRjqMTdvo9ZVk+2XuDl/aolid+6FImpvtC8fCb+SZIGI0LZnGOYT2voJcm0k
Lkf7BYZClFffuBQhERfkoxT09NUaQtzrwiXKIZEWm7VKOwkaQkwRlY3eRC0pfGVy
rXUrsilh6LkPAUYnkjiuP/N9FJcNPcQFFBYEYRqpmHgDMSDK7yef3lB06pisy0fb
DeJTsksCY61FFGoTD3yEXEdsBJ5yFdz7hdGYLkxsCBlTczc+kykY5RQXJGfhfdSb
4vaR9Vve3HkIosUrXXOtGzg29E6EzbHICmGQPKouUJlnv7UDDX2r3Ukww5Fzz7TW
LA4wzo0aA0Hu2UyPsM+DDYhQJO0CvCw8Ev0ra1dm+ypH4BEnfsiAylAxXMJvvFbu
1V9/Ny7vQHeDakmFoaa/HputmpDqi7braQAlvWOgl1pkRxFHLJr4Ct5PN7cKZUaT
0px3pe6G7kb7o0r5Vlu1tDqgQubVkbMe4DhAYsdCxB9fr0xh4ZnUNWZUlvJ7p63K
0ZNMs0fQBgl1FbLM2Gu0W76LuU6FJE+mJ+5g0r0NSCkM7hIMZkPtgvYc5giwdKF4
S8CIWTCYfI8N07ItGEE0XFqdh6pjpEQz7y4Swyl+JbMOEjWgppm5g2CJgr9y7NZh
pdOqF42fVOxOci17h/oETrUoFtkMemZ5uk6U0sIU9Skrkq/nU3Kfx9tq5X0vbEzV
yOqi5ZxUJp6yXzGKZopVCsL7jgIibC4Q+IeQQUlznTedTceGfBYCsinw8ywurblN
mlRaqHqAWbSNbrZffYsVNVp/cTgfTcOonylODhX6IH5qZuHpmVQBuX5y6AzyrPtV
5U74EDisHF97z1nKxapgxz2G7zdeyLoXJGDTpmWutxFv9IShfVOK99RPjtMcN0b2
LWVOOkiwCr+sbgjoQpC8gdbSlMiv5mI7CfgpgYaPD5kJVAV5A224JhPyZTeLEEue
uHXOpMKKYuKudV7h4lujAcdQkfabmOwy0YmTBIf+S1spWGzUxzOpA88rXJz1WDUC
6P953rSBe6+82DGziJ0Ym2frzhUwQtUZcVVICysU0XuHX8zxOmjzZthXceETIdRL
La0mPOkfyjBpj0jO7qoRUZSfpppLakaADhUzxxpjp7GW4cY9y6fcdpS2+VWGfVj+
LDZgKn/ZADkZw1xgEyd1/sS9Qa2kJfd05BVhnKOjHlPsVM7rmMAsDimn1Tywsihp
zzc1XEPvrnJcdQKhvF0X3AHAV3qCWqRfEZKWdQWc4UtRC/QtaGPsn4+tWQ4Q6CM3
PsEblQAklTSy7Cx0NgQxC/yIBWZDixRuibCqvsU636JTREWHcSwCm8VQHiWEU+lj
thi+x2pRj83Ki02gfcIgiC81HPEItScFR9FDs+VpsiKU9WRLMenB8eFNLspsaTDa
DtxJUKJqbK6rk8o3X0aFEEBi+olFU+ZSa37df68s7BbfbZYbbNxfrN9JBzfcfTzK
iKjmE/RSEfC1bYOGjt1xI+xayK5wvTAF7jFtxHBUdJMwO+6Wl+FSSJJH6Q75GW3f
UOnbtnGggReWclhFJGAfiZjBM7jNl0OfyzZyElSVbA9TplJpO0FCoUb3hYz/xAxd
Ff22u3BxTAfy2ril5ETdCWKWuHVyQLCVeFr3doi/zuldDI5uSs2S0rV/e7VfDPhD
grl6FHFhvn6wgG8UiEL5G98WrY8xEIObs1L/eUO40Bi/2SU30ESpnF42ZDfkl0l1
9nCPzNhxUK7DupImwkkqWxy2cZ3h2zQYEy6PYdTQ7zqdABmva7DOSDL36HAMu5H4
EqgGPUi1goKZ2g47hAl1h4s4dVG2OVa1vsXa0cmoDrb6MICUhXT/ZYIjAgbIP5oT
OUsWw/alvNillXGkDQ4pezoW1DOjT+o9XN4OML2GzZy9z12ckhif822AbQGHWT9f
gfWsTlVQ3LVliaUiW4t/5zbe92kTy8iAnw6M72W5dBRyDEfC/qLPC2irWWECT9vQ
FYswwuoL+QS4Znvp1y4uW2VqVvHeAglr+VuJY4nBpIOVFBZtWa3y45OeD6hACcHP
IM6od7DnRN8i9DnfvS1sHUtkzWopdm591/IndiRT/kVMFnKzNHcdUJWpS+UbfhOy
sOLu/9HsAuEwCEvOhHAByQRH8mNnjf0YSVmxXP3788iKBtqLn4ULaUefSYrTUTE2
SmQJuVZwK1LOTfZymIzffF2lgfPhailt6RRFpmlj9NyqYPyxzNTbcMYVce3mTn/f
xpNdVK8ToaoIbbfjEeK1Az/Ch8Woe2tmukcsh49MpxSTSsxsnP5uHEJYM+OUo2aL
5CZkgt2Ak7iOY9M2MkfhM//lQREOX3AOju/i4+WylH7dkQ51RLT/3qr1jOQyb7no
C253QqziOa8irOlCNr7Zzj5h2OAYM0Cks1ORBFmWp7e38ekSwpU3H1gnnHYH8D0h
bA+W1kFQeNlM6Z5OX9oduECm5bgbI2BCwVUwlmVkLJDYuJVNACUjG9J32p+Qya54
FJSo6qRJ/yxsDQHIBrKOumt/RXoXuBO4tSv5dYxoP/YOwOWIG3t4gWn/mXU/FA4Q
k/O2lqNRT9X3E9j8+9Aphb4hmlcDcCvAdPvCQtKaC+3aTxm16QzHEC6Tal1hnO2J
nu0YPBIm+wobT7SNQLiz2CBbLbLtGP4XmoTAxXQX+pX0T3aMTirYMTtPOapEv9lC
B0SRpNIu4L/tfrqjlDYFZ65mulcoB2/1eTCqclVR4wXGcCtnGKSocfulZwT6Hlhj
UkE+MIOEw6s3uFUI4nx2bgNm1UvRncVhtHtnmJUEzib5I/MrmApdQSJfVjr4k5FE
6ROec1DmZBUEZHMMkpzBKzBbVl/IguALhcYOwyCdHWPsC1m3E7QOCvHRIae9rxw4
yFxCg2ipL4y2SD/4G6jXiHG3yIPBc5Hy8Y4y61gDoONbyweOLHEN11ohYiacFVKu
MavJpz6wo+twsb65S7zHIKpPBiAYrGjFQufvHgIJ61D6obIbaDlFLpy0xMotKL7N
nTJE9UEl66rPIVzwwvQE7k9nAOJcozoUx+15/RNxzNaCHoNZ7sS1eoReWLHlibdO
PFmnC/9hVm0hZiJJ7TALVUfCWQtDFLlm9UjdeozQSyK0DcCzqxHFrINqEERRWXqA
CoVQRg5LcbWCb0oTMal3Z0k/H71vRNwuNmSilT8t1871O+lckb5sLChdB4cIvLje
wyjzgg6Z3FJTp1RMsf6FfwVsDnDdzAKPwijMWenExF8Et+wPx6unBIHen7ZJUGTa
SsnbhGht9PWuBYruVsmqFze2ww9GVHoINLUDOOCUtnlbVQrZbr4aZBeEGZ/pcQjJ
ecwwcrsvFLwhd1ireZLaawYmi8DPRMFFmUUplBqxc9RBrRS2pZ0dzjeZefDNZjbw
RjXxX9IuJIIKhOrRyjvv5GWZZgYjW+xjXmHqxw216gRJEkN9qVQZdjTePCzkufWX
xknkzfp5a0vaDWNx53+v3ixFEh4N1CdQFLweOcmGRxY=
`protect END_PROTECTED
