`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IKAc1n7iee8HTD3UgJBl2QInEwX3zE7a25xfjs3uUnQI/PIAzKLshbEKhb3pcDL5
/nXGl6ioSydoWMAwWt8Air/XZF/LVuHjSCGxfgMpYB7QbQ5cWDZDAnO/vGnuiHUB
WzxwYcIwMYFpM4K2rYjCnWHvUi7p+ARV5nMuhwbldl+C1eXj4sq79jufkoZqfzGE
213RC60pnFsF61tRpPzFRLwhRQIAVbLvOc9kuZjT08xp+J7tDRSyQOibUg7OCfNL
YMNOdxMjzxEFUeKBvB6/eH54Fo8oZvrfih3jaR3udGWINep0ka26iYLxPaYWk9uy
rICBItoD97d+K1d55mUy/ivdS3jp9GA9oyJCQ2k33eCJX6/KJrjPLf1yY17iBIDz
/+/+mRm+2q0y+QTomNUakrsdjB9LVK2aettDS56uKWX/VyG0D7iD+1CTblbT/GaA
k+St/Y/mcWKu1YFnis6vEgz4oYhnziPbOWWudtnXWNI437d/IAIqMRQUhB6xkLRB
IjavPmFs9sM0Dq0X0U0P+N8Ej1Vi6iwH98k+5V0aQrc1c0AGrEG5ds0SKYpbVOy3
TNXC756wdvT760X3lL/Q4bYpih5AOo3zkYo63qYb8akl5e0WXQksREDWV6Bd7aT8
bPSgH89DU9vhqpz7zl4boCQKQ6xFnGtZdlZfrtf8hsVWcyjfJIus78wEy2qpedez
mxh7CUbB4dNm+csZM6kyH6sqawsD4LLqe3hyRIa6QHtvGsf3soGB3YCiCo6wYMq+
oUuoGWzOobaIaXxmm8cM+Ffv+FYUeG0iPfRKwMEfwEKazGXWkhWZVhf7MEj3NjXB
lZYS9mYogqfnHtWakYMCbjS6Ig9U39NNTRyemJnkO5huqXFvKlYu9jB6d5BNH7CY
EFbi32mZPWdSpVctv3zN5/5CjgMPJ743rTw9vIWo7/0BNcbm1TSBM/aOPG3oHa7H
uIMROAFCrWoL5ED/AOFEBDYKgBWHPTYHQy3QwEBOyMm+XV1+jvT25Um38SAtD2Ir
JIioL70Kl7KeJ52r1hMzToLsPCB6tGLZKx/9Se1MsbNMG0kfIuFmlfjkg3sfXfDs
v6jY5iNPJmoHfxX+K8MVqejAOCVEDu3M18UFLu8Wq2qibCZZ3DIJRB22YwyutGcO
1kUneKyiD+ZmeozseCsgyQ0PdZBVlpTr8vXiRKNqQeesIfZ6yzuQ/bz4dSKXgzlt
Bxa+/6S2DUODgI0DJor5qW82oWvj4bMBe/Nm+wgnXK/uXz5PVb3YirYSLWYJDlNK
KMiUNctK5A8rDV+L1UQY8PATn6lIZK6shtUTs5xPGTynezKiR+GFrb1HlnLAxtsS
Qv7VjwTFHjCC0NhqVl4lXJj5aLX+jfyiuniYwff13WmuZjLAeA1eoGIuVhjWLC0C
U8ZT4PKS4aMqpIlC2t9WIdhzGjbSagkk38AbPbTUAEZuZGYOpUuMck1lN4rf/RQj
qDGoj91wivp1Y6sqV5KvHtpNJ/KhBGI5Us6ojdvuNSOVs0UwZCmNp4NVuqZNe5sw
L+e4Ro3lZ4GSTep8K88AQSFpOQCH9HnIE+kAvonbdjVTxFwNWK9PjRvgq6B3ViK/
+xnLQndnEVkc8UueN2hdtCC9Q17TMcea/q8byqZVuFYB2eIgPjGpxuE9ggRmCpi/
trrs9X/pCtCk6ASu34REMvf3Vg9CEqZd9LyEmzP6PVY0jHb7eUIy7gDwQ8EQGa/Y
DXma/kZj57cIyH3MW4W5HPORWT9sJE6oIP8QCVaRC7TBnNX6X5eEbzSG3DgaDr2A
utwC53ULBZrNQ+70PQZhysn5T9SRpQbd+PIfCTwQLSy6jO8zN2h5BBGY2SDgeZ3u
/Q7d9JwJElHxgJwKp7g77MBVCspuSLkXgvtE1k2nSVC1pKu1qIcgcUoDEscwqLt9
dgyChjYhxV2b76XiMxlbVeGyS3Q+D/NRZJZWnmMK61bt7LsYDrQ1huoFlZqHSA8u
Nhh9l7HC6yX7Qvs9lyxfj1I1xrPmFDQl/GHzhj7U/TYugi/qwoNzEM4JzvdjKuns
c0dkjuMPW50QGxCaqjLEVcQAH/rgPHICG6I7nksCLF2kxwDyYChu1AdrUCM9aIX0
XxPSn3lUYXWzqvEoaHO7b3Z4+aHPOZ9duUq5cX03GrcdFfLFrnUamJ1+4nLDqInx
mBodnU6imRZ3/UQFAdl8y928CWedj1nMO0fT0t9k9FZGgk4dzgcLdgBNV763vk2/
+VQZR/VygVWF1s203ukHMKLClGHKQNt6nttXoeFOPK3cMNhcCiwen3SLT/mlY5MK
P+cUtxmRa/iQyso04bPo2bYFFm9l3lPy4sVch85E7OCD6c6sRNTw8+gh6gQGO5kT
1y9HktsBMDjwsZVjeql5HB+Nhdbo/dadzPCGOscIjjVCTrhOyVz9wK+7y+50OH7+
/lBEoBtizZldxNtbSwT6X7L5XwM+brl6c4sDTfGbEK2xx26w1R6Og5gcs0mqhVGz
1ffJj+aoQY672i1PN6iUa4J5SLABlhLQx7qw0pAUEXTGO5raAPoxnRFYEPrJadhj
LKHDod7PRqInVO1N54KgiSIdOBpeOGqR50jc90PHI1OKgTEPuDgpc5X2pnD4VVn2
XD73YmjStKvJoCDfffA/LCmK0d13NwLMONkifnn4BuP5s9LPH/QTacAE+eXL1g0B
nqJG9eD2s6bff9kAtlMcHyl/z3dazImyYesVRKBMI+fwVTXZ+gqHY9jUTOKzJ0Z1
/YZxsnj0C0dw302UsQFwIFlBoHbuqhPyPzLjWGewNWcyf3aeZdySxIHyhf14/UWf
lbPZcnYhdYVQtzF/FfF20wAu5Fj7eSrLn9I85I+835IorHxzR4Xob2p70W8eszoB
gwCF2d7d8Rt15UjPG3a74GwYjoILl4S2mE5JPiQnuwOt4PFCeTBy5ojAJgrnHVg9
lmu8EgxS2tyEkbaiFeiGv4q02zaWBY46V2vYhv9TAo3B84vDFYa4QbXSVdgu3HGl
TJJeBgo1tfMA1OzMwb6He30VvvRdBxe5fxx4TV76KWm+tckDtNBQgMwxAJb1cCyW
3dZx0CizSNBGhWW4Qou+6h7m/xWM11YlnE8zLAdUrUW+SxI5SWpGZPI3uo3qGJDK
Y29LSgjrxbmuln5ZlszyUjQUeXlrULvzJZ2ev92cJoqdodSrJydSUMwz7WOlby34
SkfbOdp6kYnC7SEEbp8I/rVGoTd/0sVoMZFIpCblt/9BVajAARnRBZWWhbTp3TPS
xYCeZpuWlbObsGe3bs+yVvihgiNp85n0baSWAVqMqoW5ZAP9Id68EU5pZzkem1An
BobjSZYKaGWjxi9lwi0XCNJJm6+Kz6s+7XMHFLwX0FVXrwCNK61XWmo4JA/zAZus
nolQjLTIrDgEb+1m3zku3H5laJzULBT9mTE7BrCNIsSpGdkpKUKMMo3YQ7y4sfCV
Zsm+RtH36pVWkd7Y0YeKnJMw6oFepi1B1ZOJ1n3KgQYFeHf+JTwdHy6Yx982aKgm
pCtc+ZohoKvPJFvikKaA0/uaJxejtVWIYrAnpFdEtLo85wHACCfYPsBXZxWkQyLf
Unskrhs8ZXvZwNEmMuvHGlOC13Y+hnLJztWZKBxACT99zLGV7gxZwRJzo30M4sIo
7Abd9fs5k9wbjn25Feoiehq4AoxfnhqXbUcH3pNysHVZ97Kg6N/HbTj/mEN3YQc3
uPYBu0lPuVSGq5aQ/G1v8g==
`protect END_PROTECTED
