`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
50pGr7FRS+vlMShUPXWPqdhMNeubxBOVsdcqMHzkcAz8IXz/4IM7MBbu2ObLW7AX
uG5YxywF5sTlby8BORRJjwofTSmdFqv0mHwXe3swvIHlMNo0HmbxMzBwqML1mkiG
u0uQKSGXl62UKmaJhoHmpktQGnvIopMGoOGfo+62gi41+BuPS2aAzb7pzqTvmGPu
LP3dkzmdFZkhwqwDWzePeZpOGKwA1EOXtWC+OGq5mbU3f9EVmV1r93jjmr3HJYAN
2pWPv5oD0s+OBlZTGX1xgKDGp6LW2H8qtq6XnatC4poWDf2K8q95LFtG2X441771
dimCoq6uY9d+UuasW/DDvxWdP9Fl9P1u0sGZgOdiYjUFbOKswaSVmUypA+Ivx3E5
no1rnyZcHTgAUutHTDKk5i9gbBxRE2DG7W9hiI0CSsRTVlBAXB61l1k/JzCtYPAB
ihOGBSyuTI1ET5+dM1l9PNsoJR8HoNMzpBR74W21zeIaABOrt4QQ4L/rwuTUo8Ue
cOESbVSDN1tZA6lCAqelGrxc9mB4Zfbri2TrBW+MD4IW/ESkcBA9pgJUl14xckaA
J4J0L19TFn8sALXH/EwidFaes0h6xffUj23KwY/EkVXUIxAeFo68JaUlLGhIDDwU
n/WdrKFCDJEuuCrwLX/vQRs8kHFgQGuHhlJwoFy6/3TT8fcVClm4mdJ4KWYGFaW9
Sf7BhWV6+uRbc9MErP0TsQ+jZhQeeW9CIH8Q6YvID5Hjun8nnjApTRUq2fwqV2Z9
5F+wJdc/Kc7JexaJqvNO5tlu35zm4FRszCiVXWdXJbEr9NvLRoIFM7oJeQKBWbkG
`protect END_PROTECTED
