LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;

ENTITY VIRTUAL_DY IS
	PORT
	(
		nRST				: in std_logic;
		clk					: in std_logic;
	
		gen_en_sensor		: in std_logic;		---�������ʹ���ź�
		default_out			: in std_logic;		---�����������
		
		sensor_cycle		: in std_logic_vector(63 downto 0);	---����������ڣ���λ�����굥λ��
		sensor_valid_time	: in std_logic_vector(31 downto 0);	---���������Ч��ƽ����ʱ�䣨ʱ������
		SPR_XRawCoor		: in std_logic_vector(63 downto 0);	---ʵʱ����		
			
		gen_dy_out				: out std_logic		---��������ź�
	);
END ENTITY;
	
ARCHITECTURE BEHV OF VIRTUAL_DY	IS

signal gen_dy_cnt			: std_logic_vector(31 downto 0);  		
signal Pre_SPR_XRawCoor		: std_logic_vector(63 downto 0) := (others => '0');	
signal trigger				: std_logic := '0';

signal SPR_XRawCoor_r1		: std_logic_vector(63 downto 0);
signal SPR_XRawCoor_r2		: std_logic_vector(63 downto 0);

signal gen_dy				: std_logic;
signal gen_dy_r1			: std_logic;
signal gen_dy_r2			: std_logic;

signal sensor_cycle_cut		:std_logic_vector(31 downto 0);
	
BEGIN
	
	sensor_cycle_cut <= sensor_cycle(31 downto 0);
	
	process(clk) begin 
		if(clk'event and clk = '1') then 
			SPR_XRawCoor_r1 <= SPR_XRawCoor;
			SPR_XRawCoor_r2 <= SPR_XRawCoor_r1;			
		end if;		
	end process;
	
	process(clk) begin 
		if(clk'event and clk = '1') then 
			gen_dy_r1 <= gen_dy;
			gen_dy_r2 <= gen_dy_r1;			
		end if;		
	end process;
	gen_dy_out <= gen_dy_r2;
	
	
	process(clk, gen_en_sensor, nRST,default_out)
	begin
		if(clk'event and clk = '1') then
			if(nRST = '0') then
				gen_dy_cnt			<= (others => '0');
				Pre_SPR_XRawCoor 	<= SPR_XRawCoor_r2;
				trigger				<= '0';
				gen_dy 				<= default_out;	
			else	
				if(SPR_XRawCoor_r2 - Pre_SPR_XRawCoor >= sensor_cycle_cut) then
					Pre_SPR_XRawCoor	<= SPR_XRawCoor_r2;
					trigger				<=  '1';
				end if;
			
				if(trigger = '1') then
					if(gen_dy_cnt < sensor_valid_time) then		-- edge is 100us 
						gen_dy_cnt 	<= gen_dy_cnt + '1';
						gen_dy		<= not default_out; 
					else
						gen_dy_cnt 	<= (others => '0');
						gen_dy		<= default_out; 
						trigger		<= '0';
					end if;	
				
				end if;
			end if;
		end if;
	end process;
	
END BEHV;